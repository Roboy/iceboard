// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Oct 28 20:18:56 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    inout PIN_9 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    inout PIN_10 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    inout PIN_11 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_0, PIN_7_c_1, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c, ID0, ID1, ID2, n28668;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(69[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(70[12:17])
    
    wire n16011, n16007, blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(153[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(154[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(191[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(192[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(193[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(194[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(195[22:24])
    
    wire n42330;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(196[22:24])
    
    wire n74;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(198[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(199[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(200[22:35])
    
    wire n57, n15;
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(202[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(227[22:33])
    
    wire n28891;
    wire [7:0]color_23__N_164;
    
    wire n7, n3014, n28890, n3013, n3012, n3011, n3010, n3009, 
        n3008, n3007, n4683, n3006, n3005, n3004, n28889, n3003, 
        n1158, n1157, n1156, n1155, n1154, n1153, n1152, n1151, 
        n44170, n99, n98, n97, n96, n95, n94, n93, n92, n91, 
        n90, n89, n88, n87, n6106, n6107, n6108, n6109, n6110, 
        blink_N_255, n7_adj_4310, n44421, n44420;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n41694, n41690, n41654, n41650, n28764;
    wire [31:0]motor_state_23__N_106;
    wire [24:0]displacement_23__N_229;
    wire [23:0]displacement_23__N_80;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n28888, n5999, n5998, n5997, n5996, n5995, n5994, n5993, 
        n5992, n5991, n5990, n5989, n6019, n6018, n6017, n6016, 
        n7_adj_4311, n61, n17903, n63, n59, n28667, n42324, n5952, 
        n1253;
    wire [3:0]state_3__N_362;
    
    wire n6, n7_adj_4312, n28887, n8, n9, n10;
    wire [31:0]one_wire_N_513;
    
    wire n18036, n18040, n18039, n28763, n28549, n42322, n6015, 
        n6014, n6013, n6012, n6011, n6010, n6009, n6008, n6007, 
        n6006, n6028, n6027, n18038, n18037, n6026, n6025, n1252, 
        n29030, n28886, n25555, n28666, n29029, n3002, n3001, 
        n4472, n28762, n2657, n2655, n2653, n2651, n3045, n18035, 
        n28665, n28548, n28761, n28664, n5936, n36550, n4661, 
        n3000, n86, n85, n2999, n84, n83, n82, n15_adj_4313, 
        n16, n17, n18, n19, n18034, n18033, n18032, n18031, 
        n60, n2972, n2971, n16004, n81, n80, n79, n2970, n2969, 
        n2968, n2967, n2966, n2965, n2964, n2963, n2962, n2961, 
        n2960, n2959, n2958, n2957, n2956, n2955, n2954, n2953, 
        n2952, n2951, n2950, n2949, n28760, n28885, n28759, n28758, 
        n28757, n6111, n6112, n6113, n6084, n6085, n6086, n6087, 
        n6088, n6089, n6090, n6091, n6092, n6093, n6063, n558, 
        n42898, n534, n533, n532, n531, n530, n529, n528, n527, 
        n526, n525, n524, n523, n522, n521, n520, n519, n518, 
        n517, n516, n515, n514, n513, n512, n511, n34090, n28663;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n6021, n6020, n5955, n5954, n5953, n5951, n5950, n5949, 
        n5948, n5947, n5946, n5945, n5944, n5986, n5970, n5969, 
        n5968, n5967, n5966, n54, n67, n5965, n5964, n17978, 
        n18030, n5963, n18028, n75, n5962, n5961, n5960, n510, 
        n1125, n10454, n3, n4, n5, n6_adj_4314, n7_adj_4315, n8_adj_4316, 
        n9_adj_4317, n10_adj_4318, n11, n12, n13, n14, n15_adj_4319, 
        n16_adj_4320, n17_adj_4321, n18_adj_4322, n19_adj_4323, n20, 
        n21, n22, n23, n24, n25, n28884, n28756, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n28755, n28547, n28546, n28754;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(95[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n1124, n1123, n1122, n1121, n1120, n28662, n28545, n29028, 
        n29027, n29026, n28883, n28882, n28881, n122, n123, n42310, 
        n5902, n5901, n5900, n5899, n5898, n5909, n17321, n29025, 
        n29024, n29023, n28880, n28753, n24764, n29022, n42308, 
        n28879, n29021, n29020, n29019, n29018, n28878, n29017, 
        n28877, n29016, n29015, n29014, n28544, n29013, n29012, 
        n28876, n28875, n29011, n28874, n29010, n28873, n28872, 
        n29009, n29008, n42951, n28543, n28542, n6_adj_4324, n28541, 
        n737;
    wire [31:0]\FRAME_MATCHER.state_31__N_2458 ;
    
    wire n42298, n4_adj_4325, n30501, n28871, n28540, n28870, n30500, 
        n30499, n30498, n28869, n28539, n28538, n28537, n28536, 
        n43308, n53, n64, n66, n5935, n30497, n17977, n17937, 
        n17936, n30496, n17935, n30495, n17934, n17933, n17932, 
        n30494, n29007, n17931, n17930, n16001, n29006, n28868, 
        n15998, n30493, n30492, n28535, n30491, n30490, n28534, 
        n30489, n29005, n29004, n2, n29003, n29002, n15992, n30488, 
        n29001, n30487, n30486, n29000, n30485, n35428, n30484, 
        n30483, n28999, n30482, n47, n15989, n17929, n17928, n15986, 
        n42288, n46, n42286, n24670, n30481, n30480, n30479, n30478, 
        n30477, n28998, n28997, n36403, n28996, n28995, n28994, 
        n25711, n17927, n17926, n28993, n15983, n30476, n30475, 
        n28992, n42663, n15980, n30474, n30473, n30472, n30471, 
        n17925, n17924, n35419, n38981, n28991, n28990, n43465, 
        n43463, n15962, n43462, n15959, n15953, n19634, n17923, 
        n15950, n15946, n28989, n17922, n15943, n17921, n28988, 
        n28987, n28986, n17920, n2778, n28, n42280, n42278, n2855, 
        n42665, n17919, n17918, n17917, n17916, n17915, n17914, 
        n15940, n5_adj_4326, n17913, n17912, n17911, n17910, n17909, 
        n15937, n42916, n43439, n43437, n43431, n17908, n17907, 
        n43430, n28985, n3741;
    wire [31:0]\FRAME_MATCHER.state_31__N_2586 ;
    
    wire n15933, n28984, n61_adj_4327, n97_adj_4328, n28983, n28982, 
        n28981, n2_adj_4329, n28152, n28980, n43410, n43408, n43404, 
        n20_adj_4330, n18_adj_4331, n16_adj_4332, n43403, n43434, 
        n43436, n43396, n43438, n43358, n42913, n43324, n43350, 
        n43464, n42266, n43321, n17906, n43317, n4_adj_4333, n43315, 
        n43311, n43305, n42262, n17905, n17904, n42921, n36415, 
        n15912, n43300, n43297, n42246, n14_adj_4334, n43295, \FRAME_MATCHER.i_31__N_2388 , 
        \FRAME_MATCHER.i_31__N_2390 , n17902, n17901, n17900, n17899, 
        n17898, n17897, n17896, n17895, n17894, n17893, n17892, 
        n17891, n17890, n17889, n17888, n17887, n17886, n17885, 
        n17884, n17883, n17882, n17881, n17880, n17879, n17878, 
        n17877, n17876, n17875, n17874, n17873, n17872, n17871, 
        n17870, n42923, n43385, n17869, n17868, n17867, n17866, 
        n17865, n17864, n17863, n17862, n17861, n17860, n17859, 
        n17858, n17857, n17856, n17855, n17854, n17853, n17852, 
        n17851, n17850, n17849, n17848, n17847, n17846, n17845, 
        n17844, n17843, n17842, n17841, n17840, n17839, n17838, 
        n17837, n17836, n17835, n17834, n17833, n17832, n17831, 
        n17830, n17829, n17828, n17827, n17826, n17825, n17824, 
        n17823, n17822, n17821, n17820, n17819, n17818, n17817, 
        n17816, n17815, n17814, n17813, n17812, n17811, n17810, 
        n17809, n17808, n17806, n17805, n17804, n17803, n17802, 
        n17801, n17800, n17799, n17798, n17797, n17796, n17795, 
        n17794, n17793, n17792, n17791, n17790, n17789, n17788, 
        n17787, n17786, n17785, n17784, n17783, n17782, n17781, 
        n17780, n17779, n17778, n17777, n17776, n17775, n17774, 
        n17773, n17772, n17771, n17770, n17769, n17768, n17767, 
        n17766, n17765, n17764, n17763, n17762, n17761, n17760, 
        n17759, n17758, n17757, n17756, n17755, n17754, n17753, 
        n17752, n17751, n17750, n17749, n17748, n17747, n17746, 
        n17745, n17744, n17743, n17742, n17741, n17740, n17739, 
        n17738, n17737, n17736, n17735, n17734, n17733, n17732, 
        n17731, n17730, n17729, n17728, n17727, n17726, n17725, 
        n17724, n17723, n17722, n17721, n17720, n17719, n17718, 
        n17717, n17716, n17715, n17714, n17713, n17712, n17711, 
        n17710, n17709, n17708, n17707, n17706, n17705, n17704, 
        n17703, n17702, n17701, n17700, n17699, n17698, n17697, 
        n17696, n17695, n17694, n17693, n17692, n17691, n17690, 
        n17689, n17688, n17687, n17686, n17685, n17684, n17683, 
        n17682, n17681, n17680, n17679, n17678, n17677, n17676, 
        n17675, n17674, n17673, n17672, n17671, n17670, n17669, 
        n17668, n17667, n17666, n17665, n17664, n17663, n17662, 
        n1085, n44844, n393, n392, n35416, n42920, n369, n15917, 
        n42904, n1058, n1057, n1056, n1055, n1054, n1053, n1052, 
        n17661, n249, n248, n1318, n17660, n17659, n17658, n17657, 
        n17656, n17655, n17654, n17653, n17652, n17651, n17650, 
        n17649, n17648, n17647, n17646, n17645, n1320, n1321, 
        n1325, n1322, n1323, n1324, n1319, n1283, n224, n1025, 
        n1024, n1023, n1022, n1021, n1766, n1144, n29672, n42221, 
        n29671, n20_adj_4335, n21_adj_4336, n22_adj_4337, n23_adj_4338, 
        n24_adj_4339, n29670, n29669, n29668, n25_adj_4340, n1254, 
        n1255, n1256, n1257, n1258, n8_adj_4341, n43262, n29667, 
        n28979, n28978, n28977, n28976, n17976, n17975, n29666, 
        n28975, n12_adj_4342, n65, n29665, n17974, n6_adj_4343, 
        n28974, n17973, n28973, n28972, n17972, n28971, n17971, 
        n13_adj_4344, n17970, n29664, n17969, n28970, n29663, n29662, 
        n29661, n28969, n29660, n35266, n29659, n58, n28968, n28967, 
        n28966, n28965, n28964, n28963, n68, n4401, n4400, n4399, 
        n4398, n4397, n4396, n4395, n4394, n4393, n4392, n4391, 
        n4390, n4389, n4388, n4387, n4386, n4385, n4384, n4383, 
        n4382, n4381, n69, n29658, n29657, n29656, n29655, n29654, 
        n4380, n70, n29653, n29652, n29651, n29650, n29649, n29648, 
        n29647, n7821, n47_adj_4345, n46_adj_4346, n43, n42, n40, 
        n39, n38, n17644, n17643, n17642, n17641, n17640, n17639, 
        n17638, n17637, n17636, n17635, n17634, n17633, n17632, 
        n17631, n17630, n17629, n31, n17628, n17627, n17626, n17625, 
        n17624, n17623, n17621, n17620, n17619, n17618, n17617, 
        n17616, n17615, n17614, n17613, n17612, n17611, n17610, 
        n17609, n17608, n17607, n17606, n17605, n29646, n29645, 
        quadA_debounced, quadB_debounced, count_enable, n17604, n17603, 
        n17602, n17601, n17600, n17599, n17598, n17597, n17596, 
        n17595, n17594, n4379, n4378, n6_adj_4347, n29644, n42950, 
        n29643, n29642, n29641, n5895, n5894, n5893, n43476, n986, 
        n29640, n1138, quadA_debounced_adj_4348, quadB_debounced_adj_4349, 
        count_enable_adj_4350, n29639, n29638, n17593, n29637, n29636, 
        n29635, n29634, n29633, n29632, n3022, n3021, n3020, n3019, 
        n3018, n3017, n3_adj_4351, n29631, n29630, n28962, n29629, 
        n29628, n35429, n29627, n29626, n29625, n29624, n29623, 
        n17592, n17591, n29622, n62, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n29621, n29620, n34096, n34098, n29619, n29618, n17578, 
        n17576, n17575, n17574, n29617, n29616, n17573, n17572, 
        n17571, n17570, n17569, n17566, n29615, n17563, n17561, 
        n17560, n17558, n17557, n29614, n29613, n29612, n29611, 
        n29610;
    wire [2:0]r_SM_Main_adj_5026;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_5027;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_5028;   // verilog/uart_tx.v(33[16:27])
    
    wire n28961, n29609, n29608, n29607, o_Tx_Serial_N_3351, n314, 
        n315, n43392, n43165, n29606, n29605, n29604, n17555, 
        n17554, n17552, n17551, n17549, n17548, n29603, n29602, 
        n42684, n29601, n29600, n29599, n29598, n17546, n34106, 
        n34108, n17539, n29597, n320, n17538, n29596;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15_adj_4361, n34110, n3016, n34112, n29595, n4_adj_4362;
    wire [1:0]reg_B_adj_5035;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n3015, n17531, n17529, n78, n17528, n17527, n17526, n77, 
        n29594, n17968, n17967, n17312, n17966, n11_adj_4365, n17965, 
        n29593, n43227, n28960, n17525, n71, n72, n73, n29592, 
        n29591, n28959, n17523, n17522, n17521, n17520, n17519, 
        n17518, n17517, n29590, n29589, n29588, n29587, n29586, 
        n29585, n17516, n17515, n29584, n29583, n42730, n29582, 
        n43225, n29581, n29580, n29579, n17513, n17512, n17509, 
        n43298, n29578, n29577, n29576, n29575, n4_adj_4366, n29574, 
        n35088, n29573, n29572, n29571, n29570, n29569, n29568, 
        n29567, n29566, n56, n29565, n29564, n29563, n15_adj_4367, 
        n29562, n29561, n29560, n29559, n29558, n29557, n29556, 
        n29555, n29554, n35090, n29553, n55, n29552, n1224, n42686, 
        n1225, n29551, n29550, n29549, n29548, n29547, n29546, 
        n29545, n1221, n1222, n29544, n29543, n1223, n1220, n29542, 
        n29541, n4_adj_4368, n29540, n1219, n29539, n5_adj_4369, 
        n4_adj_4370, n3_adj_4371, n29538, n29537, n29536, n29535, 
        n29534, n29533, n29532, n29531, n29530, n29529, n29528, 
        n29527, n29526, n29525, n29524, n15_adj_4372, n5934, n29523, 
        n29522, n29521, n29520, n29519, n29518, n43302, n28958, 
        n29517, n29516, n29515, n34114, n29514, n29513, n17481, 
        n8_adj_4373, n9_adj_4374, n10_adj_4375, n11_adj_4376, n12_adj_4377, 
        n13_adj_4378, n14_adj_4379, n15_adj_4380, n16_adj_4381, n17_adj_4382, 
        n18_adj_4383, n19_adj_4384, n20_adj_4385, n21_adj_4386, n22_adj_4387, 
        n23_adj_4388, n24_adj_4389, n25_adj_4390, n17964, n43306, 
        n6153, n6154, n6155, n6156, n6129, n6130, n6131, n6132, 
        n6133, n6134, n958, n957, n956, n955, n954, n953, n43309, 
        n648, n649, n43202, n671, n672, n43200, n43198, n43312, 
        n43314, n783, n784, n785, n806, n807, n43192, n43190, 
        n43384, n43187, n28957, n28956, n914, n915, n916, n917, 
        n918, n28955, n28954, n938, n939, n28953, n29512, n29511, 
        n855, n852, n28952, n42911, n1043, n1044, n1045, n1046, 
        n1047, n1048, n29510, n43320, n1067, n1068, n29509, n29508, 
        n28951, n28950, n43150, n1169, n1170, n1171, n1172, n1173, 
        n1174, n1175, n1193, n1194, n5910, n5911, n5912, n5913, 
        n5914, n5915, n5916, n8_adj_4391, n28949, n43174, n28948, 
        n29507, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
        n1299, n43322, n1316, n1317, n15922, n749, n748, n746, 
        n43170, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
        n1419, n1420, n18_adj_4392, n1436, n1437, n16_adj_4393, 
        n44174, n44177, n44180, n44183, n44186, n3459, n3458, 
        n3457, n3456, n3455, n36486, n5938, n5939, n5940, n5941, 
        n13_adj_4394, n29506, n3452, n3453, n3454, n28947, n1529, 
        n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
        n1538, n17963, n28946, n1553, n1554, n28945, n43166, n43164, 
        n42910, n29505, n29504, n1643, n1644, n1645, n1646, n1647, 
        n1648, n1649, n1650, n1651, n1652, n1653, n43163, n43160, 
        n1667, n1668, n29503, n43158, n43156, n29502, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n3362, n29501, n3358, n3357, n3356, n3355, 
        n3354, n3353, n1778, n1779, n28944, n3346, n3345, n3344, 
        n3343, n3342, n5973, n5974, n5975, n5976, n5977, n5978, 
        n5979, n5980, n5981, n5982, n5983, n5984, n5985, n3330, 
        n3337, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
        n1869, n1870, n1871, n1872, n1873, n1874, n3325, n3324, 
        n3323, n3322, n3321, n3320, n3319, n1886, n1887, n43155, 
        n43326, n3317, n3316, n3315, n3314, n3313, n3312, n3311, 
        n3310, n3309, n3308, n42924, n6000, n6001, n6002, n6003, 
        n43149, n29500, n3299, n3300, n3301, n3302, n3303, n3304, 
        n3305, n3306, n3307, n1967, n1968, n1969, n1970, n1971, 
        n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n3298, n1991, n1992, n43145, n42145, n35269, n2069, 
        n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
        n2078, n2079, n2080, n2081, n2082, n2083, n3263, n2093, 
        n2094, n3258, n3257, n3256, n3255, n3254, n3253, n3252, 
        n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, 
        n6037, n6038, n6039, n6040, n6060, n3245, n3246, n3247, 
        n3248, n3249, n3250, n3251, n2168, n2169, n2170, n2171, 
        n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
        n2180, n2181, n2182, n2183, n3244, n3243, n3242, n3241, 
        n3240, n3239, n3238, n3237, n2192, n2193, n36527, n36517, 
        n6_adj_4395, n4_adj_4396, n3235, n3234, n3233, n3232, n3231, 
        n3230, n29499, n6043, n6044, n6045, n6046, n6047, n6048, 
        n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, 
        n6057, n6058, n6059, n3223, n3224, n3225, n29498, n2264, 
        n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
        n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
        n3222, n3221, n3220, n3219, n3218, n3217, n3216, n2288, 
        n2289, n3214, n3213, n3212, n3211, n3210, n3209, n29497, 
        n29496, n6064, n6065, n6066, n6067, n6068, n6069, n6070, 
        n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, 
        n6079, n6080, n6081, n3204, n3205, n3206, n3207, n3208, 
        n29495, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
        n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, 
        n2372, n2373, n2374, n3203, n3202, n3201, n3200, n3199, 
        n2381, n2382, n36500, n6094, n6095, n6096, n6097, n6098, 
        n6099, n6100, n6101, n6102, n6103, n2447, n2448, n2449, 
        n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
        n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
        n2471, n2472, n36470, n29494, n6114, n6115, n6116, n6117, 
        n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
        n6126, n29493, n2534, n2535, n2536, n2537, n2538, n2539, 
        n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
        n2548, n2549, n2550, n2551, n2552, n2553, n2558, n2559, 
        n29492, n29491, n36533, n6135, n6136, n6137, n6138, n6139, 
        n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
        n6148, n6149, n6150, n3164, n2618, n2619, n2620, n2621, 
        n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
        n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
        n2638, n29490, n2642, n2643, n29489, n3158, n36401, n6157, 
        n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
        n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
        n6174, n6175, n29488, n3157, n2699, n2700, n2701, n2702, 
        n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
        n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
        n2719, n2720, n3156, n3155, n2723, n2724, n8_adj_4397, 
        n7_adj_4398, n3154, n29487, n3153, n2777, n2798, n2799, 
        n3152, n2801, n2802, n29486, n36444, n29485, n29484, n28943, 
        n42830, n106, n35268, n29483, n29482, n3150, n3149, n3148, 
        n3147, n3146, n3145, n3144, n3143, n3142, n3141, n3140, 
        n3139, n3138, n3137, n3136, n3135, n3134, n3133, n3132, 
        n3131, n29481, n28942, n29480, n36571, n29479, n29478, 
        n29477, n29476, n29475, n29474, n29473, n3125, n29472, 
        n3124, n3123, n29471, n29470, n3122, n3121, n29469, n3120, 
        n3119, n3118, n3117, n29468, n3116, n3115, n29467, n29466, 
        n3114, n3113, n3112, n29465, n18165, n18161, n18160, n18159, 
        n18158, n18157, n18156, n18155, n18154, n18153, n18152, 
        n18151, n18150, n18149, n18148, n18147, n18146, n18145, 
        n18144, n18143, n18142, n18141, n18140, n18139, n5905, 
        n3111, n3110, n3109, n3108, n3107, n3106, n3105, n3104, 
        n29464, n3103, n3102, n3101, n3100, n29463, n18138, n18137, 
        n18136, n18135, n18134, n18133, n18132, n18131, n18130, 
        n32680, n32678, n18125, n18124, n18123, n18122, n32662, 
        n32660, n34084, n34082, n18111, n18108, n29462, n29461, 
        n29460, n29459, n29458, n29457, n29456, n29455, n29454, 
        n18105, n18101, n18097, n18096, n18095, n18094, n18093, 
        n18092, n18091, n18090, n18089, n18088, n18087, n18086, 
        n18085, n18084, n18083, n18082, n18081, n18080, n18079, 
        n18078, n18077, n18076, n63_adj_4399, n5904, n5903, n29453, 
        n18075, n35417, n18072, n18071, n18070, n18069, n18068, 
        n18067, n18066, n18065, n3065, n18064, n29452, n18063, 
        n18062, n18061, n18060, n18059, n18058, n18057, n18056, 
        n3058, n18055, n3057, n18054, n3056, n18053, n3055, n18052, 
        n3054, n18051, n3053, n18050, n3052, n18049, n3051, n18048, 
        n3050, n18047, n3049, n18046, n3048, n3047, n18045, n29451, 
        n3046, n18044, n1251, n3044, n1250, n3043, n18043, n3042, 
        n18042, n3041, n18041, n3040, n3039, n3038, n3037, n3036, 
        n28941, n3035, n3034, n3033, n3032, n28940, n28939, n28938, 
        n28937, n28936, n28935, n28934, n17466, n29450, n1184, 
        n29449, n28933, n17186, n17180, n17962, n17961, n17960, 
        n17959, n17958, n17957, n17956, n17463, n29448, n2966_adj_4400, 
        n29447, n2958_adj_4401, n2957_adj_4402, n2956_adj_4403, n2955_adj_4404, 
        n2954_adj_4405, n2953_adj_4406, n2952_adj_4407, n28932, n28931, 
        n17159, n28930, n34116, n28929, n28813, n34118, n28812, 
        n2951_adj_4408, n2950_adj_4409, n2949_adj_4410, n2948, n2947, 
        n2946, n2945, n2944, n2943, n2942, n2941, n2940, n2939, 
        n2938, n2937, n2936, n2935, n2934, n2933, n2925, n2924, 
        n2923, n2922, n34120, n28811, n17108, n17100, n29446, 
        n29445, n29444, n29443, n29442, n17955, n43025, n36306, 
        n38007, n28810, n28928, n34122, n43022, n17068, n29441, 
        n28809, n34124, n17058, n28927, n42744, n28808, n43016, 
        n28926, n32, n31_adj_4411, n30, n28925, n43010, n29, n28_adj_4412, 
        n43006, n43151, n28924, n28923, n33, n32_adj_4413, n31_adj_4414, 
        n30_adj_4415, n29_adj_4416, n28_adj_4417, n27, n26, n25_adj_4418, 
        n24_adj_4419, n23_adj_4420, n22_adj_4421, n21_adj_4422, n20_adj_4423, 
        n19_adj_4424, n18_adj_4425, n17_adj_4426, n16_adj_4427, n15_adj_4428, 
        n14_adj_4429, n13_adj_4430, n12_adj_4431, n11_adj_4432, n10_adj_4433, 
        n29440, n2921, n2920, n29439, n2919, n29438, n2918, n2917, 
        n2916, n2915, n2914, n2913, n2912, n2911, n2910, n2909, 
        n2908, n2907, n2906, n2905, n2904, n2903, n2902, n2867, 
        n29437, n29436, n29435, n29434, n29433, n29432, n42113, 
        n2858, n2857, n2856, n2855_adj_4434, n2854, n2853, n2852, 
        n2851, n2850, n2849, n2848, n2847, n2846, n2845, n2844, 
        n2843, n2842, n2841, n2840, n2839, n2838, n2837, n2836, 
        n2835, n2834, n2825, n2824, n2823, n2822, n2821, n2820, 
        n2819, n2818, n2817, n2816, n2815, n2814, n2813, n2812, 
        n2811, n2810, n2809, n2808, n2807, n2806, n2805, n2804, 
        n2803, n43003, n29431, n29430, n42702, n2768, n29429, 
        n2758, n2757, n2756, n2755, n2754, n2753, n2752, n2751, 
        n2750, n2749, n2748, n2747, n2746, n2745, n2744, n2743, 
        n2742, n2741, n2740, n2739, n2738, n2737, n2736, n2735, 
        n29428, n41591, n29427, n2725, n2724_adj_4435, n2723_adj_4436, 
        n2722, n2721, n2720_adj_4437, n2719_adj_4438, n2718_adj_4439, 
        n2717_adj_4440, n2716_adj_4441, n2715_adj_4442, n2714_adj_4443, 
        n2713_adj_4444, n2712_adj_4445, n2711_adj_4446, n2710_adj_4447, 
        n2709_adj_4448, n2708_adj_4449, n2707_adj_4450, n2706_adj_4451, 
        n2705_adj_4452, n2704_adj_4453, n29426, n36199, n1714, n1746, 
        n1715, n1747, n1716, n1748, n1717, n1749, n1718, n1750, 
        n1719, n1751, n1720, n1752, n1721, n1753, n1722, n1754_adj_4454, 
        n1723, n1755_adj_4455, n1724, n1756_adj_4456, n1725, n1757_adj_4457, 
        n1758_adj_4458, n28922, n28921, n28800, n29425, n29424, 
        n28799, n36545, n28798, n1745, n3151, n134, n135, n136, 
        n137, n138, n139, n140, n141, n142, n143, n144, n145, 
        n146, n147, n148, n149, n150, n151, n152, n153, n154, 
        n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165, n1652_adj_4459, n1653_adj_4460, n1654, n1655, 
        n1656, n1657, n1658, n29423, n29422, n29421, n28797, n29420, 
        n29419, n29418, n1679, n1621, n1622, n1623, n1624, n1625, 
        n28920, n28919, n4_adj_4461, n29417, n1646_adj_4462, n1647_adj_4463, 
        n1648_adj_4464, n1649_adj_4465, n1650_adj_4466, n1651_adj_4467, 
        n2669, n5_adj_4468, n29416, n9_adj_4469, n8_adj_4470, n7_adj_4471, 
        n6_adj_4472, n5_adj_4473, n4_adj_4474, n3_adj_4475, n28918, 
        n29415, n29414, n2658, n29413, n2656, n29412, n2654, n29411, 
        n2652, n28796, n2650, n2649, n2648, n2647, n2646, n2645, 
        n2644, n2643_adj_4476, n2642_adj_4477, n2641, n2640, n2639, 
        n2638_adj_4478, n2637_adj_4479, n2636_adj_4480, n29410, n28795, 
        n5928, n5927, n5926, n5925, n5924, n5923, n2625_adj_4481, 
        n5922, n2624_adj_4482, n5921, n2623_adj_4483, n5920, n2622_adj_4484, 
        n5919, n2621_adj_4485, n5937, n2620_adj_4486, n1547, n1548, 
        n1549, n1550, n1551, n1552, n1553_adj_4487, n1554_adj_4488, 
        n1555, n1556, n1557, n2617, n28794, n1558, n29409, n13_adj_4489, 
        n29408, n41571, n29407, n29406, n28917, n29405, n1580, 
        n1615, n41561, n1616, n11_adj_4490, n1617, n1618, n1619, 
        n1620, n2618_adj_4491, n2619_adj_4492, n41545, n41542, n1516, 
        n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
        n1525, n29404, n2616, n29403, n29402, n28916, n29401, 
        n1481, n2615, n28793, n29400, n2611, n1454, n1455, n28915, 
        n1456, n1457, n29399, n1458, n1448, n1449, n1450, n29398, 
        n1451, n1452, n1453, n2614, n2612, n2613, n34092, n34094, 
        n17390, n17389, n34126, n34128, n34130, n42993, n2608, 
        n1417_adj_4493, n1418_adj_4494, n1419_adj_4495, n1420_adj_4496, 
        n1421, n1422, n1423, n1424, n28914, n1425, n2609, n2610, 
        n29397, n1382, n2607, n34132, n34134, n34136, n34138, 
        n34140, n34142, n34144, n34146, n1358, n2606, n2605, n34148, 
        n1356, n1357, n1350, n1351, n1354, n1352, n1355, n1353, 
        n34150, n1349, n5933, n42712, n42097, n2570, n29396, n28913, 
        n29395, n29394, n2558_adj_4497, n2557, n2556, n2555, n2554, 
        n2553_adj_4498, n2552_adj_4499, n2551_adj_4500, n29393, n2550_adj_4501, 
        n2549_adj_4502, n2548_adj_4503, n2547_adj_4504, n2546_adj_4505, 
        n2545_adj_4506, n2544_adj_4507, n2543_adj_4508, n2542_adj_4509, 
        n2541_adj_4510, n2540_adj_4511, n2539_adj_4512, n2538_adj_4513, 
        n2537_adj_4514, n5932, n28912, n2525, n2524, n2523, n2522, 
        n2521, n2520, n2519, n2518, n2517, n2516, n2515, n2514, 
        n2513, n2512, n2511, n2510, n2509, n2508, n2507, n2506, 
        n42988, n42704, n2471_adj_4515, n29392, n28911, n29391, 
        n29390, n2458_adj_4516, n2457_adj_4517, n2456_adj_4518, n2_adj_4519, 
        n3_adj_4520, n4_adj_4521, n5_adj_4522, n6_adj_4523, n7_adj_4524, 
        n8_adj_4525, n9_adj_4526, n10_adj_4527, n11_adj_4528, n12_adj_4529, 
        n13_adj_4530, n14_adj_4531, n15_adj_4532, n16_adj_4533, n17_adj_4534, 
        n18_adj_4535, n19_adj_4536, n20_adj_4537, n21_adj_4538, n22_adj_4539, 
        n23_adj_4540, n24_adj_4541, n25_adj_4542, n2_adj_4543, n3_adj_4544, 
        n4_adj_4545, n5_adj_4546, n6_adj_4547, n7_adj_4548, n8_adj_4549, 
        n9_adj_4550, n10_adj_4551, n11_adj_4552, n12_adj_4553, n13_adj_4554, 
        n14_adj_4555, n15_adj_4556, n16_adj_4557, n17_adj_4558, n18_adj_4559, 
        n19_adj_4560, n20_adj_4561, n21_adj_4562, n22_adj_4563, n23_adj_4564, 
        n24_adj_4565, n25_adj_4566, n5959, n2455_adj_4567, n2454_adj_4568, 
        n2453_adj_4569, n2452_adj_4570, n2451_adj_4571, n2450_adj_4572, 
        n2449_adj_4573, n2448_adj_4574, n2447_adj_4575, n2446, n2445, 
        n2444, n2443, n2442, n2441, n2440, n2439, n2438, n28910, 
        n29389, n2425, n2424, n2423, n2422, n2421, n2420, n2419, 
        n2418, n2417, n2416, n2415, n29388, n46_adj_4576, n2414, 
        n2413, n2412, n2411, n2410, n2409, n2408, n2407, n29387, 
        n29386, n2372_adj_4577, n29385, n29384, n2358_adj_4578, n2357_adj_4579, 
        n2356, n2355, n2354, n29383, n44, n42716, n2353, n2352, 
        n2351, n2350, n2349, n2348, n2347, n2346, n42983, n2345, 
        n2344, n2343, n2342, n2341, n2340, n2339, n2325, n2324, 
        n2323, n2322, n2321, n2320, n2319, n2318, n2317, n2316, 
        n2315, n2314, n2313, n2312, n2311, n2310, n2309, n2308, 
        n29382, n42_adj_4580, n42981, n43159, n2273_adj_4581, n29381, 
        n42087, n2258, n2257, n2256, n2255, n2254, n2253, n2252, 
        n2251, n2250, n2249, n2248, n2247, n2246, n2245, n2244, 
        n2243, n2242, n29380, n40_adj_4582, n42_adj_4583, n44_adj_4584, 
        n45, n2241, n2240, n29379, n29378, n29377, n29376, n29375, 
        n2225, n2224, n2223, n2222, n2221, n2220, n2219, n2218, 
        n2217, n2216, n2215, n2214, n2213, n2212, n2211, n2210, 
        n2209, n29374, n38_adj_4585, n40_adj_4586, n42_adj_4587, n43_adj_4588, 
        n42722, n43169, n2174_adj_4589, n29373, n29372, n29371, 
        n2158, n2157, n2156, n2155, n2154, n2153, n2152, n2151, 
        n2150, n2149, n2148, n2147, n2146, n2145, n2144, n2143, 
        n2142, n29370, n36, n38_adj_4590, n40_adj_4591, n41, n43211, 
        n2141, n29369, n2125, n2124, n2123, n2122, n2121, n2120, 
        n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, 
        n2111, n2110, n43473, n29368, n41493, n34, n36_adj_4592, 
        n38_adj_4593, n39_adj_4594, n41_adj_4595, n43_adj_4596, n44_adj_4597, 
        n45_adj_4598, n42724, n42736, n2075_adj_4599, n29367, n42073, 
        n29366, n2058, n2057, n2056, n2055, n2054, n29365, n32_adj_4600, 
        n34_adj_4601, n37, n39_adj_4602, n41_adj_4603, n43_adj_4604, 
        n2053, n2052, n2051, n2050, n2049, n2048, n2047, n2046, 
        n2045, n2044, n2043, n2042, n36407, n2025, n2024, n2023, 
        n2022, n2021, n2020, n2019, n2018, n2017, n2016, n2015, 
        n29364, n30_adj_4605, n31_adj_4606, n32_adj_4607, n33_adj_4608, 
        n34_adj_4609, n35, n37_adj_4610, n39_adj_4611, n43157, n41_adj_4612, 
        n42_adj_4613, n43_adj_4614, n45_adj_4615, n2014, n2013, n2012, 
        n2011, n29363, n29362, n28_adj_4616, n29_adj_4617, n30_adj_4618, 
        n31_adj_4619, n32_adj_4620, n33_adj_4621, n35_adj_4622, n37_adj_4623, 
        n39_adj_4624, n40_adj_4625, n41_adj_4626, n43_adj_4627, n1976_adj_4628, 
        n29361, n29360, n29359, n29358, n29357, n29356, n1958, 
        n1957, n1956, n1955, n1954, n1953, n1952, n1951, n1950, 
        n1949, n1948, n1947, n1946, n1945, n29355, n26_adj_4629, 
        n27_adj_4630, n28_adj_4631, n29_adj_4632, n30_adj_4633, n31_adj_4634, 
        n33_adj_4635, n35_adj_4636, n37_adj_4637, n38_adj_4638, n39_adj_4639, 
        n41_adj_4640, n1944, n1943, n29354, n3351, n29353, n29352, 
        n1925, n1924, n1923, n1922, n1921, n1920, n1919, n1918, 
        n1917, n1916, n1915, n29351, n41477, n24_adj_4641, n25_adj_4642, 
        n26_adj_4643, n27_adj_4644, n28_adj_4645, n29_adj_4646, n30_adj_4647, 
        n31_adj_4648, n32_adj_4649, n33_adj_4650, n35_adj_4651, n36_adj_4652, 
        n37_adj_4653, n39_adj_4654, n42990, n42992, n1914, n1913, 
        n1912, n3318, n29350, n41475, n22_adj_4655, n23_adj_4656, 
        n24_adj_4657, n25_adj_4658, n26_adj_4659, n27_adj_4660, n28_adj_4661, 
        n29_adj_4662, n30_adj_4663, n31_adj_4664, n33_adj_4665, n34_adj_4666, 
        n35_adj_4667, n37_adj_4668, n39_adj_4669, n43201, n41_adj_4670, 
        n43_adj_4671, n42998, n43221, n1877, n29349, n29348, n29347, 
        n29346, n29345, n29344, n29343, n20_adj_4672, n21_adj_4673, 
        n22_adj_4674, n23_adj_4675, n24_adj_4676, n25_adj_4677, n26_adj_4678, 
        n27_adj_4679, n28_adj_4680, n29_adj_4681, n31_adj_4682, n32_adj_4683, 
        n33_adj_4684, n35_adj_4685, n37_adj_4686, n43310, n39_adj_4687, 
        n41_adj_4688, n29342, n1858, n1857, n1856, n1855, n1854, 
        n1853, n1852, n1851, n1850, n1849, n1848, n1847, n1846, 
        n1845, n1844, n29341, n41470, n18_adj_4689, n19_adj_4690, 
        n20_adj_4691, n21_adj_4692, n22_adj_4693, n23_adj_4694, n24_adj_4695, 
        n25_adj_4696, n26_adj_4697, n27_adj_4698, n29_adj_4699, n30_adj_4700, 
        n31_adj_4701, n33_adj_4702, n35_adj_4703, n37_adj_4704, n39_adj_4705, 
        n41_adj_4706, n43_adj_4707, n45_adj_4708, n43000, n29340, 
        n29339, n29338, n29337, n3236, n29336, n29335, n1825, 
        n1824, n29334, n16_adj_4709, n17_adj_4710, n18_adj_4711, n19_adj_4712, 
        n20_adj_4713, n21_adj_4714, n22_adj_4715, n23_adj_4716, n25_adj_4717, 
        n27_adj_4718, n28_adj_4719, n29_adj_4720, n31_adj_4721, n33_adj_4722, 
        n43316, n35_adj_4723, n37_adj_4724, n39_adj_4725, n41_adj_4726, 
        n43_adj_4727, n1823, n1822, n1821, n1820, n1819, n1818, 
        n3215, n1817, n1816, n1815, n1814, n1813, n29333, n41466, 
        n14_adj_4728, n16_adj_4729, n17_adj_4730, n18_adj_4731, n19_adj_4732, 
        n20_adj_4733, n21_adj_4734, n22_adj_4735, n23_adj_4736, n25_adj_4737, 
        n26_adj_4738, n27_adj_4739, n29_adj_4740, n31_adj_4741, n33_adj_4742, 
        n35_adj_4743, n37_adj_4744, n43148, n39_adj_4745, n40_adj_4746, 
        n41_adj_4747, n43_adj_4748, n45_adj_4749, n43223, n43407, 
        n29332, n12_adj_4750, n14_adj_4751, n15_adj_4752, n16_adj_4753, 
        n17_adj_4754, n18_adj_4755, n19_adj_4756, n20_adj_4757, n21_adj_4758, 
        n23_adj_4759, n24_adj_4760, n25_adj_4761, n27_adj_4762, n29_adj_4763, 
        n31_adj_4764, n33_adj_4765, n35_adj_4766, n43144, n37_adj_4767, 
        n38_adj_4768, n39_adj_4769, n41_adj_4770, n43_adj_4771, n43142, 
        n37_adj_4772, n29331, n10_adj_4773, n12_adj_4774, n13_adj_4775, 
        n14_adj_4776, n15_adj_4777, n16_adj_4778, n17_adj_4779, n18_adj_4780, 
        n19_adj_4781, n21_adj_4782, n22_adj_4783, n23_adj_4784, n25_adj_4785, 
        n27_adj_4786, n29_adj_4787, n31_adj_4788, n33_adj_4789, n43136, 
        n35_adj_4790, n36_adj_4791, n37_adj_4792, n39_adj_4793, n41_adj_4794, 
        n43230, n29330, n8_adj_4795, n10_adj_4796, n11_adj_4797, n12_adj_4798, 
        n13_adj_4799, n14_adj_4800, n15_adj_4801, n16_adj_4802, n17_adj_4803, 
        n19_adj_4804, n20_adj_4805, n21_adj_4806, n23_adj_4807, n25_adj_4808, 
        n43132, n27_adj_4809, n29_adj_4810, n31_adj_4811, n32_adj_4812, 
        n33_adj_4813, n34_adj_4814, n35_adj_4815, n37_adj_4816, n39_adj_4817, 
        n43027, n1778_adj_4818, n29329, n35_adj_4819, n6_adj_4820, 
        n8_adj_4821, n9_adj_4822, n10_adj_4823, n11_adj_4824, n12_adj_4825, 
        n13_adj_4826, n14_adj_4827, n15_adj_4828, n17_adj_4829, n19_adj_4830, 
        n21_adj_4831, n23_adj_4832, n42922, n25_adj_4833, n27_adj_4834, 
        n29_adj_4835, n31_adj_4836, n32_adj_4837, n33_adj_4838, n35_adj_4839, 
        n37_adj_4840, n29328, n29327, n4_adj_4841, n6_adj_4842, n7_adj_4843, 
        n8_adj_4844, n9_adj_4845, n10_adj_4846, n11_adj_4847, n12_adj_4848, 
        n13_adj_4849, n15_adj_4850, n16_adj_4851, n17_adj_4852, n19_adj_4853, 
        n21_adj_4854, n42912, n23_adj_4855, n24_adj_4856, n25_adj_4857, 
        n27_adj_4858, n29_adj_4859, n30_adj_4860, n31_adj_4861, n33_adj_4862, 
        n35_adj_4863, n37_adj_4864, n39_adj_4865, n41_adj_4866, n43_adj_4867, 
        n45_adj_4868, n34_adj_4869, n32_adj_4870, n17954, n31_adj_4871, 
        n29326, n29325, n17330, n29324, n28909, n29323, n29322, 
        n5890, n5891, n5892, n5881, n5882, n5883, n5884, n5885, 
        n5886, n17953, n17952, n29321, n29320, n13293, n29319, 
        n6_adj_4872, n16_adj_4873, n11_adj_4874, n10_adj_4875, n29318, 
        n29317, n25_adj_4876, n35086, n29316, n29315, n29314, n29313, 
        n29312, n29311, n29310, n29309, n44_adj_4877, n43_adj_4878, 
        n29308, n42_adj_4879, n29307, n29306, n29305, n29304, n41_adj_4880, 
        n39_adj_4881, n38_adj_4882, n42752, n10223, n10222, n10221, 
        n10220, n10219, n31_adj_4883, n10218, n26_adj_4884, n30_adj_4885, 
        n29_adj_4886, n28_adj_4887, n27_adj_4888, n25741, n42040, 
        n18_adj_4889, n28908, n19_adj_4890, n34088, n34104, n41435, 
        n11_adj_4891, n41429, n34080, n5_adj_4892, n42357, n42742, 
        n41999, n34_adj_4893, n33_adj_4894, n32_adj_4895, n31_adj_4896, 
        n30_adj_4897, n29280, n29279, n29278, n29277, n29276, n29275, 
        n29274, n41986, n41984, n29273, n29272, n25771, n43458, 
        n13_adj_4898, n35423, n34728, n11_adj_4899, n41423, n41417, 
        n17951, n18027, n17939, n41980, n41409, n42551, n41962, 
        n29271, n15977, n41960, n42756, n35418, n41958, n41956, 
        n41945, n41943, n6_adj_4900, n41937, n41934, n15930, n29270, 
        n42403, n29269, n29268, n29267, n29266, n35435, n35434, 
        n35433, n35432, n12_adj_4901, n29265, n43478, n17950, n29264, 
        n29263, n28_adj_4902, n27_adj_4903, n41915, n35431, n26_adj_4904, 
        n25_adj_4905, n42535, n41407, n43067, n29262, n29261, n41907, 
        n28907, n41405, n35430, n35422, n41903, n22916, n41897, 
        n29260, n29259, n35421, n4_adj_4906, n41891, n12_adj_4907, 
        n35420, n6_adj_4908, n42411, n41872, n29258, n42377, n17949, 
        n17240, n42415, n29257, n28906, n39157, n29256, n29255, 
        n29254, n29253, n1, n32676, n17948, n17947, n17946, n41397, 
        n17945, n41852, n41850, n41846, n41844, n43081, n43367, 
        n39099, n41842, n28905, n42405, n17944, n28_adj_4909, n26_adj_4910, 
        n2_adj_4911, n41393, n24_adj_4912, n38949, n41826, n19_adj_4913, 
        n38945, n16_adj_4914, n43137, n41818, n41806, n41804, n43133, 
        n41798, n41796, n41794, n43364, n43479, n43131, n43362, 
        n43366, n43477, n41747, n41739, n5889, n5908, n43089, 
        n5931, n41313, n5958, n41310, n6024, n41301, n41299, n41389, 
        n41297, n41296, n41295, n41363, n41294, n41293, n41355, 
        n41347, n41345, n41292, n41291, n43370, n41290, n41289, 
        n41288, n41343, n41287, n41286, n43383, n41285, n41284, 
        n41283, n17938, n41282, n41281, n41280, n41279, n41278, 
        n41277, n41276, n41275, n41274, n41273, n41272, n17943, 
        n28904, n28903, n43130, n41271, n17942, n41270, n28902, 
        n41269, n41268, n26_adj_4915, n41267, n24_adj_4916, n22_adj_4917, 
        n18_adj_4918, n41266, n36397, n43097, n2_adj_4919, n2_adj_4920, 
        n3_adj_4921, n4_adj_4922, n5_adj_4923, n6_adj_4924, n7_adj_4925, 
        n8_adj_4926, n9_adj_4927, n10_adj_4928, n11_adj_4929, n12_adj_4930, 
        n13_adj_4931, n14_adj_4932, n15_adj_4933, n16_adj_4934, n17_adj_4935, 
        n18_adj_4936, n19_adj_4937, n20_adj_4938, n21_adj_4939, n22_adj_4940, 
        n23_adj_4941, n24_adj_4942, n25_adj_4943, n26_adj_4944, n27_adj_4945, 
        n28_adj_4946, n29_adj_4947, n30_adj_4948, n31_adj_4949, n32_adj_4950, 
        n33_adj_4951, n36457, n29211, n29210, n29209, n29208, n29207, 
        n29206, n28901, n29205, n29204, n29203, n38783, n29202, 
        n29201, n29200, n28900, n541, n28683, n29199, n29198, 
        n35374, n29197, n29196, n29195, n28682, n28899, n28898, 
        n29194, n29193, n29192, n29191, n28775, n29190, n29189, 
        n29188, n28681, n29187, n29186, n29185, n41339, n29184, 
        n29183, n29182, n29181, n43129, n29180, n29179, n29178, 
        n29177, n43380, n32658, n29176, n29175, n29174, n29173, 
        n29172, n29171, n29170, n36480, n29169, n29168, n29167, 
        n29166, n29165, n38755, n29164, n42_adj_4952, n41_adj_4953, 
        n40_adj_4954, n39_adj_4955, n37_adj_4956, n41248, n36_adj_4957, 
        n29163, n29162, n29161, n29160, n29159, n41247, n29158, 
        n29157, n29_adj_4958, n42942, n29156, n29155, n36512, n29154, 
        n29153, n40_adj_4959, n39_adj_4960, n29152, n38_adj_4961, 
        n37_adj_4962, n36_adj_4963, n29151, n34_adj_4964, n29150, 
        n29149, n26_adj_4965, n29148, n29147, n29146, n29145, n29144, 
        n29143, n29142, n29141, n28774, n38_adj_4966, n29140, n37_adj_4967, 
        n29139, n29138, n29137, n36_adj_4968, n35_adj_4969, n33_adj_4970, 
        n29136, n29135, n29134, n28680, n29133, n10_adj_4971, n29132, 
        n29131, n29130, n26_adj_4972, n29129, n38713, n29128, n29127, 
        n22_adj_4973, n29126, n29125, n29124, n29123, n29122, n29121, 
        n29120, n29119, n29118, n29117, n29116, n29115, n28679, 
        n43375, n29114, n29113, n28773, n29112, n36865, n29111, 
        n29110, n42943, n43379, n24_adj_4974, n22_adj_4975, n29109, 
        n29108, n20_adj_4976, n43475, n28678, n16_adj_4977, n29107, 
        n29106, n28677, n29105, n29104, n28897, n29103, n29102, 
        n29101, n28896, n28772, n28676, n36579, n29100, n42375, 
        n29099, n29098, n29097, n29096, n29095, n28771, n28675, 
        n36465, n28674, n29094, n28770, n38657, n29093, n28895, 
        n29092, n29091, n29090, n29089, n28769, n36584, n28673, 
        n29088, n29087, n38651, n29086, n28894, n36482, n29085, 
        n29084, n29083, n29082, n36450, n29081, n29080, n28768, 
        n36409, n29079, n18029, n29078, n29077, n29076, n29075, 
        n28767, n29074, n29073, n28672, n29072, n29071, n28893, 
        n38647, n29070, n28671, n28766, n37457, n29069, n29068, 
        n29067, n29066, n36441, n29065, n29064, n29063, n29062, 
        n29061, n29060, n29059, n29058, n28892, n29057, n29056, 
        n29055, n29054, n29053, n29052, n29051, n28765, n29050, 
        n29049, n29048, n29047, n29046, n29045, n29044, n29043, 
        n29042, n29041, n29040, n29039, n29038, n29037, n29036, 
        n29035, n29034, n28670, n29033, n28669, n29032, n17941, 
        n29031, n17940, n38623, n38621, n38619, n38617, n38615, 
        n38613, n39151, n43376, n43105, n41204, n34716, n41329, 
        n40_adj_4978, n35271, n16_adj_4979, n5_adj_4980, n4_adj_4981, 
        n38565, n38563, n38561, n38059, n38559, n38557, n38551, 
        n39142, n38537, n44233, n34804, n35274, n41327, n38531, 
        n36217, n38525, n36850, n38986, n38509, n42975, n38495, 
        n38491, n39138, n38485, n43390, n38465, n38463, n34912, 
        n35270, n42884, n43389, n41323, n42890, n44228, n44224, 
        n35000, n35273, n35004, n35275, n36563, n36429, n38107, 
        n42605, n41321, n35272, n35276, n22_adj_4982, n19_adj_4983, 
        n18_adj_4984, n15_adj_4985, n36325, n36299, n37455, n37799, 
        n42972, n36150, n36148, n36146, n42627;
    
    VCC i2 (.Y(VCC_net));
    SB_IO ID1_input (.PACKAGE_PIN(PIN_10), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(ID1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID1_input.PIN_TYPE = 6'b000001;
    defparam ID1_input.PULLUP = 1'b1;
    defparam ID1_input.NEG_TRIGGER = 1'b0;
    defparam ID1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO ID2_input (.PACKAGE_PIN(PIN_11), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(ID2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID2_input.PIN_TYPE = 6'b000001;
    defparam ID2_input.PULLUP = 1'b1;
    defparam ID2_input.NEG_TRIGGER = 1'b0;
    defparam ID2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 div_46_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_1720_7 (.CI(n29479), .I0(n2554), .I1(GND_net), 
            .CO(n29480));
    SB_DFF h2_56 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_57 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF dir_61 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_IO ID0_input (.PACKAGE_PIN(PIN_9), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(ID0)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID0_input.PIN_TYPE = 6'b000001;
    defparam ID0_input.PULLUP = 1'b1;
    defparam ID0_input.NEG_TRIGGER = 1'b0;
    defparam ID0_input.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .bit_ctr({bit_ctr}), .VCC_net(VCC_net), 
            .GND_net(GND_net), .timer({timer}), .n41296(n41296), .n19(n19_adj_4890), 
            .n34116(n34116), .n34118(n34118), .n34120(n34120), .n34122(n34122), 
            .n34124(n34124), .n34090(n34090), .n34092(n34092), .n34148(n34148), 
            .n34084(n34084), .n34144(n34144), .n34146(n34146), .n34140(n34140), 
            .n34142(n34142), .n34136(n34136), .n34138(n34138), .n34132(n34132), 
            .n34134(n34134), .n34126(n34126), .n34128(n34128), .n34130(n34130), 
            .n34114(n34114), .n34112(n34112), .n34106(n34106), .n34108(n34108), 
            .n34110(n34110), .n34080(n34080), .n34082(n34082), .n34104(n34104), 
            .n34098(n34098), .n34094(n34094), .n34096(n34096), .n41295(n41295), 
            .n41284(n41284), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n41294(n41294), .n41283(n41283), .n41293(n41293), .n41292(n41292), 
            .n4(n4_adj_4906), .start(start), .\state[0] (state[0]), .n106(n106), 
            .\state[1] (state[1]), .n35266(n35266), .n41291(n41291), .n41282(n41282), 
            .n41290(n41290), .n41281(n41281), .n41289(n41289), .n41288(n41288), 
            .n34088(n34088), .n17621(n17621), .n17620(n17620), .n17619(n17619), 
            .n17618(n17618), .n17617(n17617), .n17616(n17616), .n17615(n17615), 
            .n17614(n17614), .n17613(n17613), .n17612(n17612), .n17611(n17611), 
            .n17610(n17610), .n17609(n17609), .n17608(n17608), .n41280(n41280), 
            .PIN_8_c(PIN_8_c), .n36850(n36850), .n41274(n41274), .n41273(n41273), 
            .n17607(n17607), .n41287(n41287), .n17606(n17606), .n17605(n17605), 
            .n17604(n17604), .n17603(n17603), .n41266(n41266), .n11(n11_adj_4891), 
            .n41286(n41286), .n41267(n41267), .n17058(n17058), .n17312(n17312), 
            .n41271(n41271), .n41272(n41272), .n41285(n41285), .n34150(n34150), 
            .n17389(n17389), .n17602(n17602), .n17601(n17601), .n17600(n17600), 
            .n17599(n17599), .n17598(n17598), .n17597(n17597), .n17596(n17596), 
            .n17595(n17595), .n17594(n17594), .n17593(n17593), .n17592(n17592), 
            .n17591(n17591), .n17578(n17578), .n41279(n41279), .n41278(n41278), 
            .n41277(n41277), .n41276(n41276), .\one_wire_N_513[11] (one_wire_N_513[11]), 
            .n41275(n41275), .\one_wire_N_513[8] (one_wire_N_513[8]), .n41270(n41270), 
            .\one_wire_N_513[7] (one_wire_N_513[7]), .\one_wire_N_513[6] (one_wire_N_513[6]), 
            .\one_wire_N_513[5] (one_wire_N_513[5]), .n41269(n41269), .n41268(n41268), 
            .n41297(n41297), .n25771(n25771), .n1138(n1138), .n12(n12_adj_4907), 
            .n8(n8_adj_4341), .\color[20] (color[20]), .\color[4] (color[4]), 
            .\color[10] (color[10]), .\color[11] (color[11]), .\color[9] (color[9]), 
            .\color[17] (color[17]), .\color[18] (color[18]), .\color[19] (color[19]), 
            .\color[1] (color[1]), .\color[2] (color[2]), .\color[3] (color[3]), 
            .\color[12] (color[12]), .\state_3__N_362[1] (state_3__N_362[1]), 
            .n4472(n4472), .n25711(n25711), .n36199(n36199), .n36306(n36306), 
            .n36865(n36865)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(100[10] 106[2])
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31_adj_4414), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n29478), .O(n2622_adj_4484)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_6 (.CI(n29478), .I0(n2555), .I1(GND_net), 
            .CO(n29479));
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n29477), .O(n2623_adj_4483)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1647_3_lut_3_lut (.I0(n2471), .I1(n6089), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1720_5 (.CI(n29477), .I0(n2556), .I1(VCC_net), 
            .CO(n29478));
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n29476), .O(n2624_adj_4482)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_4 (.CI(n29476), .I0(n2557), .I1(VCC_net), 
            .CO(n29477));
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4497), .I2(GND_net), 
            .I3(n29475), .O(n2625_adj_4481)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_3 (.CI(n29475), .I0(n2558_adj_4497), .I1(GND_net), 
            .CO(n29476));
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2658), .I1(VCC_net), 
            .CO(n29475));
    SB_LUT4 rem_4_add_1787_25_lut (.I0(n2669), .I1(n2636_adj_4480), .I2(VCC_net), 
            .I3(n29474), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_24_lut (.I0(GND_net), .I1(n2637_adj_4479), .I2(VCC_net), 
            .I3(n29473), .O(n2704_adj_4453)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_24 (.CI(n29473), .I0(n2637_adj_4479), .I1(VCC_net), 
            .CO(n29474));
    SB_LUT4 rem_4_add_1787_23_lut (.I0(GND_net), .I1(n2638_adj_4478), .I2(VCC_net), 
            .I3(n29472), .O(n2705_adj_4452)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_23 (.CI(n29472), .I0(n2638_adj_4478), .I1(VCC_net), 
            .CO(n29473));
    SB_LUT4 rem_4_add_1787_22_lut (.I0(GND_net), .I1(n2639), .I2(VCC_net), 
            .I3(n29471), .O(n2706_adj_4451)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_22 (.CI(n29471), .I0(n2639), .I1(VCC_net), 
            .CO(n29472));
    SB_LUT4 rem_4_add_1787_21_lut (.I0(GND_net), .I1(n2640), .I2(VCC_net), 
            .I3(n29470), .O(n2707_adj_4450)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_21 (.CI(n29470), .I0(n2640), .I1(VCC_net), 
            .CO(n29471));
    SB_LUT4 rem_4_add_1787_20_lut (.I0(GND_net), .I1(n2641), .I2(VCC_net), 
            .I3(n29469), .O(n2708_adj_4449)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_20 (.CI(n29469), .I0(n2641), .I1(VCC_net), 
            .CO(n29470));
    SB_LUT4 div_46_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1787_19_lut (.I0(GND_net), .I1(n2642_adj_4477), .I2(VCC_net), 
            .I3(n29468), .O(n2709_adj_4448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_19 (.CI(n29468), .I0(n2642_adj_4477), .I1(VCC_net), 
            .CO(n29469));
    SB_LUT4 rem_4_add_1787_18_lut (.I0(GND_net), .I1(n2643_adj_4476), .I2(VCC_net), 
            .I3(n29467), .O(n2710_adj_4447)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1645_3_lut_3_lut (.I0(n2471), .I1(n6087), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n89), .I1(n15986), .I2(GND_net), .I3(GND_net), 
            .O(n15983));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1648_3_lut_3_lut (.I0(n2471), .I1(n6090), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13086_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13293), .I3(GND_net), .O(n17831));   // verilog/coms.v(126[12] 289[6])
    defparam i13086_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF color__i9 (.Q(color[9]), .C(LED_c), .D(n18122));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i10 (.Q(color[10]), .C(LED_c), .D(n18123));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i11 (.Q(color[11]), .C(LED_c), .D(n18124));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i12 (.Q(color[12]), .C(LED_c), .D(n18125));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i17 (.Q(color[17]), .C(LED_c), .D(n36325));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i18 (.Q(color[18]), .C(LED_c), .D(n32676));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i19 (.Q(color[19]), .C(LED_c), .D(n32678));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i2 (.Q(color[2]), .C(LED_c), .D(n32658));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i20 (.Q(color[20]), .C(LED_c), .D(n32680));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i3 (.Q(color[3]), .C(LED_c), .D(n32660));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i4 (.Q(color[4]), .C(LED_c), .D(n32662));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_DFF color__i1 (.Q(color[1]), .C(LED_c), .D(n36299));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_LUT4 i13087_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13293), .I3(GND_net), .O(n17832));   // verilog/coms.v(126[12] 289[6])
    defparam i13087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1661_3_lut_3_lut (.I0(n2471), .I1(n6103), .I2(n528), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13088_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13293), .I3(GND_net), .O(n17833));   // verilog/coms.v(126[12] 289[6])
    defparam i13088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1646_3_lut_3_lut (.I0(n2471), .I1(n6088), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1598 (.I0(n92), .I1(n15946), .I2(GND_net), .I3(GND_net), 
            .O(n15980));
    defparam i1_2_lut_adj_1598.LUT_INIT = 16'hdddd;
    SB_LUT4 rem_4_i1803_3_lut (.I0(n2650), .I1(n2717_adj_4440), .I2(n2669), 
            .I3(GND_net), .O(n2749));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1797_3_lut (.I0(n2644), .I1(n2711_adj_4446), .I2(n2669), 
            .I3(GND_net), .O(n2743));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1804_3_lut (.I0(n2651), .I1(n2718_adj_4439), .I2(n2669), 
            .I3(GND_net), .O(n2750));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1806_3_lut (.I0(n2653), .I1(n2720_adj_4437), .I2(n2669), 
            .I3(GND_net), .O(n2752));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i1802_3_lut (.I0(n2649), .I1(n2716_adj_4441), .I2(n2669), 
            .I3(GND_net), .O(n2748));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1807_3_lut (.I0(n2654), .I1(n2721), .I2(n2669), .I3(GND_net), 
            .O(n2753));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1792_3_lut (.I0(n2639), .I1(n2706_adj_4451), .I2(n2669), 
            .I3(GND_net), .O(n2738));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1791_3_lut (.I0(n2638_adj_4478), .I1(n2705_adj_4452), 
            .I2(n2669), .I3(GND_net), .O(n2737));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1650_3_lut_3_lut (.I0(n2471), .I1(n6092), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1790_3_lut (.I0(n2637_adj_4479), .I1(n2704_adj_4453), 
            .I2(n2669), .I3(GND_net), .O(n2736));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1799_3_lut (.I0(n2646), .I1(n2713_adj_4444), .I2(n2669), 
            .I3(GND_net), .O(n2745));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1794_3_lut (.I0(n2641), .I1(n2708_adj_4449), .I2(n2669), 
            .I3(GND_net), .O(n2740));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1795_3_lut (.I0(n2642_adj_4477), .I1(n2709_adj_4448), 
            .I2(n2669), .I3(GND_net), .O(n2741));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1793_3_lut (.I0(n2640), .I1(n2707_adj_4450), .I2(n2669), 
            .I3(GND_net), .O(n2739));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1809_3_lut (.I0(n2656), .I1(n2723_adj_4436), .I2(n2669), 
            .I3(GND_net), .O(n2755));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1808_3_lut (.I0(n2655), .I1(n2722), .I2(n2669), .I3(GND_net), 
            .O(n2754));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1796_3_lut (.I0(n2643_adj_4476), .I1(n2710_adj_4447), 
            .I2(n2669), .I3(GND_net), .O(n2742));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1801_3_lut (.I0(n2648), .I1(n2715_adj_4442), .I2(n2669), 
            .I3(GND_net), .O(n2747));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1800_3_lut (.I0(n2647), .I1(n2714_adj_4443), .I2(n2669), 
            .I3(GND_net), .O(n2746));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1651_3_lut_3_lut (.I0(n2471), .I1(n6093), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1805_3_lut (.I0(n2652), .I1(n2719_adj_4438), .I2(n2669), 
            .I3(GND_net), .O(n2751));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i1798_3_lut (.I0(n2645), .I1(n2712_adj_4445), .I2(n2669), 
            .I3(GND_net), .O(n2744));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1656_3_lut_3_lut (.I0(n2471), .I1(n6098), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1811_3_lut (.I0(n2658), .I1(n2725), .I2(n2669), .I3(GND_net), 
            .O(n2757));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1810_3_lut (.I0(n2657), .I1(n2724_adj_4435), .I2(n2669), 
            .I3(GND_net), .O(n2756));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n36500));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut (.I0(n2744), .I1(n2751), .I2(n2746), .I3(n2747), 
            .O(n34_adj_4869));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1599 (.I0(n95), .I1(n15940), .I2(GND_net), .I3(GND_net), 
            .O(n15937));
    defparam i1_2_lut_adj_1599.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(n2742), .I1(n2754), .I2(n36500), .I3(n2755), 
            .O(n25_adj_4876));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut (.I0(n2739), .I1(n2741), .I2(n2740), .I3(n2745), 
            .O(n32_adj_4870));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1653_3_lut_3_lut (.I0(n2471), .I1(n6095), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11_4_lut (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31_adj_4871));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2753), .I1(n2748), .I2(n2752), .I3(n2750), 
            .O(n35_adj_4819));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n25_adj_4876), .I1(n34_adj_4869), .I2(n2743), 
            .I3(n2749), .O(n37_adj_4772));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37_adj_4772), .I1(n35_adj_4819), .I2(n31_adj_4871), 
            .I3(n32_adj_4870), .O(n2768));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4418), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1600 (.I0(n98), .I1(n15977), .I2(GND_net), .I3(GND_net), 
            .O(n15930));
    defparam i1_2_lut_adj_1600.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13089_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13293), .I3(GND_net), .O(n17834));   // verilog/coms.v(126[12] 289[6])
    defparam i13089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15930), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 div_46_i1652_3_lut_3_lut (.I0(n2471), .I1(n6094), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37376_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n44228));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i37376_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1660_3_lut_3_lut (.I0(n2471), .I1(n6102), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13084_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13293), .I3(GND_net), .O(n17829));   // verilog/coms.v(126[12] 289[6])
    defparam i13084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(n2254), .I1(n2246), .I2(n36545), .I3(n2255), 
            .O(n19_adj_4913));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_i1659_3_lut_3_lut (.I0(n2471), .I1(n6101), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1787_18 (.CI(n29467), .I0(n2643_adj_4476), .I1(VCC_net), 
            .CO(n29468));
    SB_LUT4 rem_4_add_1787_17_lut (.I0(GND_net), .I1(n2644), .I2(VCC_net), 
            .I3(n29466), .O(n2711_adj_4446)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1658_3_lut_3_lut (.I0(n2471), .I1(n6100), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546_adj_4505), .I1(n2613), .I2(n2570), 
            .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4939));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1657_3_lut_3_lut (.I0(n2471), .I1(n6099), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4527));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544_adj_4507), .I1(n2611), .I2(n2570), 
            .I3(GND_net), .O(n2643_adj_4476));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13216_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n35433), .I3(GND_net), .O(n17961));   // verilog/coms.v(126[12] 289[6])
    defparam i13216_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1787_17 (.CI(n29466), .I0(n2644), .I1(VCC_net), 
            .CO(n29467));
    SB_LUT4 i13229_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n35435), .I3(GND_net), .O(n17974));   // verilog/coms.v(126[12] 289[6])
    defparam i13229_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3459));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13090_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13293), .I3(GND_net), .O(n17835));   // verilog/coms.v(126[12] 289[6])
    defparam i13090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1649_3_lut_3_lut (.I0(n2471), .I1(n6091), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1654_3_lut_3_lut (.I0(n2471), .I1(n6096), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1714_3_lut_3_lut (.I0(n2558), .I1(n6121), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13091_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13293), .I3(GND_net), .O(n17836));   // verilog/coms.v(126[12] 289[6])
    defparam i13091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1601 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4914));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i1_2_lut_adj_1601.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_4912));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n19_adj_4913), .I1(n26_adj_4910), .I2(n2247), 
            .I3(n2250), .O(n28_adj_4909));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1699_3_lut_3_lut (.I0(n2558), .I1(n6106), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1701_3_lut_3_lut (.I0(n2558), .I1(n6108), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543_adj_4508), .I1(n2610), .I2(n2570), 
            .I3(GND_net), .O(n2642_adj_4477));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_31_lut (.I0(n3263), .I1(n3230), .I2(VCC_net), 
            .I3(n29211), .O(n38986)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_16_lut (.I0(GND_net), .I1(n2645), .I2(VCC_net), 
            .I3(n29465), .O(n2712_adj_4445)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_16 (.CI(n29465), .I0(n2645), .I1(VCC_net), 
            .CO(n29466));
    SB_LUT4 rem_4_add_1787_15_lut (.I0(GND_net), .I1(n2646), .I2(VCC_net), 
            .I3(n29464), .O(n2713_adj_4444)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_15 (.CI(n29464), .I0(n2646), .I1(VCC_net), 
            .CO(n29465));
    SB_LUT4 div_46_i1702_3_lut_3_lut (.I0(n2558), .I1(n6109), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32_adj_4413), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1787_14_lut (.I0(GND_net), .I1(n2647), .I2(VCC_net), 
            .I3(n29463), .O(n2714_adj_4443)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_30_lut (.I0(GND_net), .I1(n3231), .I2(VCC_net), 
            .I3(n29210), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_30 (.CI(n29210), .I0(n3231), .I1(VCC_net), 
            .CO(n29211));
    SB_LUT4 rem_4_add_2189_29_lut (.I0(GND_net), .I1(n3232), .I2(VCC_net), 
            .I3(n29209), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_29 (.CI(n29209), .I0(n3232), .I1(VCC_net), 
            .CO(n29210));
    SB_CARRY rem_4_add_1787_14 (.CI(n29463), .I0(n2647), .I1(VCC_net), 
            .CO(n29464));
    SB_LUT4 rem_4_add_1787_13_lut (.I0(GND_net), .I1(n2648), .I2(VCC_net), 
            .I3(n29462), .O(n2715_adj_4442)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(209[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1787_13 (.CI(n29462), .I0(n2648), .I1(VCC_net), 
            .CO(n29463));
    SB_LUT4 rem_4_add_2189_28_lut (.I0(GND_net), .I1(n3233), .I2(VCC_net), 
            .I3(n29208), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1602 (.I0(n2251), .I1(n28_adj_4909), .I2(n24_adj_4912), 
            .I3(n16_adj_4914), .O(n2273_adj_4581));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1787_12_lut (.I0(GND_net), .I1(n2649), .I2(VCC_net), 
            .I3(n29461), .O(n2716_adj_4441)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_12 (.CI(n29461), .I0(n2649), .I1(VCC_net), 
            .CO(n29462));
    SB_CARRY rem_4_add_2189_28 (.CI(n29208), .I0(n3233), .I1(VCC_net), 
            .CO(n29209));
    SB_LUT4 rem_4_add_1787_11_lut (.I0(GND_net), .I1(n2650), .I2(VCC_net), 
            .I3(n29460), .O(n2717_adj_4440)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_27_lut (.I0(GND_net), .I1(n3234), .I2(VCC_net), 
            .I3(n29207), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_27 (.CI(n29207), .I0(n3234), .I1(VCC_net), 
            .CO(n29208));
    SB_LUT4 rem_4_add_2189_26_lut (.I0(GND_net), .I1(n3235), .I2(VCC_net), 
            .I3(n29206), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n29460), .I0(n2650), .I1(VCC_net), 
            .CO(n29461));
    SB_CARRY rem_4_add_2189_26 (.CI(n29206), .I0(n3235), .I1(VCC_net), 
            .CO(n29207));
    SB_LUT4 rem_4_add_1787_10_lut (.I0(GND_net), .I1(n2651), .I2(VCC_net), 
            .I3(n29459), .O(n2718_adj_4439)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1700_3_lut_3_lut (.I0(n2558), .I1(n6107), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_25_lut (.I0(GND_net), .I1(n3236), .I2(VCC_net), 
            .I3(n29205), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_10 (.CI(n29459), .I0(n2651), .I1(VCC_net), 
            .CO(n29460));
    SB_LUT4 div_46_i1705_3_lut_3_lut (.I0(n2558), .I1(n6112), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1787_9_lut (.I0(GND_net), .I1(n2652), .I2(VCC_net), 
            .I3(n29458), .O(n2719_adj_4438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_25 (.CI(n29205), .I0(n3236), .I1(VCC_net), 
            .CO(n29206));
    SB_CARRY rem_4_add_1787_9 (.CI(n29458), .I0(n2652), .I1(VCC_net), 
            .CO(n29459));
    SB_LUT4 rem_4_add_1787_8_lut (.I0(GND_net), .I1(n2653), .I2(VCC_net), 
            .I3(n29457), .O(n2720_adj_4437)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_8 (.CI(n29457), .I0(n2653), .I1(VCC_net), 
            .CO(n29458));
    SB_LUT4 rem_4_add_1787_7_lut (.I0(GND_net), .I1(n2654), .I2(GND_net), 
            .I3(n29456), .O(n2721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_24_lut (.I0(GND_net), .I1(n3237), .I2(VCC_net), 
            .I3(n29204), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_24 (.CI(n29204), .I0(n3237), .I1(VCC_net), 
            .CO(n29205));
    SB_LUT4 div_46_i1703_3_lut_3_lut (.I0(n2558), .I1(n6110), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i5_4_lut_adj_1603 (.I0(n36444), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_4901));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_2189_23_lut (.I0(GND_net), .I1(n3238), .I2(VCC_net), 
            .I3(n29203), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1706_3_lut_3_lut (.I0(n2558), .I1(n6113), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut (.I0(n1453), .I1(n12_adj_4901), .I2(n1449), .I3(n1448), 
            .O(n1481));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417_adj_4493), .I2(n1382), 
            .I3(GND_net), .O(n1449));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2189_23 (.CI(n29203), .I0(n3238), .I1(VCC_net), 
            .CO(n29204));
    SB_CARRY rem_4_add_1787_7 (.CI(n29456), .I0(n2654), .I1(GND_net), 
            .CO(n29457));
    SB_LUT4 rem_4_add_1787_6_lut (.I0(GND_net), .I1(n2655), .I2(GND_net), 
            .I3(n29455), .O(n2722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_6 (.CI(n29455), .I0(n2655), .I1(GND_net), 
            .CO(n29456));
    SB_LUT4 rem_4_add_2189_22_lut (.I0(GND_net), .I1(n3239), .I2(VCC_net), 
            .I3(n29202), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_22 (.CI(n29202), .I0(n3239), .I1(VCC_net), 
            .CO(n29203));
    SB_LUT4 rem_4_add_1787_5_lut (.I0(GND_net), .I1(n2656), .I2(VCC_net), 
            .I3(n29454), .O(n2723_adj_4436)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_21_lut (.I0(GND_net), .I1(n3240), .I2(VCC_net), 
            .I3(n29201), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i37332_1_lut (.I0(n3457), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44186));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37332_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545_adj_4506), .I1(n2612), .I2(n2570), 
            .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2287_3_lut (.I0(n3358), .I1(n10223), .I2(n3362), .I3(GND_net), 
            .O(n3457));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2189_21 (.CI(n29201), .I0(n3240), .I1(VCC_net), 
            .CO(n29202));
    SB_LUT4 i1_3_lut_adj_1604 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n36441));
    defparam i1_3_lut_adj_1604.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_2189_20_lut (.I0(GND_net), .I1(n3241), .I2(VCC_net), 
            .I3(n29200), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_20 (.CI(n29200), .I0(n3241), .I1(VCC_net), 
            .CO(n29201));
    SB_LUT4 rem_4_add_2189_19_lut (.I0(GND_net), .I1(n3242), .I2(VCC_net), 
            .I3(n29199), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_19 (.CI(n29199), .I0(n3242), .I1(VCC_net), 
            .CO(n29200));
    SB_LUT4 rem_4_add_2189_18_lut (.I0(GND_net), .I1(n3243), .I2(VCC_net), 
            .I3(n29198), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut (.I0(n1554_adj_4488), .I1(n1551), .I2(n36441), .I3(n1555), 
            .O(n11_adj_4899));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i3_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_i1719_3_lut_3_lut (.I0(n2558), .I1(n6126), .I2(n529), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1787_5 (.CI(n29454), .I0(n2656), .I1(VCC_net), 
            .CO(n29455));
    SB_CARRY rem_4_add_2189_18 (.CI(n29198), .I0(n3243), .I1(VCC_net), 
            .CO(n29199));
    SB_LUT4 rem_4_add_1787_4_lut (.I0(GND_net), .I1(n2657), .I2(VCC_net), 
            .I3(n29453), .O(n2724_adj_4435)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_17_lut (.I0(GND_net), .I1(n3244), .I2(VCC_net), 
            .I3(n29197), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1704_3_lut_3_lut (.I0(n2558), .I1(n6111), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1787_4 (.CI(n29453), .I0(n2657), .I1(VCC_net), 
            .CO(n29454));
    SB_LUT4 rem_4_add_1787_3_lut (.I0(GND_net), .I1(n2658), .I2(GND_net), 
            .I3(n29452), .O(n2725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_3 (.CI(n29452), .I0(n2658), .I1(GND_net), 
            .CO(n29453));
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2758), .I1(VCC_net), 
            .CO(n29452));
    SB_CARRY rem_4_add_2189_17 (.CI(n29197), .I0(n3244), .I1(VCC_net), 
            .CO(n29198));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n29451), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4420), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558_adj_4497));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1709_3_lut_3_lut (.I0(n2558), .I1(n6116), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n29450), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut_adj_1605 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_4898));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_2189_16_lut (.I0(GND_net), .I1(n3245), .I2(VCC_net), 
            .I3(n29196), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_16 (.CI(n29196), .I0(n3245), .I1(VCC_net), 
            .CO(n29197));
    SB_CARRY rem_4_add_1854_25 (.CI(n29450), .I0(n2736), .I1(VCC_net), 
            .CO(n29451));
    SB_LUT4 i13210_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n35433), .I3(GND_net), .O(n17955));   // verilog/coms.v(126[12] 289[6])
    defparam i13210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1606 (.I0(n2356), .I1(n2358_adj_4578), .I2(GND_net), 
            .I3(GND_net), .O(n38713));
    defparam i1_2_lut_adj_1606.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_add_2189_15_lut (.I0(GND_net), .I1(n3246), .I2(VCC_net), 
            .I3(n29195), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n29449), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_15 (.CI(n29195), .I0(n3246), .I1(VCC_net), 
            .CO(n29196));
    SB_LUT4 rem_4_add_2189_14_lut (.I0(GND_net), .I1(n3247), .I2(VCC_net), 
            .I3(n29194), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_24 (.CI(n29449), .I0(n2737), .I1(VCC_net), 
            .CO(n29450));
    SB_CARRY rem_4_add_2189_14 (.CI(n29194), .I0(n3247), .I1(VCC_net), 
            .CO(n29195));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(GND_net), .I1(n3248), .I2(VCC_net), 
            .I3(n29193), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_13 (.CI(n29193), .I0(n3248), .I1(VCC_net), 
            .CO(n29194));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(GND_net), .I1(n3249), .I2(VCC_net), 
            .I3(n29192), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_12 (.CI(n29192), .I0(n3249), .I1(VCC_net), 
            .CO(n29193));
    SB_LUT4 rem_4_add_2189_11_lut (.I0(GND_net), .I1(n3250), .I2(VCC_net), 
            .I3(n29191), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1675_3_lut (.I0(n2458_adj_4516), .I1(n2525), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2557));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4938));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2189_11 (.CI(n29191), .I0(n3250), .I1(VCC_net), 
            .CO(n29192));
    SB_LUT4 rem_4_add_2189_10_lut (.I0(GND_net), .I1(n3251), .I2(VCC_net), 
            .I3(n29190), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_10 (.CI(n29190), .I0(n3251), .I1(VCC_net), 
            .CO(n29191));
    SB_LUT4 i1_4_lut (.I0(n2354), .I1(n38713), .I2(n2355), .I3(n2357_adj_4579), 
            .O(n36482));
    defparam i1_4_lut.LUT_INIT = 16'ha080;
    SB_LUT4 i13211_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n35433), .I3(GND_net), .O(n17956));   // verilog/coms.v(126[12] 289[6])
    defparam i13211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_9_lut (.I0(GND_net), .I1(n3252), .I2(VCC_net), 
            .I3(n29189), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_9 (.CI(n29189), .I0(n3252), .I1(VCC_net), 
            .CO(n29190));
    SB_LUT4 div_46_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4526));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2189_8_lut (.I0(GND_net), .I1(n3253), .I2(VCC_net), 
            .I3(n29188), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_8 (.CI(n29188), .I0(n3253), .I1(VCC_net), 
            .CO(n29189));
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n29448), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_7_lut (.I0(GND_net), .I1(n3254), .I2(GND_net), 
            .I3(n29187), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_7 (.CI(n29187), .I0(n3254), .I1(GND_net), 
            .CO(n29188));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(GND_net), .I1(n3255), .I2(GND_net), 
            .I3(n29186), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_23 (.CI(n29448), .I0(n2738), .I1(VCC_net), 
            .CO(n29449));
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n29447), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_22 (.CI(n29447), .I0(n2739), .I1(VCC_net), 
            .CO(n29448));
    SB_CARRY rem_4_add_2189_6 (.CI(n29186), .I0(n3255), .I1(GND_net), 
            .CO(n29187));
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649_adj_4465), .I1(n1716), .I2(n1679), 
            .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4937));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4525));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n29446), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648_adj_4464), .I1(n1715), .I2(n1679), 
            .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_5_lut (.I0(GND_net), .I1(n3256), .I2(VCC_net), 
            .I3(n29185), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_5 (.CI(n29185), .I0(n3256), .I1(VCC_net), 
            .CO(n29186));
    SB_LUT4 rem_4_add_2189_4_lut (.I0(GND_net), .I1(n3257), .I2(VCC_net), 
            .I3(n29184), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_4 (.CI(n29184), .I0(n3257), .I1(VCC_net), 
            .CO(n29185));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(GND_net), .I1(n3258), .I2(GND_net), 
            .I3(n29183), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4524));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2189_3 (.CI(n29183), .I0(n3258), .I1(GND_net), 
            .CO(n29184));
    SB_CARRY rem_4_add_1854_21 (.CI(n29446), .I0(n2740), .I1(VCC_net), 
            .CO(n29447));
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n29445), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_20 (.CI(n29445), .I0(n2741), .I1(VCC_net), 
            .CO(n29446));
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3358), .I1(VCC_net), 
            .CO(n29183));
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n29444), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(n13_adj_4898), .I1(n11_adj_4899), .I2(n1553_adj_4487), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1854_19 (.CI(n29444), .I0(n2742), .I1(VCC_net), 
            .CO(n29445));
    SB_LUT4 communication_counter_1199_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n29182), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1199_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n29181), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_32 (.CI(n29181), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n29182));
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n29443), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4523));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 communication_counter_1199_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n29180), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_55 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 div_46_i1708_3_lut_3_lut (.I0(n2558), .I1(n6115), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY communication_counter_1199_add_4_31 (.CI(n29180), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n29181));
    SB_LUT4 communication_counter_1199_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n29179), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_30 (.CI(n29179), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n29180));
    SB_LUT4 communication_counter_1199_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n29178), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4428), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758_adj_4458));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_29 (.CI(n29178), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n29179));
    SB_LUT4 communication_counter_1199_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n29177), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4522));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4936));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4521));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37329_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44183));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37329_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n10222), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY communication_counter_1199_add_4_28 (.CI(n29177), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n29178));
    SB_CARRY rem_4_add_1854_18 (.CI(n29443), .I0(n2743), .I1(VCC_net), 
            .CO(n29444));
    SB_LUT4 communication_counter_1199_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n29176), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_27 (.CI(n29176), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n29177));
    SB_LUT4 communication_counter_1199_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n29175), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_26 (.CI(n29175), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n29176));
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n29442), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1199_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n29174), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_25 (.CI(n29174), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n29175));
    SB_LUT4 communication_counter_1199_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n29173), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_24 (.CI(n29173), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n29174));
    SB_LUT4 communication_counter_1199_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n29172), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4520));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13085_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13293), .I3(GND_net), .O(n17830));   // verilog/coms.v(126[12] 289[6])
    defparam i13085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1062_rep_69_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), 
            .I3(GND_net), .O(n1656));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1062_rep_69_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1854_17 (.CI(n29442), .I0(n2744), .I1(VCC_net), 
            .CO(n29443));
    SB_LUT4 div_46_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4519));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37326_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44180));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37326_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n29441), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_23 (.CI(n29172), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n29173));
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164), .I3(GND_net), 
            .O(n3235));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4566));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4935));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4565));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n10221), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1717_3_lut_3_lut (.I0(n2558), .I1(n6124), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1199_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n29171), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164), .I3(GND_net), 
            .O(n3233));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1718_3_lut_3_lut (.I0(n2558), .I1(n6125), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1199_add_4_22 (.CI(n29171), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n29172));
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164), .I3(GND_net), 
            .O(n3234));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n29170), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_21 (.CI(n29170), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n29171));
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164), .I3(GND_net), 
            .O(n3232));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF communication_counter_1199__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4318));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4934));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1854_16 (.CI(n29441), .I0(n2745), .I1(VCC_net), 
            .CO(n29442));
    SB_LUT4 i37323_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44177));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37323_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1199_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n29169), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_20 (.CI(n29169), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n29170));
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n29440), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_15 (.CI(n29440), .I0(n2746), .I1(VCC_net), 
            .CO(n29441));
    SB_LUT4 communication_counter_1199_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n29168), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_19 (.CI(n29168), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n29169));
    SB_LUT4 communication_counter_1199_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n29167), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_18 (.CI(n29167), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n29168));
    SB_LUT4 add_577_24_lut (.I0(duty[22]), .I1(n44224), .I2(n3), .I3(n28683), 
            .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n29439), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_14 (.CI(n29439), .I0(n2747), .I1(VCC_net), 
            .CO(n29440));
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214), .I2(n3164), .I3(GND_net), 
            .O(n3246));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_577_23_lut (.I0(duty[21]), .I1(n44224), .I2(n4), .I3(n28682), 
            .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n10220), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_577_23 (.CI(n28682), .I0(n44224), .I1(n4), .CO(n28683));
    SB_LUT4 add_577_22_lut (.I0(duty[20]), .I1(n44224), .I2(n5), .I3(n28681), 
            .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_577_22 (.CI(n28681), .I0(n44224), .I1(n5), .CO(n28682));
    SB_LUT4 add_577_21_lut (.I0(duty[19]), .I1(n44224), .I2(n6_adj_4314), 
            .I3(n28680), .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213), .I2(n3164), .I3(GND_net), 
            .O(n3245));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n29166), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_21 (.CI(n28680), .I0(n44224), .I1(n6_adj_4314), .CO(n28681));
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n29438), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_577_20_lut (.I0(duty[18]), .I1(n44224), .I2(n7_adj_4315), 
            .I3(n28679), .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_577_20 (.CI(n28679), .I0(n44224), .I1(n7_adj_4315), .CO(n28680));
    SB_CARRY rem_4_add_1854_13 (.CI(n29438), .I0(n2748), .I1(VCC_net), 
            .CO(n29439));
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210), .I2(n3164), .I3(GND_net), 
            .O(n3242));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4564));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n29437), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_12 (.CI(n29437), .I0(n2749), .I1(VCC_net), 
            .CO(n29438));
    SB_LUT4 add_577_19_lut (.I0(duty[17]), .I1(n44224), .I2(n8_adj_4316), 
            .I3(n28678), .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_1199_add_4_17 (.CI(n29166), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n29167));
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209), .I2(n3164), .I3(GND_net), 
            .O(n3241));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1058_3_lut (.I0(n1553_adj_4487), .I1(n1620), .I2(n1580), 
            .I3(GND_net), .O(n1652_adj_4459));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n29436), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_11 (.CI(n29436), .I0(n2750), .I1(VCC_net), 
            .CO(n29437));
    SB_CARRY add_577_19 (.CI(n28678), .I0(n44224), .I1(n8_adj_4316), .CO(n28679));
    SB_LUT4 i13227_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n35435), .I3(GND_net), .O(n17972));   // verilog/coms.v(126[12] 289[6])
    defparam i13227_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4563));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1199_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n29165), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164), .I3(GND_net), 
            .O(n3239));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1712_3_lut_3_lut (.I0(n2558), .I1(n6119), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164), .I3(GND_net), 
            .O(n3237));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4933));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37320_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44174));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37320_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n10219), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164), .I3(GND_net), 
            .O(n3238));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4562));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649_adj_4465));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13190_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n35428), .I3(GND_net), .O(n17935));   // verilog/coms.v(126[12] 289[6])
    defparam i13190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164), .I3(GND_net), 
            .O(n3236));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n29435), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2215_3_lut (.I0(n3254), .I1(n3321), .I2(n3263), .I3(GND_net), 
            .O(n3353));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2217_3_lut (.I0(n3256), .I1(n3323), .I2(n3263), .I3(GND_net), 
            .O(n3355));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648_adj_4464));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4932));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4931));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_1199_add_4_16 (.CI(n29165), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n29166));
    SB_LUT4 communication_counter_1199_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n29164), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_15 (.CI(n29164), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n29165));
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4930));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2138_3_lut (.I0(n3145), .I1(n3212), .I2(n3164), .I3(GND_net), 
            .O(n3244));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2143_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2216_3_lut (.I0(n3255), .I1(n3322), .I2(n3263), .I3(GND_net), 
            .O(n3354));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4323));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4561));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2144_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4429), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164), .I3(GND_net), 
            .O(n3231));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4560));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211), .I2(n3164), .I3(GND_net), 
            .O(n3243));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2219_3_lut (.I0(n3258), .I1(n3325), .I2(n3263), .I3(GND_net), 
            .O(n3357));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_10 (.CI(n29435), .I0(n2751), .I1(VCC_net), 
            .CO(n29436));
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n29434), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2142_3_lut (.I0(n3149), .I1(n3216), .I2(n3164), .I3(GND_net), 
            .O(n3248));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2218_3_lut (.I0(n3257), .I1(n3324), .I2(n3263), .I3(GND_net), 
            .O(n3356));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2206_3_lut (.I0(n3245), .I1(n3312), .I2(n3263), .I3(GND_net), 
            .O(n3344));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2208_3_lut (.I0(n3247), .I1(n3314), .I2(n3263), .I3(GND_net), 
            .O(n3346));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2213_3_lut (.I0(n3252), .I1(n3319), .I2(n3263), .I3(GND_net), 
            .O(n3351));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4929));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215), .I2(n3164), .I3(GND_net), 
            .O(n3247));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1734_3_lut (.I0(n2549_adj_4502), .I1(n2616), .I2(n2570), 
            .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221), .I2(n3164), .I3(GND_net), 
            .O(n3253));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220), .I2(n3164), .I3(GND_net), 
            .O(n3252));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i994_rep_71_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), 
            .I3(GND_net), .O(n1556));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i994_rep_71_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223), .I2(n3164), .I3(GND_net), 
            .O(n3255));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4322));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222), .I2(n3164), .I3(GND_net), 
            .O(n3254));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164), .I3(GND_net), 
            .O(n3240));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2077_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2077_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_9 (.CI(n29434), .I0(n2752), .I1(VCC_net), 
            .CO(n29435));
    SB_LUT4 communication_counter_1199_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n29163), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_14 (.CI(n29163), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n29164));
    SB_LUT4 communication_counter_1199_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n29162), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n3249), .I1(n3351), .I2(n3316), .I3(n3263), 
            .O(n38613));
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'hfcee;
    SB_CARRY communication_counter_1199_add_4_13 (.CI(n29162), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n29163));
    SB_LUT4 div_46_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4559));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1199_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n29161), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_12 (.CI(n29161), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n29162));
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n29160), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n38613), .I1(n3251), .I2(n3318), .I3(n3263), 
            .O(n38615));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'hfaee;
    SB_LUT4 div_46_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4558));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n29433), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2071_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_8 (.CI(n29433), .I0(n2753), .I1(VCC_net), 
            .CO(n29434));
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4928));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n29432), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_11 (.CI(n29160), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n29161));
    SB_LUT4 communication_counter_1199_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n29159), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_10 (.CI(n29159), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n29160));
    SB_LUT4 rem_4_i2058_rep_78_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), 
            .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2058_rep_78_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n29158), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13212_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n35433), .I3(GND_net), .O(n17957));   // verilog/coms.v(126[12] 289[6])
    defparam i13212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12879_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17624));   // verilog/coms.v(126[12] 289[6])
    defparam i12879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12880_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17625));   // verilog/coms.v(126[12] 289[6])
    defparam i12880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(n3242), .I1(n38615), .I2(n3309), .I3(n3263), 
            .O(n38617));
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_9 (.CI(n29158), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n29159));
    SB_LUT4 i1_4_lut_adj_1610 (.I0(n3240), .I1(n38617), .I2(n3307), .I3(n3263), 
            .O(n38619));
    defparam i1_4_lut_adj_1610.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n29157), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_8 (.CI(n29157), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n29158));
    SB_LUT4 communication_counter_1199_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n29156), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2075_3_lut (.I0(n3050), .I1(n3117), .I2(n3065), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_7 (.CI(n29156), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n29157));
    SB_LUT4 i12881_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17626));   // verilog/coms.v(126[12] 289[6])
    defparam i12881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2076_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1611 (.I0(n3239), .I1(n38619), .I2(n3306), .I3(n3263), 
            .O(n38621));
    defparam i1_4_lut_adj_1611.LUT_INIT = 16'hfcee;
    SB_LUT4 communication_counter_1199_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n29155), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12882_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17627));   // verilog/coms.v(126[12] 289[6])
    defparam i12882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554_adj_4488));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_6 (.CI(n29155), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n29156));
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2207_3_lut (.I0(n3246), .I1(n3313), .I2(n3263), .I3(GND_net), 
            .O(n3345));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(n3253), .I1(n3344), .I2(n3320), .I3(n3263), 
            .O(n38551));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'hfcee;
    SB_LUT4 i12883_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17628));   // verilog/coms.v(126[12] 289[6])
    defparam i12883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12884_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17629));   // verilog/coms.v(126[12] 289[6])
    defparam i12884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2204_3_lut (.I0(n3243), .I1(n3310), .I2(n3263), .I3(GND_net), 
            .O(n3342));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12885_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17630));   // verilog/coms.v(126[12] 289[6])
    defparam i12885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2205_3_lut (.I0(n3244), .I1(n3311), .I2(n3263), .I3(GND_net), 
            .O(n3343));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1613 (.I0(n3356), .I1(n3357), .I2(n3358), .I3(GND_net), 
            .O(n36533));
    defparam i1_3_lut_adj_1613.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(n3343), .I1(n3342), .I2(n38551), .I3(n3345), 
            .O(n38557));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i12886_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17631));   // verilog/coms.v(126[12] 289[6])
    defparam i12886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12887_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17632));   // verilog/coms.v(126[12] 289[6])
    defparam i12887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12888_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17633));   // verilog/coms.v(126[12] 289[6])
    defparam i12888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(n3354), .I1(n38557), .I2(n36533), .I3(n3355), 
            .O(n38559));
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n3241), .I1(n38559), .I2(n3308), .I3(n3263), 
            .O(n38561));
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i991_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), .I3(GND_net), 
            .O(n1553_adj_4487));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(n3237), .I1(n38561), .I2(n3304), .I3(n3263), 
            .O(n38563));
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1618 (.I0(n3236), .I1(n38621), .I2(n3303), .I3(n3263), 
            .O(n38623));
    defparam i1_4_lut_adj_1618.LUT_INIT = 16'hfcee;
    SB_LUT4 div_46_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4557));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12889_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17634));   // verilog/coms.v(126[12] 289[6])
    defparam i12889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1619 (.I0(n3353), .I1(n3250), .I2(n3317), .I3(n3263), 
            .O(n38651));
    defparam i1_4_lut_adj_1619.LUT_INIT = 16'hfaee;
    SB_LUT4 i12890_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17635));   // verilog/coms.v(126[12] 289[6])
    defparam i12890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_7 (.CI(n29432), .I0(n2754), .I1(GND_net), 
            .CO(n29433));
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n29431), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12891_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17636));   // verilog/coms.v(126[12] 289[6])
    defparam i12891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1620 (.I0(n3248), .I1(n3346), .I2(n3315), .I3(n3263), 
            .O(n28));
    defparam i3_4_lut_adj_1620.LUT_INIT = 16'hfcee;
    SB_LUT4 i12892_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17637));   // verilog/coms.v(126[12] 289[6])
    defparam i12892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_6 (.CI(n29431), .I0(n2755), .I1(GND_net), 
            .CO(n29432));
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n29430), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2069_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), .I3(GND_net), 
            .O(n3143));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12893_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17638));   // verilog/coms.v(126[12] 289[6])
    defparam i12893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_5 (.CI(n29430), .I0(n2756), .I1(VCC_net), 
            .CO(n29431));
    SB_LUT4 i12894_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17639));   // verilog/coms.v(126[12] 289[6])
    defparam i12894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n29154), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n29429), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_4 (.CI(n29429), .I0(n2757), .I1(VCC_net), 
            .CO(n29430));
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n29428), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(n38623), .I1(n3235), .I2(n3302), .I3(n3263), 
            .O(n46));
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'hfaee;
    SB_LUT4 i12895_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17640));   // verilog/coms.v(126[12] 289[6])
    defparam i12895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12896_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17641));   // verilog/coms.v(126[12] 289[6])
    defparam i12896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_3 (.CI(n29428), .I0(n2758), .I1(GND_net), 
            .CO(n29429));
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1622 (.I0(n38563), .I1(n3233), .I2(n3300), .I3(n3263), 
            .O(n47));
    defparam i1_4_lut_adj_1622.LUT_INIT = 16'hfaee;
    SB_LUT4 i12897_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17642));   // verilog/coms.v(126[12] 289[6])
    defparam i12897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12898_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17643));   // verilog/coms.v(126[12] 289[6])
    defparam i12898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12899_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17644));   // verilog/coms.v(126[12] 289[6])
    defparam i12899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1623 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n36579));
    defparam i1_3_lut_adj_1623.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i2199_3_lut (.I0(n3238), .I1(n3305), .I2(n3263), .I3(GND_net), 
            .O(n3337));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12900_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17645));   // verilog/coms.v(126[12] 289[6])
    defparam i12900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1624 (.I0(n3054), .I1(n3042), .I2(n36579), .I3(n3055), 
            .O(n29_adj_4958));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i6_4_lut_adj_1624.LUT_INIT = 16'heccc;
    SB_LUT4 i14_4_lut_adj_1625 (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37_adj_4956));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 add_577_18_lut (.I0(duty[16]), .I1(n44224), .I2(n9_adj_4317), 
            .I3(n28677), .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2858), .I1(VCC_net), 
            .CO(n29428));
    SB_LUT4 i13_4_lut_adj_1626 (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36_adj_4957));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i12901_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[19] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17646));   // verilog/coms.v(126[12] 289[6])
    defparam i12901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12902_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[19] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17647));   // verilog/coms.v(126[12] 289[6])
    defparam i12902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550_adj_4501), .I1(n2617), .I2(n2570), 
            .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut_adj_1627 (.I0(n37_adj_4956), .I1(n29_adj_4958), .I2(n3043), 
            .I3(n3048), .O(n42_adj_4952));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i19_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1628 (.I0(n3234), .I1(n3337), .I2(n3301), .I3(n3263), 
            .O(n38463));
    defparam i1_4_lut_adj_1628.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_add_1921_27_lut (.I0(n2867), .I1(n2834), .I2(VCC_net), 
            .I3(n29427), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i17_4_lut_adj_1629 (.I0(n3045), .I1(n3053), .I2(n3047), .I3(n3050), 
            .O(n40_adj_4954));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i17_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i12903_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[19] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17648));   // verilog/coms.v(126[12] 289[6])
    defparam i12903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut (.I0(n3044), .I1(n36_adj_4957), .I2(n3033), .I3(n3032), 
            .O(n41_adj_4953));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1921_26_lut (.I0(GND_net), .I1(n2835), .I2(VCC_net), 
            .I3(n29426), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12904_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[19] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17649));   // verilog/coms.v(126[12] 289[6])
    defparam i12904_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_26 (.CI(n29426), .I0(n2835), .I1(VCC_net), 
            .CO(n29427));
    SB_CARRY add_577_18 (.CI(n28677), .I0(n44224), .I1(n9_adj_4317), .CO(n28678));
    SB_LUT4 i12905_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[19] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17650));   // verilog/coms.v(126[12] 289[6])
    defparam i12905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2836), .I2(VCC_net), 
            .I3(n29425), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_5 (.CI(n29154), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n29155));
    SB_CARRY rem_4_add_1921_25 (.CI(n29425), .I0(n2836), .I1(VCC_net), 
            .CO(n29426));
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2837), .I2(VCC_net), 
            .I3(n29424), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_24 (.CI(n29424), .I0(n2837), .I1(VCC_net), 
            .CO(n29425));
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2838), .I2(VCC_net), 
            .I3(n29423), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2192_3_lut (.I0(n3231), .I1(n3298), .I2(n3263), .I3(GND_net), 
            .O(n3330));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut (.I0(n3046), .I1(n3051), .I2(n3049), .I3(n3052), 
            .O(n39_adj_4955));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4955), .I1(n41_adj_4953), .I2(n40_adj_4954), 
            .I3(n42_adj_4952), .O(n3065));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12906_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[19] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17651));   // verilog/coms.v(126[12] 289[6])
    defparam i12906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1199_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n29153), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(n47), .I1(n46), .I2(n28), .I3(n38651), 
            .O(n38657));
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28_adj_4417), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1631 (.I0(n3232), .I1(n38463), .I2(n3299), .I3(n3263), 
            .O(n38465));
    defparam i1_4_lut_adj_1631.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(n38986), .I1(n38465), .I2(n38657), 
            .I3(n3330), .O(n3362));
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i12907_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[19] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17652));   // verilog/coms.v(126[12] 289[6])
    defparam i12907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4556));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_23 (.CI(n29423), .I0(n2838), .I1(VCC_net), 
            .CO(n29424));
    SB_LUT4 i12908_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[18] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17653));   // verilog/coms.v(126[12] 289[6])
    defparam i12908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12909_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[18] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17654));   // verilog/coms.v(126[12] 289[6])
    defparam i12909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37319_2_lut (.I0(n3362), .I1(n10218), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37319_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12910_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[18] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17655));   // verilog/coms.v(126[12] 289[6])
    defparam i12910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1633 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n36527));
    defparam i1_3_lut_adj_1633.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2839), .I2(VCC_net), 
            .I3(n29422), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1634 (.I0(n3154), .I1(n3142), .I2(n36527), .I3(n3155), 
            .O(n31_adj_4883));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i7_4_lut_adj_1634.LUT_INIT = 16'heccc;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4920));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1707_3_lut_3_lut (.I0(n2558), .I1(n6114), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551_adj_4500), .I1(n2618_adj_4491), 
            .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_22 (.CI(n29422), .I0(n2839), .I1(VCC_net), 
            .CO(n29423));
    SB_CARRY communication_counter_1199_add_4_4 (.CI(n29153), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n29154));
    SB_LUT4 communication_counter_1199_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n29152), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n29421), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1199_add_4_3 (.CI(n29152), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n29153));
    SB_LUT4 communication_counter_1199_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1199_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_21 (.CI(n29421), .I0(n2840), .I1(VCC_net), 
            .CO(n29422));
    SB_LUT4 i12911_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[18] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17656));   // verilog/coms.v(126[12] 289[6])
    defparam i12911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12912_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[18] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17657));   // verilog/coms.v(126[12] 289[6])
    defparam i12912_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1199_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n29152));
    SB_LUT4 i12913_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[18] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17658));   // verilog/coms.v(126[12] 289[6])
    defparam i12913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13213_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n35433), .I3(GND_net), .O(n17958));   // verilog/coms.v(126[12] 289[6])
    defparam i13213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12914_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[18] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17659));   // verilog/coms.v(126[12] 289[6])
    defparam i12914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12915_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[18] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17660));   // verilog/coms.v(126[12] 289[6])
    defparam i12915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12916_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[17] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17661));   // verilog/coms.v(126[12] 289[6])
    defparam i12916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12917_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[17] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17662));   // verilog/coms.v(126[12] 289[6])
    defparam i12917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12918_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[17] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17663));   // verilog/coms.v(126[12] 289[6])
    defparam i12918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_4_lut_adj_1635 (.I0(n3137), .I1(n3138), .I2(n3143), .I3(n3140), 
            .O(n39_adj_4881));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i15_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i12919_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[17] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17664));   // verilog/coms.v(126[12] 289[6])
    defparam i12919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3139), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4884));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12920_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[17] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17665));   // verilog/coms.v(126[12] 289[6])
    defparam i12920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12921_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[17] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17666));   // verilog/coms.v(126[12] 289[6])
    defparam i12921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1636 (.I0(n3134), .I1(n3135), .I2(n3136), .I3(n3141), 
            .O(n38_adj_4882));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n39_adj_4881), .I1(n31_adj_4883), .I2(n3152), 
            .I3(n3150), .O(n44_adj_4877));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1637 (.I0(n3149), .I1(n3148), .I2(n3153), .I3(n3146), 
            .O(n42_adj_4879));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i18_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i12922_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[17] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17667));   // verilog/coms.v(126[12] 289[6])
    defparam i12922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12923_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[17] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17668));   // verilog/coms.v(126[12] 289[6])
    defparam i12923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12924_3_lut (.I0(Kp[1]), .I1(\data_in_frame[2] [1]), .I2(n17068), 
            .I3(GND_net), .O(n17669));   // verilog/coms.v(126[12] 289[6])
    defparam i12924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13214_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n35433), .I3(GND_net), .O(n17959));   // verilog/coms.v(126[12] 289[6])
    defparam i13214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19_4_lut_adj_1638 (.I0(n3132), .I1(n38_adj_4882), .I2(n26_adj_4884), 
            .I3(n3131), .O(n43_adj_4878));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i19_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n44170), .I1(n2_adj_4920), .I2(n3452), 
            .I3(n29151), .O(color_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n29420), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_20 (.CI(n29420), .I0(n2841), .I1(VCC_net), 
            .CO(n29421));
    SB_LUT4 i12925_3_lut (.I0(Kp[2]), .I1(\data_in_frame[2] [2]), .I2(n17068), 
            .I3(GND_net), .O(n17670));   // verilog/coms.v(126[12] 289[6])
    defparam i12925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n29419), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n44174), .I1(n2_adj_4920), .I2(n3453), 
            .I3(n29150), .O(color_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_8 (.CI(n29150), .I0(n2_adj_4920), .I1(n3453), 
            .CO(n29151));
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n44177), .I1(n2_adj_4920), .I2(n3454), 
            .I3(n29149), .O(color_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1921_19 (.CI(n29419), .I0(n2842), .I1(VCC_net), 
            .CO(n29420));
    SB_LUT4 add_577_17_lut (.I0(duty[15]), .I1(n44224), .I2(n10_adj_4318), 
            .I3(n28676), .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4555));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1639 (.I0(n3147), .I1(n3145), .I2(n3144), .I3(n3151), 
            .O(n41_adj_4880));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i17_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_2298_7 (.CI(n29149), .I0(n2_adj_4920), .I1(n3454), 
            .CO(n29150));
    SB_LUT4 i12926_3_lut (.I0(Kp[3]), .I1(\data_in_frame[2] [3]), .I2(n17068), 
            .I3(GND_net), .O(n17671));   // verilog/coms.v(126[12] 289[6])
    defparam i12926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n44180), .I1(n2_adj_4920), .I2(n3455), 
            .I3(n29148), .O(color_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i23_4_lut (.I0(n41_adj_4880), .I1(n43_adj_4878), .I2(n42_adj_4879), 
            .I3(n44_adj_4877), .O(n3164));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12927_3_lut (.I0(Kp[4]), .I1(\data_in_frame[2] [4]), .I2(n17068), 
            .I3(GND_net), .O(n17672));   // verilog/coms.v(126[12] 289[6])
    defparam i12927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12928_3_lut (.I0(Kp[5]), .I1(\data_in_frame[2] [5]), .I2(n17068), 
            .I3(GND_net), .O(n17673));   // verilog/coms.v(126[12] 289[6])
    defparam i12928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13215_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n35433), .I3(GND_net), .O(n17960));   // verilog/coms.v(126[12] 289[6])
    defparam i13215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4416), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12929_3_lut (.I0(Kp[6]), .I1(\data_in_frame[2] [6]), .I2(n17068), 
            .I3(GND_net), .O(n17674));   // verilog/coms.v(126[12] 289[6])
    defparam i12929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12930_3_lut (.I0(Kp[7]), .I1(\data_in_frame[2] [7]), .I2(n17068), 
            .I3(GND_net), .O(n17675));   // verilog/coms.v(126[12] 289[6])
    defparam i12930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12931_3_lut (.I0(Ki[1]), .I1(\data_in_frame[3] [1]), .I2(n17068), 
            .I3(GND_net), .O(n17676));   // verilog/coms.v(126[12] 289[6])
    defparam i12931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1716_3_lut_3_lut (.I0(n2558), .I1(n6123), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1869_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), .I3(GND_net), 
            .O(n2847));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1872_3_lut (.I0(n2751), .I1(n2818), .I2(n2768), .I3(GND_net), 
            .O(n2850));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1873_3_lut (.I0(n2752), .I1(n2819), .I2(n2768), .I3(GND_net), 
            .O(n2851));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12932_3_lut (.I0(Ki[2]), .I1(\data_in_frame[3] [2]), .I2(n17068), 
            .I3(GND_net), .O(n17677));   // verilog/coms.v(126[12] 289[6])
    defparam i12932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12933_3_lut (.I0(Ki[3]), .I1(\data_in_frame[3] [3]), .I2(n17068), 
            .I3(GND_net), .O(n17678));   // verilog/coms.v(126[12] 289[6])
    defparam i12933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4927));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2298_6 (.CI(n29148), .I0(n2_adj_4920), .I1(n3455), 
            .CO(n29149));
    SB_LUT4 rem_4_i1868_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548_adj_4503), .I1(n2615), .I2(n2570), 
            .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30_adj_4415), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225), .I2(n3164), .I3(GND_net), 
            .O(n3257));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224), .I2(n3164), .I3(GND_net), 
            .O(n3256));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1640 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n36584));
    defparam i1_3_lut_adj_1640.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n44183), .I1(n2_adj_4920), .I2(n3456), 
            .I3(n29147), .O(color_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552_adj_4499), .I1(n2619_adj_4492), 
            .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1871_3_lut (.I0(n2750), .I1(n2817), .I2(n2768), .I3(GND_net), 
            .O(n2849));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547_adj_4504), .I1(n2614), .I2(n2570), 
            .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1739_3_lut (.I0(n2554), .I1(n2621_adj_4485), .I2(n2570), 
            .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538_adj_4513), .I1(n2605), .I2(n2570), 
            .I3(GND_net), .O(n2637_adj_4479));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553_adj_4498), .I1(n2620_adj_4486), 
            .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558_adj_4497), .I1(n2625_adj_4481), 
            .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4483), .I2(n2570), 
            .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4484), .I2(n2570), 
            .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4482), .I2(n2570), 
            .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1662_3_lut (.I0(n2445), .I1(n2512), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2544_adj_4507));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1661_3_lut (.I0(n2444), .I1(n2511), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2543_adj_4508));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1659_3_lut (.I0(n2442), .I1(n2509), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2541_adj_4510));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1668_3_lut (.I0(n2451_adj_4571), .I1(n2518), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2550_adj_4501));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1670_3_lut (.I0(n2453_adj_4569), .I1(n2520), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2552_adj_4499));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1669_3_lut (.I0(n2452_adj_4570), .I1(n2519), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2551_adj_4500));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1666_3_lut (.I0(n2449_adj_4573), .I1(n2516), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2548_adj_4503));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1667_3_lut (.I0(n2450_adj_4572), .I1(n2517), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2549_adj_4502));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1665_3_lut (.I0(n2448_adj_4574), .I1(n2515), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2547_adj_4504));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1671_3_lut (.I0(n2454_adj_4568), .I1(n2521), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2553_adj_4498));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1663_3_lut (.I0(n2446), .I1(n2513), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2545_adj_4506));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1664_3_lut (.I0(n2447_adj_4575), .I1(n2514), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2546_adj_4505));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1658_3_lut (.I0(n2441), .I1(n2508), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2540_adj_4511));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n29418), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_18 (.CI(n29418), .I0(n2843), .I1(VCC_net), 
            .CO(n29419));
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n29417), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_17 (.CI(n29417), .I0(n2844), .I1(VCC_net), 
            .CO(n29418));
    SB_CARRY rem_4_add_2298_5 (.CI(n29147), .I0(n2_adj_4920), .I1(n3456), 
            .CO(n29148));
    SB_LUT4 i17_4_lut_adj_1641 (.I0(n3252), .I1(n3253), .I2(n3247), .I3(n3248), 
            .O(n42));
    defparam i17_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1711_3_lut_3_lut (.I0(n2558), .I1(n6118), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1874_3_lut (.I0(n2753), .I1(n2820), .I2(n2768), .I3(GND_net), 
            .O(n2852));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n44186), .I1(n2_adj_4920), .I2(n3457), 
            .I3(n29146), .O(color_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n29416), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12934_3_lut (.I0(Ki[4]), .I1(\data_in_frame[3] [4]), .I2(n17068), 
            .I3(GND_net), .O(n17679));   // verilog/coms.v(126[12] 289[6])
    defparam i12934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12935_3_lut (.I0(Ki[5]), .I1(\data_in_frame[3] [5]), .I2(n17068), 
            .I3(GND_net), .O(n17680));   // verilog/coms.v(126[12] 289[6])
    defparam i12935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12936_3_lut (.I0(Ki[6]), .I1(\data_in_frame[3] [6]), .I2(n17068), 
            .I3(GND_net), .O(n17681));   // verilog/coms.v(126[12] 289[6])
    defparam i12936_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_16 (.CI(n29416), .I0(n2845), .I1(VCC_net), 
            .CO(n29417));
    SB_LUT4 i12937_3_lut (.I0(Ki[7]), .I1(\data_in_frame[3] [7]), .I2(n17068), 
            .I3(GND_net), .O(n17682));   // verilog/coms.v(126[12] 289[6])
    defparam i12937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12938_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17683));   // verilog/coms.v(126[12] 289[6])
    defparam i12938_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13157_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n35418), 
            .I3(GND_net), .O(n17902));   // verilog/coms.v(126[12] 289[6])
    defparam i13157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1674_3_lut (.I0(n2457_adj_4517), .I1(n2524), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2556));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32201_2_lut (.I0(start), .I1(one_wire_N_513[6]), .I2(GND_net), 
            .I3(GND_net), .O(n38981));
    defparam i32201_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32318_4_lut (.I0(one_wire_N_513[11]), .I1(one_wire_N_513[7]), 
            .I2(one_wire_N_513[8]), .I3(n38981), .O(n39099));
    defparam i32318_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n4_adj_4906), .I1(n39099), .I2(n106), .I3(one_wire_N_513[5]), 
            .O(n35266));
    defparam i8_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 div_46_i1710_3_lut_3_lut (.I0(n2558), .I1(n6117), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12939_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17684));   // verilog/coms.v(126[12] 289[6])
    defparam i12939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816), .I2(n2768), .I3(GND_net), 
            .O(n2848));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1642 (.I0(n3240), .I1(n3254), .I2(n36584), .I3(n3255), 
            .O(n31));
    defparam i6_4_lut_adj_1642.LUT_INIT = 16'heaaa;
    SB_LUT4 i13_3_lut (.I0(n3243), .I1(n3231), .I2(n3230), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1643 (.I0(n3250), .I1(n3251), .I2(n3249), .I3(n3244), 
            .O(n43));
    defparam i18_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1644 (.I0(n3236), .I1(n3238), .I2(n3237), .I3(n3239), 
            .O(n40));
    defparam i15_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n29415), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821), .I2(n2768), .I3(GND_net), 
            .O(n2853));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1645 (.I0(n2349), .I1(n2348), .I2(n2353), .I3(n2350), 
            .O(n28_adj_4902));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_2298_4 (.CI(n29146), .I0(n2_adj_4920), .I1(n3457), 
            .CO(n29147));
    SB_CARRY rem_4_add_1921_15 (.CI(n29415), .I0(n2846), .I1(VCC_net), 
            .CO(n29416));
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n36482), 
            .O(n26_adj_4904));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1646 (.I0(n1647_adj_4463), .I1(n1646_adj_4462), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4875));
    defparam i1_2_lut_adj_1646.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1647 (.I0(n2346), .I1(n2351), .I2(n2347), .I3(n2352), 
            .O(n27_adj_4903));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1713_3_lut_3_lut (.I0(n2558), .I1(n6120), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_4920), 
            .I2(n3458), .I3(n29145), .O(color_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n29414), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_14 (.CI(n29414), .I0(n2847), .I1(VCC_net), 
            .CO(n29415));
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2298_3 (.CI(n29145), .I0(n2_adj_4920), .I1(n3458), 
            .CO(n29146));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_4920), 
            .I2(n3459), .I3(VCC_net), .O(color_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_4920), .I1(n3459), 
            .CO(n29145));
    SB_CARRY add_577_17 (.CI(n28676), .I0(n44224), .I1(n10_adj_4318), 
            .CO(n28677));
    SB_LUT4 div_46_i1715_3_lut_3_lut (.I0(n2558), .I1(n6122), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_577_16_lut (.I0(duty[14]), .I1(n44224), .I2(n11), .I3(n28675), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n29413), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12940_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17685));   // verilog/coms.v(126[12] 289[6])
    defparam i12940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12941_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17686));   // verilog/coms.v(126[12] 289[6])
    defparam i12941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_13 (.CI(n29413), .I0(n2848), .I1(VCC_net), 
            .CO(n29414));
    SB_LUT4 i12942_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17687));   // verilog/coms.v(126[12] 289[6])
    defparam i12942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12943_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17688));   // verilog/coms.v(126[12] 289[6])
    defparam i12943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_577_16 (.CI(n28675), .I0(n44224), .I1(n11), .CO(n28676));
    SB_LUT4 add_2297_25_lut (.I0(n249), .I1(n44228), .I2(n248), .I3(n29144), 
            .O(displacement_23__N_229[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_577_15_lut (.I0(duty[13]), .I1(n44224), .I2(n12), .I3(n28674), 
            .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2297_24_lut (.I0(n393), .I1(n44228), .I2(n392), .I3(n29143), 
            .O(displacement_23__N_229[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12944_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17689));   // verilog/coms.v(126[12] 289[6])
    defparam i12944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12945_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17690));   // verilog/coms.v(126[12] 289[6])
    defparam i12945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12946_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17691));   // verilog/coms.v(126[12] 289[6])
    defparam i12946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4554));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n29412), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_12 (.CI(n29412), .I0(n2849), .I1(VCC_net), 
            .CO(n29413));
    SB_CARRY add_2297_24 (.CI(n29143), .I0(n44228), .I1(n392), .CO(n29144));
    SB_LUT4 add_2297_23_lut (.I0(n534), .I1(n44228), .I2(n533), .I3(n29142), 
            .O(displacement_23__N_229[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12947_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17692));   // verilog/coms.v(126[12] 289[6])
    defparam i12947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n29411), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_23 (.CI(n29142), .I0(n44228), .I1(n533), .CO(n29143));
    SB_LUT4 i21_4_lut (.I0(n31), .I1(n42), .I2(n3241), .I3(n3242), .O(n46_adj_4346));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2297_22_lut (.I0(n672), .I1(n44228), .I2(n671), .I3(n29141), 
            .O(displacement_23__N_229[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12948_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17693));   // verilog/coms.v(126[12] 289[6])
    defparam i12948_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_11 (.CI(n29411), .I0(n2850), .I1(VCC_net), 
            .CO(n29412));
    SB_LUT4 i12949_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17694));   // verilog/coms.v(126[12] 289[6])
    defparam i12949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1648 (.I0(n3232), .I1(n3234), .I2(n3233), .I3(n3235), 
            .O(n39));
    defparam i14_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i12950_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17695));   // verilog/coms.v(126[12] 289[6])
    defparam i12950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825), .I2(n2768), .I3(GND_net), 
            .O(n2857));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12951_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17696));   // verilog/coms.v(126[12] 289[6])
    defparam i12951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_4_lut_adj_1649 (.I0(n43), .I1(n3245), .I2(n38), .I3(n3246), 
            .O(n47_adj_4345));
    defparam i22_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4345), .I1(n39), .I2(n46_adj_4346), 
            .I3(n40), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4553));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824), .I2(n2768), .I3(GND_net), 
            .O(n2856));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12952_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17697));   // verilog/coms.v(126[12] 289[6])
    defparam i12952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12953_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17698));   // verilog/coms.v(126[12] 289[6])
    defparam i12953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12954_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17699));   // verilog/coms.v(126[12] 289[6])
    defparam i12954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n29410), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_10 (.CI(n29410), .I0(n2851), .I1(VCC_net), 
            .CO(n29411));
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n29409), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_9 (.CI(n29409), .I0(n2852), .I1(VCC_net), 
            .CO(n29410));
    SB_CARRY add_577_15 (.CI(n28674), .I0(n44224), .I1(n12), .CO(n28675));
    SB_CARRY add_2297_22 (.CI(n29141), .I0(n44228), .I1(n671), .CO(n29142));
    SB_LUT4 i12955_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17700));   // verilog/coms.v(126[12] 289[6])
    defparam i12955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13092_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13293), .I3(GND_net), .O(n17837));   // verilog/coms.v(126[12] 289[6])
    defparam i13092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13093_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13293), .I3(GND_net), .O(n17838));   // verilog/coms.v(126[12] 289[6])
    defparam i13093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13094_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13293), .I3(GND_net), .O(n17839));   // verilog/coms.v(126[12] 289[6])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13095_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13293), .I3(GND_net), .O(n17840));   // verilog/coms.v(126[12] 289[6])
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13096_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13293), .I3(GND_net), .O(n17841));   // verilog/coms.v(126[12] 289[6])
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13097_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13293), .I3(GND_net), .O(n17842));   // verilog/coms.v(126[12] 289[6])
    defparam i13097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13098_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13293), .I3(GND_net), .O(n17843));   // verilog/coms.v(126[12] 289[6])
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13228_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n35435), .I3(GND_net), .O(n17973));   // verilog/coms.v(126[12] 289[6])
    defparam i13228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823), .I2(n2768), .I3(GND_net), 
            .O(n2855_adj_4434));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12956_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17701));   // verilog/coms.v(126[12] 289[6])
    defparam i12956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12957_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17702));   // verilog/coms.v(126[12] 289[6])
    defparam i12957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13099_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13293), .I3(GND_net), .O(n17844));   // verilog/coms.v(126[12] 289[6])
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822), .I2(n2768), .I3(GND_net), 
            .O(n2854));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12958_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17703));   // verilog/coms.v(126[12] 289[6])
    defparam i12958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n29408), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13100_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17845));   // verilog/coms.v(126[12] 289[6])
    defparam i13100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1650 (.I0(n2856), .I1(n2857), .I2(n2858), .I3(GND_net), 
            .O(n36571));
    defparam i1_3_lut_adj_1650.LUT_INIT = 16'hfefe;
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4321));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12959_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17704));   // verilog/coms.v(126[12] 289[6])
    defparam i12959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12960_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17705));   // verilog/coms.v(126[12] 289[6])
    defparam i12960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12961_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17706));   // verilog/coms.v(126[12] 289[6])
    defparam i12961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12962_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17707));   // verilog/coms.v(126[12] 289[6])
    defparam i12962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_577_14_lut (.I0(duty[12]), .I1(n44224), .I2(n13), .I3(n28673), 
            .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12963_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17708));   // verilog/coms.v(126[12] 289[6])
    defparam i12963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12964_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17709));   // verilog/coms.v(126[12] 289[6])
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13101_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n17068), .I3(GND_net), .O(n17846));   // verilog/coms.v(126[12] 289[6])
    defparam i13101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12965_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17710));   // verilog/coms.v(126[12] 289[6])
    defparam i12965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13102_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n17068), .I3(GND_net), .O(n17847));   // verilog/coms.v(126[12] 289[6])
    defparam i13102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2297_21_lut (.I0(n807), .I1(n44228), .I2(n806), .I3(n29140), 
            .O(displacement_23__N_229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13217_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n35433), .I3(GND_net), .O(n17962));   // verilog/coms.v(126[12] 289[6])
    defparam i13217_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2297_21 (.CI(n29140), .I0(n44228), .I1(n806), .CO(n29141));
    SB_LUT4 i1_3_lut_adj_1651 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n36457));
    defparam i1_3_lut_adj_1651.LUT_INIT = 16'hfefe;
    SB_CARRY add_577_14 (.CI(n28673), .I0(n44224), .I1(n13), .CO(n28674));
    SB_CARRY rem_4_add_1921_8 (.CI(n29408), .I0(n2853), .I1(VCC_net), 
            .CO(n29409));
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4552));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1652 (.I0(n1653_adj_4460), .I1(n1652_adj_4459), 
            .I2(n1651_adj_4467), .I3(n10_adj_4875), .O(n16_adj_4873));
    defparam i7_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2297_20_lut (.I0(n939), .I1(n44228), .I2(n938), .I3(n29139), 
            .O(displacement_23__N_229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_983_13_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n29672), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_983_12_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n29671), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12966_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17711));   // verilog/coms.v(126[12] 289[6])
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1653 (.I0(n2842), .I1(n2854), .I2(n36571), .I3(n2855_adj_4434), 
            .O(n26_adj_4972));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_4_lut_adj_1653.LUT_INIT = 16'heaaa;
    SB_LUT4 i12967_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17712));   // verilog/coms.v(126[12] 289[6])
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1654 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_4905));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i9_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i12968_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17713));   // verilog/coms.v(126[12] 289[6])
    defparam i12968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1655 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33_adj_4970));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_983_12 (.CI(n29671), .I0(n1449), .I1(VCC_net), 
            .CO(n29672));
    SB_LUT4 i12969_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID0), .I2(n13293), 
            .I3(GND_net), .O(n17714));   // verilog/coms.v(126[12] 289[6])
    defparam i12969_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2297_20 (.CI(n29139), .I0(n44228), .I1(n938), .CO(n29140));
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n29407), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2297_19_lut (.I0(n1068), .I1(n44228), .I2(n1067), .I3(n29138), 
            .O(displacement_23__N_229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n29670), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2297_19 (.CI(n29138), .I0(n44228), .I1(n1067), .CO(n29139));
    SB_CARRY rem_4_add_983_11 (.CI(n29670), .I0(n1450), .I1(VCC_net), 
            .CO(n29671));
    SB_LUT4 i13103_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n17068), .I3(GND_net), .O(n17848));   // verilog/coms.v(126[12] 289[6])
    defparam i13103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n29669), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4973));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_983_10 (.CI(n29669), .I0(n1451), .I1(VCC_net), 
            .CO(n29670));
    SB_LUT4 div_46_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4551));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13104_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n17068), .I3(GND_net), .O(n17849));   // verilog/coms.v(126[12] 289[6])
    defparam i13104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4926));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1657 (.I0(n33_adj_4970), .I1(n2840), .I2(n26_adj_4972), 
            .I3(n2841), .O(n38_adj_4966));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i17_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i13105_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n17068), .I3(GND_net), .O(n17850));   // verilog/coms.v(126[12] 289[6])
    defparam i13105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n29668), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_9 (.CI(n29668), .I0(n1452), .I1(VCC_net), .CO(n29669));
    SB_CARRY rem_4_add_1921_7 (.CI(n29407), .I0(n2854), .I1(GND_net), 
            .CO(n29408));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n29667), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_8 (.CI(n29667), .I0(n1453), .I1(VCC_net), .CO(n29668));
    SB_LUT4 i13106_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n17068), .I3(GND_net), .O(n17851));   // verilog/coms.v(126[12] 289[6])
    defparam i13106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2855_adj_4434), .I2(GND_net), 
            .I3(n29406), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_CARRY rem_4_add_1921_6 (.CI(n29406), .I0(n2855_adj_4434), .I1(GND_net), 
            .CO(n29407));
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4320));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1658 (.I0(n2853), .I1(n2848), .I2(n2845), .I3(n2852), 
            .O(n36_adj_4968));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i15_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4550));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13107_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n35419), 
            .I3(GND_net), .O(n17852));   // verilog/coms.v(126[12] 289[6])
    defparam i13107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1659 (.I0(n2851), .I1(n2850), .I2(n2847), .I3(n22_adj_4973), 
            .O(n37_adj_4967));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i16_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4925));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4924));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4549));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_LUT4 i13108_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n35419), 
            .I3(GND_net), .O(n17853));   // verilog/coms.v(126[12] 289[6])
    defparam i13108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4548));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13109_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n35419), 
            .I3(GND_net), .O(n17854));   // verilog/coms.v(126[12] 289[6])
    defparam i13109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4923));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13110_3_lut (.I0(\data_in_frame[0] [4]), .I1(rx_data[4]), .I2(n35419), 
            .I3(GND_net), .O(n17855));   // verilog/coms.v(126[12] 289[6])
    defparam i13110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut_adj_1660 (.I0(n2843), .I1(n2849), .I2(n2844), .I3(n2846), 
            .O(n35_adj_4969));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1661 (.I0(n1648_adj_4464), .I1(n1654), .I2(n36457), 
            .I3(n1655), .O(n11_adj_4874));
    defparam i2_4_lut_adj_1661.LUT_INIT = 16'heaaa;
    SB_LUT4 i12970_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID1), .I2(n13293), 
            .I3(GND_net), .O(n17715));   // verilog/coms.v(126[12] 289[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13111_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n35419), 
            .I3(GND_net), .O(n17856));   // verilog/coms.v(126[12] 289[6])
    defparam i13111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12971_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID2), .I2(n13293), 
            .I3(GND_net), .O(n17716));   // verilog/coms.v(126[12] 289[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12972_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13293), .I3(GND_net), .O(n17717));   // verilog/coms.v(126[12] 289[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_4_lut_adj_1662 (.I0(n35_adj_4969), .I1(n37_adj_4967), .I2(n36_adj_4968), 
            .I3(n38_adj_4966), .O(n2867));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i20_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1768_3_lut_3_lut (.I0(n2642), .I1(n6143), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12973_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13293), .I3(GND_net), .O(n17718));   // verilog/coms.v(126[12] 289[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13112_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n35419), 
            .I3(GND_net), .O(n17857));   // verilog/coms.v(126[12] 289[6])
    defparam i13112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12974_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13293), .I3(GND_net), .O(n17719));   // verilog/coms.v(126[12] 289[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_LUT4 add_577_13_lut (.I0(duty[11]), .I1(n44224), .I2(n14), .I3(n28672), 
            .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_13_lut.LUT_INIT = 16'h8BB8;
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_LUT4 add_2297_18_lut (.I0(n1194), .I1(n44228), .I2(n1193), .I3(n29137), 
            .O(displacement_23__N_229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_18_lut.LUT_INIT = 16'h8BB8;
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_LUT4 div_46_i1755_3_lut_3_lut (.I0(n2642), .I1(n6130), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_LUT4 i13113_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n35419), 
            .I3(GND_net), .O(n17858));   // verilog/coms.v(126[12] 289[6])
    defparam i13113_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(251[10] 253[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_CARRY add_2297_18 (.CI(n29137), .I0(n44228), .I1(n1193), .CO(n29138));
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_CARRY add_577_13 (.CI(n28672), .I0(n44224), .I1(n14), .CO(n28673));
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 i12975_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13293), .I3(GND_net), .O(n17720));   // verilog/coms.v(126[12] 289[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 add_2297_17_lut (.I0(n1317), .I1(n44228), .I2(n1316), .I3(n29136), 
            .O(displacement_23__N_229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_17_lut.LUT_INIT = 16'h8BB8;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 add_577_12_lut (.I0(duty[10]), .I1(n44224), .I2(n15_adj_4319), 
            .I3(n28671), .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_12_lut.LUT_INIT = 16'h8BB8;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_CARRY add_2297_17 (.CI(n29136), .I0(n44228), .I1(n1316), .CO(n29137));
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n29405), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2297_16_lut (.I0(n1437), .I1(n44228), .I2(n1436), .I3(n29135), 
            .O(displacement_23__N_229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_16_lut.LUT_INIT = 16'h8BB8;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(163[10] 176[6])
    SB_LUT4 i13218_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n35434), .I3(GND_net), .O(n17963));   // verilog/coms.v(126[12] 289[6])
    defparam i13218_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2297_16 (.CI(n29135), .I0(n44228), .I1(n1436), .CO(n29136));
    SB_LUT4 add_2297_15_lut (.I0(n1554), .I1(n44228), .I2(n1553), .I3(n29134), 
            .O(displacement_23__N_229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_15 (.CI(n29134), .I0(n44228), .I1(n1553), .CO(n29135));
    SB_LUT4 i13282_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[7] [1]), 
            .I2(n17068), .I3(GND_net), .O(n18027));   // verilog/coms.v(126[12] 289[6])
    defparam i13282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13283_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[7] [2]), 
            .I2(n17068), .I3(GND_net), .O(n18028));   // verilog/coms.v(126[12] 289[6])
    defparam i13283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13284_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[7] [3]), 
            .I2(n17068), .I3(GND_net), .O(n18029));   // verilog/coms.v(126[12] 289[6])
    defparam i13284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n29666), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_5 (.CI(n29405), .I0(n2856), .I1(VCC_net), 
            .CO(n29406));
    SB_LUT4 i13285_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[7] [4]), 
            .I2(n17068), .I3(GND_net), .O(n18030));   // verilog/coms.v(126[12] 289[6])
    defparam i13285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2297_14_lut (.I0(n1668), .I1(n44228), .I2(n1667), .I3(n29133), 
            .O(displacement_23__N_229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13286_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[7] [5]), 
            .I2(n17068), .I3(GND_net), .O(n18031));   // verilog/coms.v(126[12] 289[6])
    defparam i13286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1673_3_lut (.I0(n2456_adj_4518), .I1(n2523), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2555));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2297_14 (.CI(n29133), .I0(n44228), .I1(n1667), .CO(n29134));
    SB_LUT4 add_2297_13_lut (.I0(n1779), .I1(n44228), .I2(n1778), .I3(n29132), 
            .O(displacement_23__N_229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13287_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[7] [6]), 
            .I2(n17068), .I3(GND_net), .O(n18032));   // verilog/coms.v(126[12] 289[6])
    defparam i13287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13288_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[7] [7]), 
            .I2(n17068), .I3(GND_net), .O(n18033));   // verilog/coms.v(126[12] 289[6])
    defparam i13288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13289_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[6] [0]), 
            .I2(n17068), .I3(GND_net), .O(n18034));   // verilog/coms.v(126[12] 289[6])
    defparam i13289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13290_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[6] [1]), 
            .I2(n17068), .I3(GND_net), .O(n18035));   // verilog/coms.v(126[12] 289[6])
    defparam i13290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13114_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n35420), 
            .I3(GND_net), .O(n17859));   // verilog/coms.v(126[12] 289[6])
    defparam i13114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1657_3_lut (.I0(n2440), .I1(n2507), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2539_adj_4512));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1656_3_lut (.I0(n2439), .I1(n2506), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2538_adj_4513));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1663 (.I0(n2538_adj_4513), .I1(n2539_adj_4512), 
            .I2(n2537_adj_4514), .I3(n2540_adj_4511), .O(n28_adj_4412));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1664 (.I0(n2556), .I1(n2558_adj_4497), .I2(GND_net), 
            .I3(GND_net), .O(n38755));
    defparam i1_2_lut_adj_1664.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1665 (.I0(n2554), .I1(n38755), .I2(n2555), .I3(n2557), 
            .O(n36486));
    defparam i1_4_lut_adj_1665.LUT_INIT = 16'ha080;
    SB_LUT4 i14_3_lut (.I0(n2547_adj_4504), .I1(n28_adj_4412), .I2(n2549_adj_4502), 
            .I3(GND_net), .O(n32));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_2297_13 (.CI(n29132), .I0(n44228), .I1(n1778), .CO(n29133));
    SB_LUT4 i13115_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n35420), 
            .I3(GND_net), .O(n17860));   // verilog/coms.v(126[12] 289[6])
    defparam i13115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1666 (.I0(n36486), .I1(n2546_adj_4505), .I2(n2545_adj_4506), 
            .I3(n2553_adj_4498), .O(n30));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2297_12_lut (.I0(n1887), .I1(n44228), .I2(n1886), .I3(n29131), 
            .O(displacement_23__N_229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13_4_lut_adj_1667 (.I0(n2548_adj_4503), .I1(n2551_adj_4500), 
            .I2(n2552_adj_4499), .I3(n2550_adj_4501), .O(n31_adj_4411));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2857), .I2(VCC_net), 
            .I3(n29404), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_12 (.CI(n29131), .I0(n44228), .I1(n1886), .CO(n29132));
    SB_CARRY rem_4_add_1921_4 (.CI(n29404), .I0(n2857), .I1(VCC_net), 
            .CO(n29405));
    SB_LUT4 add_2297_11_lut (.I0(n1992), .I1(n44228), .I2(n1991), .I3(n29130), 
            .O(displacement_23__N_229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_11 (.CI(n29130), .I0(n44228), .I1(n1991), .CO(n29131));
    SB_LUT4 add_2297_10_lut (.I0(n2094), .I1(n44228), .I2(n2093), .I3(n29129), 
            .O(displacement_23__N_229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_10 (.CI(n29129), .I0(n44228), .I1(n2093), .CO(n29130));
    SB_LUT4 add_2297_9_lut (.I0(n2193), .I1(n44228), .I2(n2192), .I3(n29128), 
            .O(displacement_23__N_229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_983_7 (.CI(n29666), .I0(n1454), .I1(GND_net), .CO(n29667));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2858), .I2(GND_net), 
            .I3(n29403), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_9 (.CI(n29128), .I0(n44228), .I1(n2192), .CO(n29129));
    SB_LUT4 add_2297_8_lut (.I0(n2289), .I1(n44228), .I2(n2288), .I3(n29127), 
            .O(displacement_23__N_229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_8 (.CI(n29127), .I0(n44228), .I1(n2288), .CO(n29128));
    SB_LUT4 add_2297_7_lut (.I0(n2382), .I1(n44228), .I2(n2381), .I3(n29126), 
            .O(displacement_23__N_229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1921_3 (.CI(n29403), .I0(n2858), .I1(GND_net), 
            .CO(n29404));
    SB_LUT4 i13116_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n35420), 
            .I3(GND_net), .O(n17861));   // verilog/coms.v(126[12] 289[6])
    defparam i13116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2297_7 (.CI(n29126), .I0(n44228), .I1(n2381), .CO(n29127));
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2958_adj_4401), .I1(VCC_net), 
            .CO(n29403));
    SB_LUT4 add_2297_6_lut (.I0(n2472), .I1(n44228), .I2(n2471), .I3(n29125), 
            .O(displacement_23__N_229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_6 (.CI(n29125), .I0(n44228), .I1(n2471), .CO(n29126));
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n29665), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2297_5_lut (.I0(n2559), .I1(n44228), .I2(n2558), .I3(n29124), 
            .O(displacement_23__N_229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4543), .I3(n29402), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2297_5 (.CI(n29124), .I0(n44228), .I1(n2558), .CO(n29125));
    SB_LUT4 add_2297_4_lut (.I0(n2643), .I1(n44228), .I2(n2642), .I3(n29123), 
            .O(displacement_23__N_229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2297_4 (.CI(n29123), .I0(n44228), .I1(n2642), .CO(n29124));
    SB_LUT4 div_46_i1754_3_lut_3_lut (.I0(n2642), .I1(n6129), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2297_3_lut (.I0(n2724), .I1(n44228), .I2(n2723), .I3(n29122), 
            .O(displacement_23__N_229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4544), .I3(n29401), .O(n3_adj_4371)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_1668 (.I0(n11_adj_4874), .I1(n16_adj_4873), .I2(n1649_adj_4465), 
            .I3(n1650_adj_4466), .O(n1679));
    defparam i8_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_CARRY add_2297_3 (.CI(n29122), .I0(n44228), .I1(n2723), .CO(n29123));
    SB_CARRY div_46_unary_minus_2_add_3_24 (.CI(n29401), .I0(GND_net), .I1(n3_adj_4544), 
            .CO(n29402));
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_4920), .I3(n30501), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4921), .I3(n30500), .O(n3_adj_4475)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n30500), .I0(GND_net), .I1(n3_adj_4921), 
            .CO(n30501));
    SB_CARRY rem_4_add_983_6 (.CI(n29665), .I0(n1455), .I1(GND_net), .CO(n29666));
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2858));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4317));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4545), .I3(n29400), .O(n4_adj_4370)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n29664), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_23 (.CI(n29400), .I0(GND_net), .I1(n4_adj_4545), 
            .CO(n29401));
    SB_CARRY rem_4_add_983_5 (.CI(n29664), .I0(n1456), .I1(VCC_net), .CO(n29665));
    SB_LUT4 div_46_i1756_3_lut_3_lut (.I0(n2642), .I1(n6131), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4546), .I3(n29399), .O(n5_adj_4369)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_22 (.CI(n29399), .I0(GND_net), .I1(n5_adj_4546), 
            .CO(n29400));
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n29663), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_4 (.CI(n29663), .I0(n1457), .I1(VCC_net), .CO(n29664));
    SB_LUT4 add_2297_2_lut (.I0(n2802), .I1(n44228), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4547), .I3(n29398), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13117_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n35420), 
            .I3(GND_net), .O(n17862));   // verilog/coms.v(126[12] 289[6])
    defparam i13117_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2297_2 (.CI(VCC_net), .I0(n44228), .I1(n2801), .CO(n29122));
    SB_LUT4 i11_4_lut_adj_1669 (.I0(n2541_adj_4510), .I1(n2543_adj_4508), 
            .I2(n2542_adj_4509), .I3(n2544_adj_4507), .O(n29));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2296_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n29121), 
            .O(n6153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4922), .I3(n30499), .O(n4_adj_4474)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13118_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n35420), 
            .I3(GND_net), .O(n17863));   // verilog/coms.v(126[12] 289[6])
    defparam i13118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(n29662), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13119_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n35420), 
            .I3(GND_net), .O(n17864));   // verilog/coms.v(126[12] 289[6])
    defparam i13119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1758_3_lut_3_lut (.I0(n2642), .I1(n6133), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13120_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n35420), 
            .I3(GND_net), .O(n17865));   // verilog/coms.v(126[12] 289[6])
    defparam i13120_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n30499), .I0(GND_net), .I1(n4_adj_4922), 
            .CO(n30500));
    SB_CARRY div_46_unary_minus_2_add_3_21 (.CI(n29398), .I0(GND_net), .I1(n6_adj_4547), 
            .CO(n29399));
    SB_LUT4 add_2296_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n29120), 
            .O(n6154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1670 (.I0(n25_adj_4905), .I1(n27_adj_4903), .I2(n26_adj_4904), 
            .I3(n28_adj_4902), .O(n2372_adj_4577));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i15_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1757_3_lut_3_lut (.I0(n2642), .I1(n6132), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4923), .I3(n30498), .O(n5_adj_4473)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_24 (.CI(n29120), .I0(n2700), .I1(n79), .CO(n29121));
    SB_LUT4 add_2296_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n29119), 
            .O(n6155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4548), .I3(n29397), .O(n7_adj_4312)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_20 (.CI(n29397), .I0(GND_net), .I1(n7_adj_4548), 
            .CO(n29398));
    SB_LUT4 div_46_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4549), .I3(n29396), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n30498), .I0(GND_net), .I1(n5_adj_4923), 
            .CO(n30499));
    SB_CARRY add_2296_23 (.CI(n29119), .I0(n2701), .I1(n80), .CO(n29120));
    SB_LUT4 add_2296_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n29118), 
            .O(n6156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1761_3_lut_3_lut (.I0(n2642), .I1(n6136), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4924), .I3(n30497), .O(n6_adj_4472)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n30497), .I0(GND_net), .I1(n6_adj_4924), 
            .CO(n30498));
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4925), .I3(n30496), .O(n7_adj_4471)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13159_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n35418), 
            .I3(GND_net), .O(n17904));   // verilog/coms.v(126[12] 289[6])
    defparam i13159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1762_3_lut_3_lut (.I0(n2642), .I1(n6137), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13160_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n35418), 
            .I3(GND_net), .O(n17905));   // verilog/coms.v(126[12] 289[6])
    defparam i13160_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_983_3 (.CI(n29662), .I0(n1458), .I1(GND_net), .CO(n29663));
    SB_CARRY add_2296_22 (.CI(n29118), .I0(n2702), .I1(n81), .CO(n29119));
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1558), .I1(VCC_net), 
            .CO(n29662));
    SB_LUT4 i13161_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n35418), 
            .I3(GND_net), .O(n17906));   // verilog/coms.v(126[12] 289[6])
    defparam i13161_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_2_add_3_19 (.CI(n29396), .I0(GND_net), .I1(n8_adj_4549), 
            .CO(n29397));
    SB_LUT4 i13162_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n35423), 
            .I3(GND_net), .O(n17907));   // verilog/coms.v(126[12] 289[6])
    defparam i13162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4550), .I3(n29395), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_18 (.CI(n29395), .I0(GND_net), .I1(n9_adj_4550), 
            .CO(n29396));
    SB_LUT4 i13163_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n35423), 
            .I3(GND_net), .O(n17908));   // verilog/coms.v(126[12] 289[6])
    defparam i13163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1050_14_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n29661), .O(n1646_adj_4462)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n30496), .I0(GND_net), .I1(n7_adj_4925), 
            .CO(n30497));
    SB_CARRY add_577_12 (.CI(n28671), .I0(n44224), .I1(n15_adj_4319), 
            .CO(n28672));
    SB_LUT4 rem_4_add_1050_13_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n29660), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_577_11_lut (.I0(duty[9]), .I1(n44224), .I2(n16_adj_4320), 
            .I3(n28670), .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4926), .I3(n30495), .O(n8_adj_4470)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4551), .I3(n29394), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_13 (.CI(n29660), .I0(n1548), .I1(VCC_net), 
            .CO(n29661));
    SB_LUT4 add_2296_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n29117), 
            .O(n6157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13164_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n35423), 
            .I3(GND_net), .O(n17909));   // verilog/coms.v(126[12] 289[6])
    defparam i13164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13165_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n35423), 
            .I3(GND_net), .O(n17910));   // verilog/coms.v(126[12] 289[6])
    defparam i13165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13166_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n35423), 
            .I3(GND_net), .O(n17911));   // verilog/coms.v(126[12] 289[6])
    defparam i13166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1759_3_lut_3_lut (.I0(n2642), .I1(n6134), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n29659), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_12 (.CI(n29659), .I0(n1549), .I1(VCC_net), 
            .CO(n29660));
    SB_LUT4 i13167_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n35423), 
            .I3(GND_net), .O(n17912));   // verilog/coms.v(126[12] 289[6])
    defparam i13167_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_2_add_3_17 (.CI(n29394), .I0(GND_net), .I1(n10_adj_4551), 
            .CO(n29395));
    SB_LUT4 i13168_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n35423), 
            .I3(GND_net), .O(n17913));   // verilog/coms.v(126[12] 289[6])
    defparam i13168_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_21 (.CI(n29117), .I0(n2703), .I1(n82), .CO(n29118));
    SB_LUT4 add_2296_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n29116), 
            .O(n6158)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13169_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n35423), 
            .I3(GND_net), .O(n17914));   // verilog/coms.v(126[12] 289[6])
    defparam i13169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4552), .I3(n29393), .O(n11_adj_4365)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n29658), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13170_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n35430), 
            .I3(GND_net), .O(n17915));   // verilog/coms.v(126[12] 289[6])
    defparam i13170_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_20 (.CI(n29116), .I0(n2704), .I1(n83), .CO(n29117));
    SB_LUT4 i13171_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n35430), 
            .I3(GND_net), .O(n17916));   // verilog/coms.v(126[12] 289[6])
    defparam i13171_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n30495), .I0(GND_net), .I1(n8_adj_4926), 
            .CO(n30496));
    SB_CARRY add_577_11 (.CI(n28670), .I0(n44224), .I1(n16_adj_4320), 
            .CO(n28671));
    SB_LUT4 i13172_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n35430), 
            .I3(GND_net), .O(n17917));   // verilog/coms.v(126[12] 289[6])
    defparam i13172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13173_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n35430), 
            .I3(GND_net), .O(n17918));   // verilog/coms.v(126[12] 289[6])
    defparam i13173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1760_3_lut_3_lut (.I0(n2642), .I1(n6135), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2296_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n29115), 
            .O(n6159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13174_3_lut (.I0(\data_in_frame[8] [4]), .I1(rx_data[4]), .I2(n35430), 
            .I3(GND_net), .O(n17919));   // verilog/coms.v(126[12] 289[6])
    defparam i13174_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_19 (.CI(n29115), .I0(n2705), .I1(n84), .CO(n29116));
    SB_LUT4 i13175_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n35430), 
            .I3(GND_net), .O(n17920));   // verilog/coms.v(126[12] 289[6])
    defparam i13175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2296_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n29114), 
            .O(n6160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_577_10_lut (.I0(duty[8]), .I1(n44224), .I2(n17_adj_4321), 
            .I3(n28669), .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13176_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n35430), 
            .I3(GND_net), .O(n17921));   // verilog/coms.v(126[12] 289[6])
    defparam i13176_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_18 (.CI(n29114), .I0(n2706), .I1(n85), .CO(n29115));
    SB_LUT4 i13177_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n35430), 
            .I3(GND_net), .O(n17922));   // verilog/coms.v(126[12] 289[6])
    defparam i13177_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_2_add_3_16 (.CI(n29393), .I0(GND_net), .I1(n11_adj_4552), 
            .CO(n29394));
    SB_LUT4 add_2296_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n29113), 
            .O(n6161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13121_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n35420), 
            .I3(GND_net), .O(n17866));   // verilog/coms.v(126[12] 289[6])
    defparam i13121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4553), .I3(n29392), .O(n12_adj_4342)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13122_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n35416), 
            .I3(GND_net), .O(n17867));   // verilog/coms.v(126[12] 289[6])
    defparam i13122_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_17 (.CI(n29113), .I0(n2707), .I1(n86), .CO(n29114));
    SB_LUT4 i13123_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n35416), 
            .I3(GND_net), .O(n17868));   // verilog/coms.v(126[12] 289[6])
    defparam i13123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13178_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n35429), 
            .I3(GND_net), .O(n17923));   // verilog/coms.v(126[12] 289[6])
    defparam i13178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13124_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n35416), 
            .I3(GND_net), .O(n17869));   // verilog/coms.v(126[12] 289[6])
    defparam i13124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13179_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n35429), 
            .I3(GND_net), .O(n17924));   // verilog/coms.v(126[12] 289[6])
    defparam i13179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13125_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n35416), 
            .I3(GND_net), .O(n17870));   // verilog/coms.v(126[12] 289[6])
    defparam i13125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1775_3_lut_3_lut (.I0(n2642), .I1(n6150), .I2(n530), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2296_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n29112), 
            .O(n6162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13126_3_lut (.I0(\data_in_frame[2] [4]), .I1(rx_data[4]), .I2(n35416), 
            .I3(GND_net), .O(n17871));   // verilog/coms.v(126[12] 289[6])
    defparam i13126_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_16 (.CI(n29112), .I0(n2708), .I1(n87), .CO(n29113));
    SB_LUT4 div_46_i1765_3_lut_3_lut (.I0(n2642), .I1(n6140), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_46_unary_minus_2_add_3_15 (.CI(n29392), .I0(GND_net), .I1(n12_adj_4553), 
            .CO(n29393));
    SB_LUT4 i13127_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n35416), 
            .I3(GND_net), .O(n17872));   // verilog/coms.v(126[12] 289[6])
    defparam i13127_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1050_11 (.CI(n29658), .I0(n1550), .I1(VCC_net), 
            .CO(n29659));
    SB_LUT4 add_2296_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n29111), 
            .O(n6163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13128_3_lut (.I0(\data_in_frame[2] [6]), .I1(rx_data[6]), .I2(n35416), 
            .I3(GND_net), .O(n17873));   // verilog/coms.v(126[12] 289[6])
    defparam i13128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13129_3_lut (.I0(\data_in_frame[2] [7]), .I1(rx_data[7]), .I2(n35416), 
            .I3(GND_net), .O(n17874));   // verilog/coms.v(126[12] 289[6])
    defparam i13129_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_577_10 (.CI(n28669), .I0(n44224), .I1(n17_adj_4321), 
            .CO(n28670));
    SB_LUT4 i13219_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n35434), .I3(GND_net), .O(n17964));   // verilog/coms.v(126[12] 289[6])
    defparam i13219_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_15 (.CI(n29111), .I0(n2709), .I1(n88), .CO(n29112));
    SB_LUT4 i13130_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n35417), 
            .I3(GND_net), .O(n17875));   // verilog/coms.v(126[12] 289[6])
    defparam i13130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13131_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n35417), 
            .I3(GND_net), .O(n17876));   // verilog/coms.v(126[12] 289[6])
    defparam i13131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1764_3_lut_3_lut (.I0(n2642), .I1(n6139), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2296_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n29110), 
            .O(n6164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4316));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n29657), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4554), .I3(n29391), .O(n13_adj_4344)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13132_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n35417), 
            .I3(GND_net), .O(n17877));   // verilog/coms.v(126[12] 289[6])
    defparam i13132_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_14 (.CI(n29110), .I0(n2710), .I1(n89), .CO(n29111));
    SB_LUT4 i13133_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n35417), 
            .I3(GND_net), .O(n17878));   // verilog/coms.v(126[12] 289[6])
    defparam i13133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13220_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n35434), .I3(GND_net), .O(n17965));   // verilog/coms.v(126[12] 289[6])
    defparam i13220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13134_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n35417), 
            .I3(GND_net), .O(n17879));   // verilog/coms.v(126[12] 289[6])
    defparam i13134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2296_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n29109), 
            .O(n6165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13135_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n35417), 
            .I3(GND_net), .O(n17880));   // verilog/coms.v(126[12] 289[6])
    defparam i13135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13136_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n35417), 
            .I3(GND_net), .O(n17881));   // verilog/coms.v(126[12] 289[6])
    defparam i13136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13137_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n35417), 
            .I3(GND_net), .O(n17882));   // verilog/coms.v(126[12] 289[6])
    defparam i13137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13138_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n35421), 
            .I3(GND_net), .O(n17883));   // verilog/coms.v(126[12] 289[6])
    defparam i13138_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_13 (.CI(n29109), .I0(n2711), .I1(n90), .CO(n29110));
    SB_LUT4 i13139_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n35421), 
            .I3(GND_net), .O(n17884));   // verilog/coms.v(126[12] 289[6])
    defparam i13139_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13140_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n35421), 
            .I3(GND_net), .O(n17885));   // verilog/coms.v(126[12] 289[6])
    defparam i13140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13141_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n35421), 
            .I3(GND_net), .O(n17886));   // verilog/coms.v(126[12] 289[6])
    defparam i13141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13142_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n35421), 
            .I3(GND_net), .O(n17887));   // verilog/coms.v(126[12] 289[6])
    defparam i13142_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2296_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n29108), 
            .O(n6166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13143_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n35421), 
            .I3(GND_net), .O(n17888));   // verilog/coms.v(126[12] 289[6])
    defparam i13143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13144_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n35421), 
            .I3(GND_net), .O(n17889));   // verilog/coms.v(126[12] 289[6])
    defparam i13144_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_12 (.CI(n29108), .I0(n2712), .I1(n91), .CO(n29109));
    SB_LUT4 div_46_i1773_3_lut_3_lut (.I0(n2642), .I1(n6148), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13145_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n35421), 
            .I3(GND_net), .O(n17890));   // verilog/coms.v(126[12] 289[6])
    defparam i13145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13300_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[5] [3]), 
            .I2(n17068), .I3(GND_net), .O(n18045));   // verilog/coms.v(126[12] 289[6])
    defparam i13300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13299_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[5] [2]), 
            .I2(n17068), .I3(GND_net), .O(n18044));   // verilog/coms.v(126[12] 289[6])
    defparam i13299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13298_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[5] [1]), 
            .I2(n17068), .I3(GND_net), .O(n18043));   // verilog/coms.v(126[12] 289[6])
    defparam i13298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13146_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n35422), 
            .I3(GND_net), .O(n17891));   // verilog/coms.v(126[12] 289[6])
    defparam i13146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2296_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n29107), 
            .O(n6167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13302_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[5] [5]), 
            .I2(n17068), .I3(GND_net), .O(n18047));   // verilog/coms.v(126[12] 289[6])
    defparam i13302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13301_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[5] [4]), 
            .I2(n17068), .I3(GND_net), .O(n18046));   // verilog/coms.v(126[12] 289[6])
    defparam i13301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13304_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[5] [7]), 
            .I2(n17068), .I3(GND_net), .O(n18049));   // verilog/coms.v(126[12] 289[6])
    defparam i13304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13303_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[5] [6]), 
            .I2(n17068), .I3(GND_net), .O(n18048));   // verilog/coms.v(126[12] 289[6])
    defparam i13303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13306_3_lut (.I0(encoder0_position[2]), .I1(n3020), .I2(count_enable), 
            .I3(GND_net), .O(n18051));   // quad.v(35[10] 41[6])
    defparam i13306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13305_3_lut (.I0(encoder0_position[1]), .I1(n3021), .I2(count_enable), 
            .I3(GND_net), .O(n18050));   // quad.v(35[10] 41[6])
    defparam i13305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4927), .I3(n30494), .O(n9_adj_4469)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13308_3_lut (.I0(encoder0_position[4]), .I1(n3018), .I2(count_enable), 
            .I3(GND_net), .O(n18053));   // quad.v(35[10] 41[6])
    defparam i13308_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_14 (.CI(n29391), .I0(GND_net), .I1(n13_adj_4554), 
            .CO(n29392));
    SB_CARRY add_2296_11 (.CI(n29107), .I0(n2713), .I1(n92), .CO(n29108));
    SB_LUT4 i13307_3_lut (.I0(encoder0_position[3]), .I1(n3019), .I2(count_enable), 
            .I3(GND_net), .O(n18052));   // quad.v(35[10] 41[6])
    defparam i13307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13310_3_lut (.I0(encoder0_position[6]), .I1(n3016), .I2(count_enable), 
            .I3(GND_net), .O(n18055));   // quad.v(35[10] 41[6])
    defparam i13310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13309_3_lut (.I0(encoder0_position[5]), .I1(n3017), .I2(count_enable), 
            .I3(GND_net), .O(n18054));   // quad.v(35[10] 41[6])
    defparam i13309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13147_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n35422), 
            .I3(GND_net), .O(n17892));   // verilog/coms.v(126[12] 289[6])
    defparam i13147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13148_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n35422), 
            .I3(GND_net), .O(n17893));   // verilog/coms.v(126[12] 289[6])
    defparam i13148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13149_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n35422), 
            .I3(GND_net), .O(n17894));   // verilog/coms.v(126[12] 289[6])
    defparam i13149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1774_3_lut_3_lut (.I0(n2642), .I1(n6149), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2296_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n29106), 
            .O(n6168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13221_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n35434), .I3(GND_net), .O(n17966));   // verilog/coms.v(126[12] 289[6])
    defparam i13221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13222_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n35434), .I3(GND_net), .O(n17967));   // verilog/coms.v(126[12] 289[6])
    defparam i13222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13223_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n35434), .I3(GND_net), .O(n17968));   // verilog/coms.v(126[12] 289[6])
    defparam i13223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13224_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n35434), .I3(GND_net), .O(n17969));   // verilog/coms.v(126[12] 289[6])
    defparam i13224_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2296_10 (.CI(n29106), .I0(n2714), .I1(n93), .CO(n29107));
    SB_LUT4 i13225_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n35434), .I3(GND_net), .O(n17970));   // verilog/coms.v(126[12] 289[6])
    defparam i13225_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13226_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n35435), .I3(GND_net), .O(n17971));   // verilog/coms.v(126[12] 289[6])
    defparam i13226_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13321_3_lut (.I0(encoder0_position[17]), .I1(n3005), .I2(count_enable), 
            .I3(GND_net), .O(n18066));   // quad.v(35[10] 41[6])
    defparam i13321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2296_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n29105), 
            .O(n6169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13320_3_lut (.I0(encoder0_position[16]), .I1(n3006), .I2(count_enable), 
            .I3(GND_net), .O(n18065));   // quad.v(35[10] 41[6])
    defparam i13320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13319_3_lut (.I0(encoder0_position[15]), .I1(n3007), .I2(count_enable), 
            .I3(GND_net), .O(n18064));   // quad.v(35[10] 41[6])
    defparam i13319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13318_3_lut (.I0(encoder0_position[14]), .I1(n3008), .I2(count_enable), 
            .I3(GND_net), .O(n18063));   // quad.v(35[10] 41[6])
    defparam i13318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13317_3_lut (.I0(encoder0_position[13]), .I1(n3009), .I2(count_enable), 
            .I3(GND_net), .O(n18062));   // quad.v(35[10] 41[6])
    defparam i13317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13316_3_lut (.I0(encoder0_position[12]), .I1(n3010), .I2(count_enable), 
            .I3(GND_net), .O(n18061));   // quad.v(35[10] 41[6])
    defparam i13316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13315_3_lut (.I0(encoder0_position[11]), .I1(n3011), .I2(count_enable), 
            .I3(GND_net), .O(n18060));   // quad.v(35[10] 41[6])
    defparam i13315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13314_3_lut (.I0(encoder0_position[10]), .I1(n3012), .I2(count_enable), 
            .I3(GND_net), .O(n18059));   // quad.v(35[10] 41[6])
    defparam i13314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13313_3_lut (.I0(encoder0_position[9]), .I1(n3013), .I2(count_enable), 
            .I3(GND_net), .O(n18058));   // quad.v(35[10] 41[6])
    defparam i13313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(n5_adj_4468), .I1(n122), .I2(n2778), 
            .I3(n63_adj_4399), .O(n6_adj_4872));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'heaaa;
    SB_LUT4 i2_3_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2388 ), .I2(n7_adj_4311), 
            .I3(GND_net), .O(n7_adj_4310));   // verilog/coms.v(126[12] 289[6])
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i4_4_lut_adj_1672 (.I0(n7_adj_4310), .I1(\FRAME_MATCHER.state_31__N_2586 [2]), 
            .I2(n6_adj_4872), .I3(n61_adj_4327), .O(n44421));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1672.LUT_INIT = 16'hfafe;
    SB_LUT4 div_46_i1766_3_lut_3_lut (.I0(n2642), .I1(n6141), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1050_10 (.CI(n29657), .I0(n1551), .I1(VCC_net), 
            .CO(n29658));
    SB_LUT4 div_46_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4555), .I3(n29390), .O(n14_adj_4334)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n29656), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1767_3_lut_3_lut (.I0(n2642), .I1(n6142), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_46_unary_minus_2_add_3_13 (.CI(n29390), .I0(GND_net), .I1(n14_adj_4555), 
            .CO(n29391));
    SB_LUT4 div_46_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4556), .I3(n29389), .O(n15_adj_4361)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_9 (.CI(n29656), .I0(n1552), .I1(VCC_net), 
            .CO(n29657));
    SB_LUT4 div_46_i1772_3_lut_3_lut (.I0(n2642), .I1(n6147), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_46_unary_minus_2_add_3_12 (.CI(n29389), .I0(GND_net), .I1(n15_adj_4556), 
            .CO(n29390));
    SB_LUT4 div_46_i1770_3_lut_3_lut (.I0(n2642), .I1(n6145), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4557), .I3(n29388), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1553_adj_4487), .I2(VCC_net), 
            .I3(n29655), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n30494), .I0(GND_net), .I1(n9_adj_4927), 
            .CO(n30495));
    SB_CARRY rem_4_add_1050_8 (.CI(n29655), .I0(n1553_adj_4487), .I1(VCC_net), 
            .CO(n29656));
    SB_LUT4 div_46_i1769_3_lut_3_lut (.I0(n2642), .I1(n6144), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1554_adj_4488), .I2(GND_net), 
            .I3(n29654), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_11 (.CI(n29388), .I0(GND_net), .I1(n16_adj_4557), 
            .CO(n29389));
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n16_adj_4979), .I1(n2778), .I2(n61_adj_4327), 
            .I3(n3741), .O(n5_adj_4326));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'heeef;
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4928), .I3(n30493), .O(n10_adj_4433)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut_adj_1674 (.I0(n29), .I1(n31_adj_4411), .I2(n30), 
            .I3(n32), .O(n2570));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i17_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1050_7 (.CI(n29654), .I0(n1554_adj_4488), .I1(GND_net), 
            .CO(n29655));
    SB_LUT4 div_46_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4558), .I3(n29387), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n29653), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_10 (.CI(n29387), .I0(GND_net), .I1(n17_adj_4558), 
            .CO(n29388));
    SB_LUT4 div_46_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4559), .I3(n29386), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_9 (.CI(n29105), .I0(n2715), .I1(n94), .CO(n29106));
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_577_9_lut (.I0(duty[7]), .I1(n44224), .I2(n18_adj_4322), 
            .I3(n28668), .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4315));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4314));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1763_3_lut_3_lut (.I0(n2642), .I1(n6138), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12976_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13293), .I3(GND_net), .O(n17721));   // verilog/coms.v(126[12] 289[6])
    defparam i12976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4431), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12977_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13293), .I3(GND_net), .O(n17722));   // verilog/coms.v(126[12] 289[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12978_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13293), .I3(GND_net), .O(n17723));   // verilog/coms.v(126[12] 289[6])
    defparam i12978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12979_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13293), .I3(GND_net), .O(n17724));   // verilog/coms.v(126[12] 289[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12980_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13293), .I3(GND_net), .O(n17725));   // verilog/coms.v(126[12] 289[6])
    defparam i12980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12981_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13293), .I3(GND_net), .O(n17726));   // verilog/coms.v(126[12] 289[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12982_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13293), .I3(GND_net), .O(n17727));   // verilog/coms.v(126[12] 289[6])
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12983_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13293), .I3(GND_net), .O(n17728));   // verilog/coms.v(126[12] 289[6])
    defparam i12983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12984_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13293), .I3(GND_net), .O(n17729));   // verilog/coms.v(126[12] 289[6])
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12985_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13293), .I3(GND_net), .O(n17730));   // verilog/coms.v(126[12] 289[6])
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1771_3_lut_3_lut (.I0(n2642), .I1(n6146), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12986_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13293), .I3(GND_net), .O(n17731));   // verilog/coms.v(126[12] 289[6])
    defparam i12986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12987_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13293), .I3(GND_net), .O(n17732));   // verilog/coms.v(126[12] 289[6])
    defparam i12987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12988_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13293), .I3(GND_net), .O(n17733));   // verilog/coms.v(126[12] 289[6])
    defparam i12988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12989_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13293), .I3(GND_net), .O(n17734));   // verilog/coms.v(126[12] 289[6])
    defparam i12989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12990_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13293), .I3(GND_net), .O(n17735));   // verilog/coms.v(126[12] 289[6])
    defparam i12990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12991_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13293), .I3(GND_net), .O(n17736));   // verilog/coms.v(126[12] 289[6])
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12992_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13293), .I3(GND_net), .O(n17737));   // verilog/coms.v(126[12] 289[6])
    defparam i12992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12993_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13293), .I3(GND_net), .O(n17738));   // verilog/coms.v(126[12] 289[6])
    defparam i12993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12994_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13293), .I3(GND_net), .O(n17739));   // verilog/coms.v(126[12] 289[6])
    defparam i12994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12995_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13293), .I3(GND_net), .O(n17740));   // verilog/coms.v(126[12] 289[6])
    defparam i12995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12996_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13293), .I3(GND_net), .O(n17741));   // verilog/coms.v(126[12] 289[6])
    defparam i12996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12997_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13293), .I3(GND_net), .O(n17742));   // verilog/coms.v(126[12] 289[6])
    defparam i12997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12998_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13293), .I3(GND_net), .O(n17743));   // verilog/coms.v(126[12] 289[6])
    defparam i12998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12999_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13293), .I3(GND_net), .O(n17744));   // verilog/coms.v(126[12] 289[6])
    defparam i12999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13000_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13293), .I3(GND_net), .O(n17745));   // verilog/coms.v(126[12] 289[6])
    defparam i13000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13001_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13293), .I3(GND_net), .O(n17746));   // verilog/coms.v(126[12] 289[6])
    defparam i13001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13002_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13293), .I3(GND_net), .O(n17747));   // verilog/coms.v(126[12] 289[6])
    defparam i13002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13003_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13293), .I3(GND_net), .O(n17748));   // verilog/coms.v(126[12] 289[6])
    defparam i13003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13004_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13293), .I3(GND_net), .O(n17749));   // verilog/coms.v(126[12] 289[6])
    defparam i13004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13005_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13293), .I3(GND_net), .O(n17750));   // verilog/coms.v(126[12] 289[6])
    defparam i13005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13006_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13293), .I3(GND_net), .O(n17751));   // verilog/coms.v(126[12] 289[6])
    defparam i13006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13007_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13293), .I3(GND_net), .O(n17752));   // verilog/coms.v(126[12] 289[6])
    defparam i13007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4922));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13008_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13293), .I3(GND_net), .O(n17753));   // verilog/coms.v(126[12] 289[6])
    defparam i13008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4547));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6156), 
            .I3(n2724), .O(n41_adj_4866));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6157), 
            .I3(n2724), .O(n39_adj_4865));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4340), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n532));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(\FRAME_MATCHER.i_31__N_2390 ), .I1(n63_adj_4399), 
            .I2(n2855), .I3(n123), .O(n4_adj_4981));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'haaa2;
    SB_LUT4 div_46_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6154), 
            .I3(n2724), .O(n45_adj_4868));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6155), 
            .I3(n2724), .O(n43_adj_4867));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n4_adj_4981), .I1(n123), .I2(n5_adj_4326), 
            .I3(n63_adj_4399), .O(n5_adj_4980));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'heafa;
    SB_LUT4 div_46_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6162), 
            .I3(n2724), .O(n29_adj_4859));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i3_4_lut_adj_1677 (.I0(n5_adj_4980), .I1(\FRAME_MATCHER.state_31__N_2458 [1]), 
            .I2(\FRAME_MATCHER.i_31__N_2388 ), .I3(n97_adj_4328), .O(n44420));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1677.LUT_INIT = 16'hfafe;
    SB_LUT4 div_46_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6161), 
            .I3(n2724), .O(n31_adj_4861));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6158), 
            .I3(n2724), .O(n37_adj_4864));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i23748_2_lut_3_lut (.I0(n28152), .I1(n746), .I2(n855), .I3(GND_net), 
            .O(n957));
    defparam i23748_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 div_46_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6166), 
            .I3(n2724), .O(n21_adj_4854));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13339_3_lut (.I0(encoder1_position[10]), .I1(n2962), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18084));   // quad.v(35[10] 41[6])
    defparam i13339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6165), 
            .I3(n2724), .O(n23_adj_4855));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6164), 
            .I3(n2724), .O(n25_adj_4857));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13338_3_lut (.I0(encoder1_position[9]), .I1(n2963), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18083));   // quad.v(35[10] 41[6])
    defparam i13338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6168), 
            .I3(n2724), .O(n17_adj_4852));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6167), 
            .I3(n2724), .O(n19_adj_4853));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6172), 
            .I3(n2724), .O(n9_adj_4845));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6173), 
            .I3(n2724), .O(n7_adj_4843));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6159), 
            .I3(n2724), .O(n35_adj_4863));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6160), 
            .I3(n2724), .O(n33_adj_4862));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13337_3_lut (.I0(encoder1_position[8]), .I1(n2964), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18082));   // quad.v(35[10] 41[6])
    defparam i13337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6171), 
            .I3(n2724), .O(n11_adj_4847));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6170), 
            .I3(n2724), .O(n13_adj_4849));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13150_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n35422), 
            .I3(GND_net), .O(n17895));   // verilog/coms.v(126[12] 289[6])
    defparam i13150_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6169), 
            .I3(n2724), .O(n15_adj_4850));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6163), 
            .I3(n2724), .O(n27_adj_4858));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13341_3_lut (.I0(encoder1_position[12]), .I1(n2960), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18086));   // quad.v(35[10] 41[6])
    defparam i13341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34990_4_lut (.I0(n27_adj_4858), .I1(n15_adj_4850), .I2(n13_adj_4849), 
            .I3(n11_adj_4847), .O(n41844));
    defparam i34990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4862), 
            .I3(GND_net), .O(n12_adj_4848));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13340_3_lut (.I0(encoder1_position[11]), .I1(n2961), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18085));   // quad.v(35[10] 41[6])
    defparam i13340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n28152), .I1(n746), .I2(n4_adj_4396), 
            .I3(n748), .O(n955));
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 rem_4_i586_3_lut_4_lut (.I0(n28152), .I1(n746), .I2(n855), 
            .I3(n749), .O(n956));
    defparam rem_4_i586_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 i13291_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[6] [2]), 
            .I2(n17068), .I3(GND_net), .O(n18036));   // verilog/coms.v(126[12] 289[6])
    defparam i13291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4424), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4425), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4423), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2357_adj_4579));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4421), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458_adj_4516));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357_adj_4579), .I1(n2424), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2456_adj_4518));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4472), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34964_2_lut (.I0(n33_adj_4862), .I1(n15_adj_4850), .I2(GND_net), 
            .I3(GND_net), .O(n41818));
    defparam i34964_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13343_3_lut (.I0(encoder1_position[14]), .I1(n2958), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18088));   // quad.v(35[10] 41[6])
    defparam i13343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4849), 
            .I3(GND_net), .O(n10_adj_4846));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i30_3_lut (.I0(n12_adj_4848), .I1(n83), 
            .I2(n35_adj_4863), .I3(GND_net), .O(n30_adj_4860));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13342_3_lut (.I0(encoder1_position[13]), .I1(n2959), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18087));   // quad.v(35[10] 41[6])
    defparam i13342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13345_3_lut (.I0(encoder1_position[16]), .I1(n2956), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18090));   // quad.v(35[10] 41[6])
    defparam i13345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13344_3_lut (.I0(encoder1_position[15]), .I1(n2957), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18089));   // quad.v(35[10] 41[6])
    defparam i13344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1828_3_lut (.I0(n2720), .I1(n6174), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35061_3_lut (.I0(n7_adj_4843), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n41915));
    defparam i35061_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420_adj_4496), .I2(n1382), 
            .I3(GND_net), .O(n1452));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650_adj_4466));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650_adj_4466), .I1(n1717), .I2(n1679), 
            .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1257_3_lut (.I0(n1848), .I1(n1915), .I2(n1877), .I3(GND_net), 
            .O(n1947));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4471), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i722_rep_77_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), 
            .I3(GND_net), .O(n1156));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i722_rep_77_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i990_rep_70_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), 
            .I3(GND_net), .O(n1552));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i990_rep_70_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651_adj_4467));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651_adj_4467), .I1(n1718), .I2(n1679), 
            .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1258_3_lut (.I0(n1849), .I1(n1916), .I2(n1877), .I3(GND_net), 
            .O(n1948));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13347_3_lut (.I0(encoder1_position[18]), .I1(n2954), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18092));   // quad.v(35[10] 41[6])
    defparam i13347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35697_4_lut (.I0(n13_adj_4849), .I1(n11_adj_4847), .I2(n9_adj_4845), 
            .I3(n41915), .O(n42551));
    defparam i35697_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35681_4_lut (.I0(n19_adj_4853), .I1(n17_adj_4852), .I2(n15_adj_4850), 
            .I3(n42551), .O(n42535));
    defparam i35681_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i13346_3_lut (.I0(encoder1_position[17]), .I1(n2955), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18091));   // quad.v(35[10] 41[6])
    defparam i13346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36408_4_lut (.I0(n25_adj_4857), .I1(n23_adj_4855), .I2(n21_adj_4854), 
            .I3(n42535), .O(n43262));
    defparam i36408_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35976_4_lut (.I0(n31_adj_4861), .I1(n29_adj_4859), .I2(n27_adj_4858), 
            .I3(n43262), .O(n42830));
    defparam i35976_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4430), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756_adj_4456));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756_adj_4456), .I1(n1823), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1264_3_lut (.I0(n1855), .I1(n1922), .I2(n1877), .I3(GND_net), 
            .O(n1954));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1398_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1602_3_lut (.I0(n2353), .I1(n2420), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2452_adj_4570));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35385_3_lut (.I0(n2250), .I1(n2317), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35386_3_lut (.I0(n2349), .I1(n2416), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2448_adj_4574));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1597_3_lut (.I0(n2348), .I1(n2415), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2447_adj_4575));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36091_3_lut (.I0(n2251), .I1(n2318), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2350));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35875_3_lut (.I0(n2350), .I1(n2417), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2449_adj_4573));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35551_3_lut (.I0(n1877), .I1(n1778_adj_4818), .I2(n1679), 
            .I3(GND_net), .O(n42405));
    defparam i35551_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1059_3_lut (.I0(n1554_adj_4488), .I1(n1621), .I2(n1580), 
            .I3(GND_net), .O(n1653_adj_4460));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1126_rep_59_3_lut (.I0(n1720), .I1(n1819), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n39157));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1126_rep_59_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1193_rep_53_3_lut (.I0(n39157), .I1(n1918), .I2(n1877), 
            .I3(GND_net), .O(n39151));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1193_rep_53_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36179_3_lut (.I0(n39151), .I1(n1653_adj_4460), .I2(n42405), 
            .I3(GND_net), .O(n1950));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13349_3_lut (.I0(encoder1_position[20]), .I1(n2952), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18094));   // quad.v(35[10] 41[6])
    defparam i13349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36510_4_lut (.I0(n37_adj_4864), .I1(n35_adj_4863), .I2(n33_adj_4862), 
            .I3(n42830), .O(n43364));
    defparam i36510_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13348_3_lut (.I0(encoder1_position[19]), .I1(n2953), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18093));   // quad.v(35[10] 41[6])
    defparam i13348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4867), 
            .I3(GND_net), .O(n16_adj_4851));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13151_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n35422), 
            .I3(GND_net), .O(n17896));   // verilog/coms.v(126[12] 289[6])
    defparam i13151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4843), 
            .I3(GND_net), .O(n6_adj_4842));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i36180_3_lut (.I0(n1950), .I1(n2017), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36186_3_lut (.I0(n1652_adj_4459), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1192_3_lut (.I0(n1751), .I1(n1818), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1259_3_lut (.I0(n1850), .I1(n1917), .I2(n1877), .I3(GND_net), 
            .O(n1949));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2346));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4475), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1678 (.I0(n957), .I1(n956), .I2(n958), .I3(GND_net), 
            .O(n36409));
    defparam i1_3_lut_adj_1678.LUT_INIT = 16'hfefe;
    SB_LUT4 i20977_4_lut (.I0(n954), .I1(n953), .I2(n36409), .I3(n955), 
            .O(n986));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i20977_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_1679 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n36407));
    defparam i1_3_lut_adj_1679.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1680 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n38491));
    defparam i1_2_lut_adj_1680.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n1052), .I1(n38491), .I2(n1053), .I3(n36407), 
            .O(n1085));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'hfefa;
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1682 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n38495));
    defparam i1_2_lut_adj_1682.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(n1154), .I1(n38495), .I2(n1155), .I3(n1157), 
            .O(n36403));
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'ha080;
    SB_LUT4 i36058_3_lut (.I0(n6_adj_4842), .I1(n90), .I2(n21_adj_4854), 
            .I3(GND_net), .O(n42912));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36058_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36059_3_lut (.I0(n42912), .I1(n89), .I2(n23_adj_4855), .I3(GND_net), 
            .O(n42913));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36059_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35018_4_lut (.I0(n21_adj_4854), .I1(n19_adj_4853), .I2(n17_adj_4852), 
            .I3(n9_adj_4845), .O(n41872));
    defparam i35018_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1050_6 (.CI(n29653), .I0(n1555), .I1(GND_net), 
            .CO(n29654));
    SB_LUT4 i34885_2_lut (.I0(n43_adj_4867), .I1(n19_adj_4853), .I2(GND_net), 
            .I3(GND_net), .O(n41739));
    defparam i34885_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13152_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n35422), 
            .I3(GND_net), .O(n17897));   // verilog/coms.v(126[12] 289[6])
    defparam i13152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n29652), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n30493), .I0(GND_net), .I1(n10_adj_4928), 
            .CO(n30494));
    SB_CARRY add_577_9 (.CI(n28668), .I0(n44224), .I1(n18_adj_4322), .CO(n28669));
    SB_CARRY rem_4_add_1050_5 (.CI(n29652), .I0(n1556), .I1(VCC_net), 
            .CO(n29653));
    SB_LUT4 div_46_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4852), 
            .I3(GND_net), .O(n8_adj_4844));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i24_3_lut (.I0(n16_adj_4851), .I1(n78), 
            .I2(n45_adj_4868), .I3(GND_net), .O(n24_adj_4856));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34893_4_lut (.I0(n43_adj_4867), .I1(n25_adj_4857), .I2(n23_adj_4855), 
            .I3(n41872), .O(n41747));
    defparam i34893_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35890_4_lut (.I0(n24_adj_4856), .I1(n8_adj_4844), .I2(n45_adj_4868), 
            .I3(n41739), .O(n42744));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35890_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4929), .I3(n30492), .O(n11_adj_4432)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n29651), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35468_3_lut (.I0(n42913), .I1(n88), .I2(n25_adj_4857), .I3(GND_net), 
            .O(n42322));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35468_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1829_3_lut (.I0(n531), .I1(n6175), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13153_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n35422), 
            .I3(GND_net), .O(n17898));   // verilog/coms.v(126[12] 289[6])
    defparam i13153_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1050_4 (.CI(n29651), .I0(n1557), .I1(VCC_net), 
            .CO(n29652));
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(n29650), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_9 (.CI(n29386), .I0(GND_net), .I1(n18_adj_4559), 
            .CO(n29387));
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n30492), .I0(GND_net), .I1(n11_adj_4929), 
            .CO(n30493));
    SB_CARRY rem_4_add_1050_3 (.CI(n29650), .I0(n1558), .I1(GND_net), 
            .CO(n29651));
    SB_LUT4 div_46_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4560), .I3(n29385), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n29104), 
            .O(n6170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1658), .I1(VCC_net), 
            .CO(n29650));
    SB_CARRY div_46_unary_minus_2_add_3_8 (.CI(n29385), .I0(GND_net), .I1(n19_adj_4560), 
            .CO(n29386));
    SB_LUT4 div_46_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4561), .I3(n29384), .O(n20_adj_4335)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_8 (.CI(n29104), .I0(n2716), .I1(n95), .CO(n29105));
    SB_LUT4 add_577_8_lut (.I0(duty[6]), .I1(n44224), .I2(n19_adj_4323), 
            .I3(n28667), .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_LessThan_1830_i4_4_lut (.I0(n532), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4841));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_2296_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n29103), 
            .O(n6171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4930), .I3(n30491), .O(n12_adj_4431)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_7 (.CI(n29103), .I0(n2717), .I1(n96), .CO(n29104));
    SB_CARRY div_46_unary_minus_2_add_3_7 (.CI(n29384), .I0(GND_net), .I1(n20_adj_4561), 
            .CO(n29385));
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4462), .I2(VCC_net), 
            .I3(n29649), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n30491), .I0(GND_net), .I1(n12_adj_4930), 
            .CO(n30492));
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4931), .I3(n30490), .O(n13_adj_4430)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4463), .I2(VCC_net), 
            .I3(n29648), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_14 (.CI(n29648), .I0(n1647_adj_4463), .I1(VCC_net), 
            .CO(n29649));
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n30490), .I0(GND_net), .I1(n13_adj_4931), 
            .CO(n30491));
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4932), .I3(n30489), .O(n14_adj_4429)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13352_3_lut (.I0(encoder1_position[23]), .I1(n2949), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18097));   // quad.v(35[10] 41[6])
    defparam i13352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36093_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35873_3_lut (.I0(n2351), .I1(n2418), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2450_adj_4572));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647_adj_4463));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2453_adj_4569));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36056_3_lut (.I0(n4_adj_4841), .I1(n87), .I2(n27_adj_4858), 
            .I3(GND_net), .O(n42910));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36056_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36057_3_lut (.I0(n42910), .I1(n86), .I2(n29_adj_4859), .I3(GND_net), 
            .O(n42911));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36057_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13351_3_lut (.I0(encoder1_position[22]), .I1(n2950), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18096));   // quad.v(35[10] 41[6])
    defparam i13351_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n30489), .I0(GND_net), .I1(n14_adj_4932), 
            .CO(n30490));
    SB_LUT4 i34972_4_lut (.I0(n33_adj_4862), .I1(n31_adj_4861), .I2(n29_adj_4859), 
            .I3(n41844), .O(n41826));
    defparam i34972_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36472_4_lut (.I0(n30_adj_4860), .I1(n10_adj_4846), .I2(n35_adj_4863), 
            .I3(n41818), .O(n43326));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36472_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4464), .I2(VCC_net), 
            .I3(n29647), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13350_3_lut (.I0(encoder1_position[21]), .I1(n2951), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18095));   // quad.v(35[10] 41[6])
    defparam i13350_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_13 (.CI(n29647), .I0(n1648_adj_4464), .I1(VCC_net), 
            .CO(n29648));
    SB_LUT4 i13297_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[5] [0]), 
            .I2(n17068), .I3(GND_net), .O(n18042));   // verilog/coms.v(126[12] 289[6])
    defparam i13297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4465), .I2(VCC_net), 
            .I3(n29646), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4562), .I3(n29383), .O(n21_adj_4336)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4933), .I3(n30488), .O(n15_adj_4428)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_12 (.CI(n29646), .I0(n1649_adj_4465), .I1(VCC_net), 
            .CO(n29647));
    SB_CARRY div_46_unary_minus_2_add_3_6 (.CI(n29383), .I0(GND_net), .I1(n21_adj_4562), 
            .CO(n29384));
    SB_LUT4 add_2296_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n29102), 
            .O(n6172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4466), .I2(VCC_net), 
            .I3(n29645), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4563), .I3(n29382), .O(n22_adj_4337)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_11 (.CI(n29645), .I0(n1650_adj_4466), .I1(VCC_net), 
            .CO(n29646));
    SB_CARRY div_46_unary_minus_2_add_3_5 (.CI(n29382), .I0(GND_net), .I1(n22_adj_4563), 
            .CO(n29383));
    SB_CARRY add_2296_6 (.CI(n29102), .I0(n2718), .I1(n97), .CO(n29103));
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n30488), .I0(GND_net), .I1(n15_adj_4933), 
            .CO(n30489));
    SB_LUT4 i13296_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[6] [7]), 
            .I2(n17068), .I3(GND_net), .O(n18041));   // verilog/coms.v(126[12] 289[6])
    defparam i13296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35470_3_lut (.I0(n42911), .I1(n85), .I2(n31_adj_4861), .I3(GND_net), 
            .O(n42324));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35470_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36582_4_lut (.I0(n42324), .I1(n43326), .I2(n35_adj_4863), 
            .I3(n41826), .O(n43436));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36582_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4467), .I2(VCC_net), 
            .I3(n29644), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_10 (.CI(n29644), .I0(n1651_adj_4467), .I1(VCC_net), 
            .CO(n29645));
    SB_LUT4 add_2296_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n29101), 
            .O(n6173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_5 (.CI(n29101), .I0(n2719), .I1(n98), .CO(n29102));
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4459), .I2(VCC_net), 
            .I3(n29643), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_8 (.CI(n28667), .I0(n44224), .I1(n19_adj_4323), .CO(n28668));
    SB_LUT4 div_46_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4564), .I3(n29381), .O(n23_adj_4338)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_4 (.CI(n29381), .I0(GND_net), .I1(n23_adj_4564), 
            .CO(n29382));
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4934), .I3(n30487), .O(n16_adj_4427)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n30487), .I0(GND_net), .I1(n16_adj_4934), 
            .CO(n30488));
    SB_LUT4 add_2296_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n29100), 
            .O(n6174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36583_3_lut (.I0(n43436), .I1(n82), .I2(n37_adj_4864), .I3(GND_net), 
            .O(n43437));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36583_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36542_3_lut (.I0(n43437), .I1(n81), .I2(n39_adj_4865), .I3(GND_net), 
            .O(n43396));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36542_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34940_4_lut (.I0(n43_adj_4867), .I1(n41_adj_4866), .I2(n39_adj_4865), 
            .I3(n43364), .O(n41794));
    defparam i34940_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36376_4_lut (.I0(n42322), .I1(n42744), .I2(n45_adj_4868), 
            .I3(n41747), .O(n43230));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36376_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13295_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[6] [6]), 
            .I2(n17068), .I3(GND_net), .O(n18040));   // verilog/coms.v(126[12] 289[6])
    defparam i13295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35476_3_lut (.I0(n43396), .I1(n80), .I2(n41_adj_4866), .I3(GND_net), 
            .O(n42330));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35476_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_577_7_lut (.I0(duty[5]), .I1(n44224), .I2(n20), .I3(n28666), 
            .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1117_9 (.CI(n29643), .I0(n1652_adj_4459), .I1(VCC_net), 
            .CO(n29644));
    SB_CARRY add_2296_4 (.CI(n29100), .I0(n2720), .I1(n99), .CO(n29101));
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4460), .I2(VCC_net), 
            .I3(n29642), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_3_lut (.I0(GND_net), .I1(n531), .I2(n558), .I3(n29099), 
            .O(n6175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4565), .I3(n29380), .O(n24_adj_4339)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_7 (.CI(n28666), .I0(n44224), .I1(n20), .CO(n28667));
    SB_LUT4 rem_4_i584_3_lut_4_lut (.I0(n28152), .I1(n746), .I2(n6_adj_4343), 
            .I3(n852), .O(n954));
    defparam rem_4_i584_3_lut_4_lut.LUT_INIT = 16'h7f08;
    SB_LUT4 i13294_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[6] [5]), 
            .I2(n17068), .I3(GND_net), .O(n18039));   // verilog/coms.v(126[12] 289[6])
    defparam i13294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13293_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[6] [4]), 
            .I2(n17068), .I3(GND_net), .O(n18038));   // verilog/coms.v(126[12] 289[6])
    defparam i13293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1807_3_lut (.I0(n2699), .I1(n6153), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_8 (.CI(n29642), .I0(n1653_adj_4460), .I1(VCC_net), 
            .CO(n29643));
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n29641), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_3 (.CI(n29380), .I0(GND_net), .I1(n24_adj_4565), 
            .CO(n29381));
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4935), .I3(n30486), .O(n17_adj_4426)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_7 (.CI(n29641), .I0(n1654), .I1(GND_net), 
            .CO(n29642));
    SB_LUT4 div_46_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4566), .I3(VCC_net), .O(n25_adj_4340)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_3 (.CI(n29099), .I0(n531), .I1(n558), .CO(n29100));
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n29640), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4566), 
            .CO(n29380));
    SB_CARRY rem_4_add_1117_6 (.CI(n29640), .I0(n1655), .I1(GND_net), 
            .CO(n29641));
    SB_LUT4 div_46_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4519), .I3(n29379), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2296_2 (.CI(VCC_net), .I0(n532), .I1(VCC_net), .CO(n29099));
    SB_LUT4 add_577_6_lut (.I0(duty[4]), .I1(n44224), .I2(n21), .I3(n28665), 
            .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n29639), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4520), .I3(n29378), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_6 (.CI(n28665), .I0(n44224), .I1(n21), .CO(n28666));
    SB_LUT4 rem_4_add_916_11_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n28549), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n30486), .I0(GND_net), .I1(n17_adj_4935), 
            .CO(n30487));
    SB_CARRY rem_4_add_1117_5 (.CI(n29639), .I0(n1656), .I1(VCC_net), 
            .CO(n29640));
    SB_CARRY div_46_unary_minus_4_add_3_24 (.CI(n29378), .I0(GND_net), .I1(n3_adj_4520), 
            .CO(n29379));
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n29638), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_4 (.CI(n29638), .I0(n1657), .I1(VCC_net), 
            .CO(n29639));
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n29637), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4521), .I3(n29377), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2295_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n29098), 
            .O(n6129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_23 (.CI(n29377), .I0(GND_net), .I1(n4_adj_4521), 
            .CO(n29378));
    SB_LUT4 add_2295_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n29097), 
            .O(n6130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4936), .I3(n30485), .O(n18_adj_4425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_3 (.CI(n29637), .I0(n1658), .I1(GND_net), 
            .CO(n29638));
    SB_LUT4 div_46_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4522), .I3(n29376), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_22 (.CI(n29097), .I0(n2619), .I1(n80), .CO(n29098));
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n28548), .O(n1417_adj_4493)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4458), .I1(VCC_net), 
            .CO(n29637));
    SB_CARRY div_46_unary_minus_4_add_3_22 (.CI(n29376), .I0(GND_net), .I1(n5_adj_4522), 
            .CO(n29377));
    SB_LUT4 rem_4_add_1184_16_lut (.I0(n1778_adj_4818), .I1(n1745), .I2(VCC_net), 
            .I3(n29636), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4523), .I3(n29375), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_15_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n29635), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_21 (.CI(n29375), .I0(GND_net), .I1(n6_adj_4523), 
            .CO(n29376));
    SB_LUT4 add_2295_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n29096), 
            .O(n6131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_577_5_lut (.I0(duty[3]), .I1(n44224), .I2(n22), .I3(n28664), 
            .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2295_21 (.CI(n29096), .I0(n2620), .I1(n81), .CO(n29097));
    SB_LUT4 add_2295_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n29095), 
            .O(n6132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36504_4_lut (.I0(n42330), .I1(n43230), .I2(n45_adj_4868), 
            .I3(n41794), .O(n43358));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36504_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2295_20 (.CI(n29095), .I0(n2621), .I1(n82), .CO(n29096));
    SB_LUT4 add_2295_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n29094), 
            .O(n6133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_19 (.CI(n29094), .I0(n2622), .I1(n83), .CO(n29095));
    SB_LUT4 add_2295_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n29093), 
            .O(n6134)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_18 (.CI(n29093), .I0(n2623), .I1(n84), .CO(n29094));
    SB_LUT4 add_2295_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n29092), 
            .O(n6135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_17 (.CI(n29092), .I0(n2624), .I1(n85), .CO(n29093));
    SB_LUT4 add_2295_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n29091), 
            .O(n6136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_16 (.CI(n29091), .I0(n2625), .I1(n86), .CO(n29092));
    SB_CARRY rem_4_add_916_10 (.CI(n28548), .I0(n1350), .I1(VCC_net), 
            .CO(n28549));
    SB_LUT4 add_2295_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n29090), 
            .O(n6137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36505_3_lut (.I0(n43358), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36505_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n30485), .I0(GND_net), .I1(n18_adj_4936), 
            .CO(n30486));
    SB_CARRY rem_4_add_1184_15 (.CI(n29635), .I0(n1746), .I1(VCC_net), 
            .CO(n29636));
    SB_LUT4 div_46_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4524), .I3(n29374), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n29634), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_20 (.CI(n29374), .I0(GND_net), .I1(n7_adj_4524), 
            .CO(n29375));
    SB_CARRY add_2295_15 (.CI(n29090), .I0(n2626), .I1(n87), .CO(n29091));
    SB_LUT4 div_46_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4525), .I3(n29373), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n29634), .I0(n1747), .I1(VCC_net), 
            .CO(n29635));
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4937), .I3(n30484), .O(n19_adj_4424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n29633), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_19 (.CI(n29373), .I0(GND_net), .I1(n8_adj_4525), 
            .CO(n29374));
    SB_CARRY rem_4_add_1184_13 (.CI(n29633), .I0(n1748), .I1(VCC_net), 
            .CO(n29634));
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n29632), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4526), .I3(n29372), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2295_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n29089), 
            .O(n6138)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_18 (.CI(n29372), .I0(GND_net), .I1(n9_adj_4526), 
            .CO(n29373));
    SB_CARRY rem_4_add_1184_12 (.CI(n29632), .I0(n1749), .I1(VCC_net), 
            .CO(n29633));
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n30484), .I0(GND_net), .I1(n19_adj_4937), 
            .CO(n30485));
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n29631), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4938), .I3(n30483), .O(n20_adj_4423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4432), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4546));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4433), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_11 (.CI(n29631), .I0(n1750), .I1(VCC_net), 
            .CO(n29632));
    SB_LUT4 div_46_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4527), .I3(n29371), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n30483), .I0(GND_net), .I1(n20_adj_4938), 
            .CO(n30484));
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4939), .I3(n30482), .O(n21_adj_4422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_14 (.CI(n29089), .I0(n2627), .I1(n88), .CO(n29090));
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n28547), .O(n1418_adj_4494)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2295_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n29088), 
            .O(n6139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_17 (.CI(n29371), .I0(GND_net), .I1(n10_adj_4527), 
            .CO(n29372));
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n29630), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2295_13 (.CI(n29088), .I0(n2628), .I1(n89), .CO(n29089));
    SB_LUT4 div_46_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4528), .I3(n29370), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_16 (.CI(n29370), .I0(GND_net), .I1(n11_adj_4528), 
            .CO(n29371));
    SB_CARRY rem_4_add_1184_10 (.CI(n29630), .I0(n1751), .I1(VCC_net), 
            .CO(n29631));
    SB_CARRY rem_4_add_916_9 (.CI(n28547), .I0(n1351), .I1(VCC_net), .CO(n28548));
    SB_LUT4 div_46_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4529), .I3(n29369), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n29629), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_9 (.CI(n29629), .I0(n1752), .I1(VCC_net), 
            .CO(n29630));
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n30482), .I0(GND_net), .I1(n21_adj_4939), 
            .CO(n30483));
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n29628), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n29628), .I0(n1753), .I1(VCC_net), 
            .CO(n29629));
    SB_LUT4 rem_4_i926_rep_74_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), 
            .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i926_rep_74_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2295_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n29087), 
            .O(n6140)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1754_adj_4454), .I2(GND_net), 
            .I3(n29627), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4940), .I3(n30481), .O(n22_adj_4421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4545));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4921));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13292_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[6] [3]), 
            .I2(n17068), .I3(GND_net), .O(n18037));   // verilog/coms.v(126[12] 289[6])
    defparam i13292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4544));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13154_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n35418), 
            .I3(GND_net), .O(n17899));   // verilog/coms.v(126[12] 289[6])
    defparam i13154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4838));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4836));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4840));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4839));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4339), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n531));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4833));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4834));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4822));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4831));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4832));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4826));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4828));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4829));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4835));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4824));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4830));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35104_4_lut (.I0(n29_adj_4835), .I1(n17_adj_4829), .I2(n15_adj_4828), 
            .I3(n13_adj_4826), .O(n41958));
    defparam i35104_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35773_4_lut (.I0(n11_adj_4824), .I1(n9_adj_4822), .I2(n2719), 
            .I3(n98), .O(n42627));
    defparam i35773_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i36036_4_lut (.I0(n17_adj_4829), .I1(n15_adj_4828), .I2(n13_adj_4826), 
            .I3(n42627), .O(n42890));
    defparam i36036_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36030_4_lut (.I0(n23_adj_4832), .I1(n21_adj_4831), .I2(n19_adj_4830), 
            .I3(n42890), .O(n42884));
    defparam i36030_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_577_5 (.CI(n28664), .I0(n44224), .I1(n22), .CO(n28665));
    SB_LUT4 i35106_4_lut (.I0(n29_adj_4835), .I1(n27_adj_4834), .I2(n25_adj_4833), 
            .I3(n42884), .O(n41960));
    defparam i35106_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1777_i6_4_lut (.I0(n531), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4820));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i13363_4_lut (.I0(n38107), .I1(byte_transmit_counter[0]), .I2(n7821), 
            .I3(n17100), .O(n18108));   // verilog/coms.v(126[12] 289[6])
    defparam i13363_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY add_2295_12 (.CI(n29087), .I0(n2629), .I1(n90), .CO(n29088));
    SB_LUT4 i13360_3_lut (.I0(n17330), .I1(r_Bit_Index_adj_5028[0]), .I2(n17186), 
            .I3(GND_net), .O(n18105));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13360_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 add_2295_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n29086), 
            .O(n6141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36066_3_lut (.I0(n6_adj_4820), .I1(n87), .I2(n29_adj_4835), 
            .I3(GND_net), .O(n42920));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36066_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_46_unary_minus_4_add_3_15 (.CI(n29369), .I0(GND_net), .I1(n12_adj_4529), 
            .CO(n29370));
    SB_CARRY add_2295_11 (.CI(n29086), .I0(n2630), .I1(n91), .CO(n29087));
    SB_CARRY rem_4_add_1184_7 (.CI(n29627), .I0(n1754_adj_4454), .I1(GND_net), 
            .CO(n29628));
    SB_LUT4 add_2295_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n29085), 
            .O(n6142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_10 (.CI(n29085), .I0(n2631), .I1(n92), .CO(n29086));
    SB_LUT4 add_2295_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n29084), 
            .O(n6143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4530), .I3(n29368), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_9 (.CI(n29084), .I0(n2632), .I1(n93), .CO(n29085));
    SB_CARRY div_46_unary_minus_4_add_3_14 (.CI(n29368), .I0(GND_net), .I1(n13_adj_4530), 
            .CO(n29369));
    SB_LUT4 div_46_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4531), .I3(n29367), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1777_i32_3_lut (.I0(n14_adj_4827), .I1(n83), 
            .I2(n37_adj_4840), .I3(GND_net), .O(n32_adj_4837));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36067_3_lut (.I0(n42920), .I1(n86), .I2(n31_adj_4836), .I3(GND_net), 
            .O(n42921));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36067_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35089_4_lut (.I0(n35_adj_4839), .I1(n33_adj_4838), .I2(n31_adj_4836), 
            .I3(n41958), .O(n41943));
    defparam i35089_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36470_4_lut (.I0(n32_adj_4837), .I1(n12_adj_4825), .I2(n37_adj_4840), 
            .I3(n41934), .O(n43324));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36470_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35456_3_lut (.I0(n42921), .I1(n85), .I2(n33_adj_4838), .I3(GND_net), 
            .O(n42310));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35456_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36068_3_lut (.I0(n8_adj_4821), .I1(n90), .I2(n23_adj_4832), 
            .I3(GND_net), .O(n42922));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36068_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36069_3_lut (.I0(n42922), .I1(n89), .I2(n25_adj_4833), .I3(GND_net), 
            .O(n42923));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36069_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35751_4_lut (.I0(n25_adj_4833), .I1(n23_adj_4832), .I2(n21_adj_4831), 
            .I3(n41984), .O(n42605));
    defparam i35751_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37343_4_lut (.I0(r_SM_Main[2]), .I1(n41247), .I2(n41248), 
            .I3(r_SM_Main[1]), .O(n25741));
    defparam i37343_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i35888_3_lut (.I0(n10_adj_4823), .I1(n91), .I2(n21_adj_4831), 
            .I3(GND_net), .O(n42742));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35888_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35454_3_lut (.I0(n42923), .I1(n88), .I2(n27_adj_4834), .I3(GND_net), 
            .O(n42308));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35454_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36251_4_lut (.I0(n35_adj_4839), .I1(n33_adj_4838), .I2(n31_adj_4836), 
            .I3(n41960), .O(n43105));
    defparam i36251_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36580_4_lut (.I0(n42310), .I1(n43324), .I2(n37_adj_4840), 
            .I3(n41943), .O(n43434));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36580_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36062_4_lut (.I0(n42308), .I1(n42742), .I2(n27_adj_4834), 
            .I3(n42605), .O(n42916));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36062_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36624_4_lut (.I0(n42916), .I1(n43434), .I2(n37_adj_4840), 
            .I3(n43105), .O(n43478));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36624_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36625_3_lut (.I0(n43478), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n43479));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36625_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36621_3_lut (.I0(n43479), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n43475));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36621_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36296_3_lut (.I0(n43475), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n43150));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36296_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36297_3_lut (.I0(n43150), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n43151));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36297_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i2018_4_lut (.I0(n43151), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i2018_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i13009_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13293), .I3(GND_net), .O(n17754));   // verilog/coms.v(126[12] 289[6])
    defparam i13009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4815));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4817));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4813));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4338), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n530));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4816));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1755_adj_4455), .I2(GND_net), 
            .I3(n29626), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_6 (.CI(n29626), .I0(n1755_adj_4455), .I1(GND_net), 
            .CO(n29627));
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n30481), .I0(GND_net), .I1(n22_adj_4940), 
            .CO(n30482));
    SB_LUT4 div_46_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4809));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n28546), .O(n1419_adj_4495)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2295_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n29083), 
            .O(n6144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4941), .I3(n30480), .O(n23_adj_4420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4810));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4797));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4807));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4808));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4799));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13356_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n37457), 
            .I3(GND_net), .O(n18101));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13356_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1756_adj_4456), .I2(VCC_net), 
            .I3(n29625), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_13 (.CI(n29367), .I0(GND_net), .I1(n14_adj_4531), 
            .CO(n29368));
    SB_LUT4 div_46_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4801));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n30480), .I0(GND_net), .I1(n23_adj_4941), 
            .CO(n30481));
    SB_LUT4 rem_4_i1660_3_lut (.I0(n2443), .I1(n2510), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2542_adj_4509));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_5 (.CI(n29625), .I0(n1756_adj_4456), .I1(VCC_net), 
            .CO(n29626));
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4942), .I3(n30479), .O(n24_adj_4419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1757_adj_4457), .I2(VCC_net), 
            .I3(n29624), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_4 (.CI(n29624), .I0(n1757_adj_4457), .I1(VCC_net), 
            .CO(n29625));
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n30479), .I0(GND_net), .I1(n24_adj_4942), 
            .CO(n30480));
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4943), .I3(n30478), .O(n25_adj_4418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_8 (.CI(n29083), .I0(n2633), .I1(n94), .CO(n29084));
    SB_LUT4 div_46_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4803));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4804));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4811));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4806));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34490_4_lut (.I0(n31_adj_4811), .I1(n19_adj_4804), .I2(n17_adj_4803), 
            .I3(n15_adj_4801), .O(n41343));
    defparam i34490_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35233_4_lut (.I0(n13_adj_4799), .I1(n11_adj_4797), .I2(n2637), 
            .I3(n98), .O(n42087));
    defparam i35233_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i35811_4_lut (.I0(n19_adj_4804), .I1(n17_adj_4803), .I2(n15_adj_4801), 
            .I3(n42087), .O(n42665));
    defparam i35811_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35809_4_lut (.I0(n25_adj_4808), .I1(n23_adj_4807), .I2(n21_adj_4806), 
            .I3(n42665), .O(n42663));
    defparam i35809_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1758_adj_4458), .I2(GND_net), 
            .I3(n29623), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4532), .I3(n29366), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n30478), .I0(GND_net), .I1(n25_adj_4943), 
            .CO(n30479));
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_4944), .I3(n30477), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542_adj_4509), .I1(n2609), .I2(n2570), 
            .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_3 (.CI(n29623), .I0(n1758_adj_4458), .I1(GND_net), 
            .CO(n29624));
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1858), .I1(VCC_net), 
            .CO(n29623));
    SB_LUT4 i34494_4_lut (.I0(n31_adj_4811), .I1(n29_adj_4810), .I2(n27_adj_4809), 
            .I3(n42663), .O(n41347));
    defparam i34494_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n30477), .I0(GND_net), .I1(n26_adj_4944), 
            .CO(n30478));
    SB_CARRY div_46_unary_minus_4_add_3_12 (.CI(n29366), .I0(GND_net), .I1(n15_adj_4532), 
            .CO(n29367));
    SB_LUT4 div_46_LessThan_1722_i8_4_lut (.I0(n530), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4795));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36276_3_lut (.I0(n8_adj_4795), .I1(n87), .I2(n31_adj_4811), 
            .I3(GND_net), .O(n43130));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36276_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2295_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n29082), 
            .O(n6145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_7 (.CI(n29082), .I0(n2634), .I1(n95), .CO(n29083));
    SB_LUT4 add_2295_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n29081), 
            .O(n6146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_6 (.CI(n29081), .I0(n2635), .I1(n96), .CO(n29082));
    SB_LUT4 add_2295_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n29080), 
            .O(n6147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_5 (.CI(n29080), .I0(n2636), .I1(n97), .CO(n29081));
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_4945), .I3(n30476), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2295_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n29079), 
            .O(n6148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_17_lut (.I0(n1877), .I1(n1844), .I2(VCC_net), 
            .I3(n29622), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4533), .I3(n29365), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_16_lut (.I0(GND_net), .I1(n1845), .I2(VCC_net), 
            .I3(n29621), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36277_3_lut (.I0(n43130), .I1(n86), .I2(n33_adj_4813), .I3(GND_net), 
            .O(n43131));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36277_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2295_4 (.CI(n29079), .I0(n2637), .I1(n98), .CO(n29080));
    SB_LUT4 add_2295_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n29078), 
            .O(n6149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_11 (.CI(n29365), .I0(GND_net), .I1(n16_adj_4533), 
            .CO(n29366));
    SB_CARRY rem_4_add_1251_16 (.CI(n29621), .I0(n1845), .I1(VCC_net), 
            .CO(n29622));
    SB_CARRY add_2295_3 (.CI(n29078), .I0(n2638), .I1(n99), .CO(n29079));
    SB_LUT4 add_2295_2_lut (.I0(GND_net), .I1(n530), .I2(n558), .I3(VCC_net), 
            .O(n6150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2295_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2295_2 (.CI(VCC_net), .I0(n530), .I1(n558), .CO(n29078));
    SB_LUT4 add_2294_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n29077), 
            .O(n6106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4534), .I3(n29364), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2294_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n29076), 
            .O(n6107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i34_3_lut (.I0(n16_adj_4802), .I1(n83), 
            .I2(n39_adj_4817), .I3(GND_net), .O(n34_adj_4814));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n30476), .I0(GND_net), .I1(n27_adj_4945), 
            .CO(n30477));
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_4946), .I3(n30475), .O(n28_adj_4417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n30475), .I0(GND_net), .I1(n28_adj_4946), 
            .CO(n30476));
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_4947), .I3(n30474), .O(n29_adj_4416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n30474), .I0(GND_net), .I1(n29_adj_4947), 
            .CO(n30475));
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_4948), .I3(n30473), .O(n30_adj_4415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34474_4_lut (.I0(n37_adj_4816), .I1(n35_adj_4815), .I2(n33_adj_4813), 
            .I3(n41343), .O(n41327));
    defparam i34474_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36468_4_lut (.I0(n34_adj_4814), .I1(n14_adj_4800), .I2(n39_adj_4817), 
            .I3(n41323), .O(n43322));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36468_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36170_3_lut (.I0(n43131), .I1(n85), .I2(n35_adj_4815), .I3(GND_net), 
            .O(n32_adj_4812));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36170_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36278_3_lut (.I0(n10_adj_4796), .I1(n90), .I2(n25_adj_4808), 
            .I3(GND_net), .O(n43132));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36278_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1251_15_lut (.I0(GND_net), .I1(n1846), .I2(VCC_net), 
            .I3(n29620), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_10 (.CI(n29364), .I0(GND_net), .I1(n17_adj_4534), 
            .CO(n29365));
    SB_CARRY add_2294_21 (.CI(n29076), .I0(n2535), .I1(n81), .CO(n29077));
    SB_CARRY rem_4_add_1251_15 (.CI(n29620), .I0(n1846), .I1(VCC_net), 
            .CO(n29621));
    SB_LUT4 div_46_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4535), .I3(n29363), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_14_lut (.I0(GND_net), .I1(n1847), .I2(VCC_net), 
            .I3(n29619), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_9 (.CI(n29363), .I0(GND_net), .I1(n18_adj_4535), 
            .CO(n29364));
    SB_LUT4 add_2294_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n29075), 
            .O(n6108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_577_4_lut (.I0(duty[2]), .I1(n44224), .I2(n23), .I3(n28663), 
            .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2294_20 (.CI(n29075), .I0(n2536), .I1(n82), .CO(n29076));
    SB_CARRY rem_4_add_1251_14 (.CI(n29619), .I0(n1847), .I1(VCC_net), 
            .CO(n29620));
    SB_LUT4 div_46_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4536), .I3(n29362), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2294_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n29074), 
            .O(n6109)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_19 (.CI(n29074), .I0(n2537), .I1(n83), .CO(n29075));
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n30473), .I0(GND_net), .I1(n30_adj_4948), 
            .CO(n30474));
    SB_LUT4 rem_4_add_1251_13_lut (.I0(GND_net), .I1(n1848), .I2(VCC_net), 
            .I3(n29618), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_8 (.CI(n29362), .I0(GND_net), .I1(n19_adj_4536), 
            .CO(n29363));
    SB_CARRY rem_4_add_1251_13 (.CI(n29618), .I0(n1848), .I1(VCC_net), 
            .CO(n29619));
    SB_LUT4 rem_4_add_1251_12_lut (.I0(GND_net), .I1(n1849), .I2(VCC_net), 
            .I3(n29617), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4537), .I3(n29361), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2294_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n29073), 
            .O(n6110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_18 (.CI(n29073), .I0(n2538), .I1(n84), .CO(n29074));
    SB_CARRY rem_4_add_1251_12 (.CI(n29617), .I0(n1849), .I1(VCC_net), 
            .CO(n29618));
    SB_CARRY div_46_unary_minus_4_add_3_7 (.CI(n29361), .I0(GND_net), .I1(n20_adj_4537), 
            .CO(n29362));
    SB_LUT4 add_2294_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n29072), 
            .O(n6111)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_11_lut (.I0(GND_net), .I1(n1850), .I2(VCC_net), 
            .I3(n29616), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4538), .I3(n29360), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_4949), .I3(n30472), .O(n31_adj_4414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_11 (.CI(n29616), .I0(n1850), .I1(VCC_net), 
            .CO(n29617));
    SB_CARRY div_46_unary_minus_4_add_3_6 (.CI(n29360), .I0(GND_net), .I1(n21_adj_4538), 
            .CO(n29361));
    SB_CARRY add_2294_17 (.CI(n29072), .I0(n2539), .I1(n85), .CO(n29073));
    SB_LUT4 rem_4_add_1251_10_lut (.I0(GND_net), .I1(n1851), .I2(VCC_net), 
            .I3(n29615), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4539), .I3(n29359), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2294_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n29071), 
            .O(n6112)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_4 (.CI(n28663), .I0(n44224), .I1(n23), .CO(n28664));
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n30472), .I0(GND_net), .I1(n31_adj_4949), 
            .CO(n30473));
    SB_CARRY rem_4_add_1251_10 (.CI(n29615), .I0(n1851), .I1(VCC_net), 
            .CO(n29616));
    SB_CARRY div_46_unary_minus_4_add_3_5 (.CI(n29359), .I0(GND_net), .I1(n22_adj_4539), 
            .CO(n29360));
    SB_LUT4 rem_4_add_1251_9_lut (.I0(GND_net), .I1(n1852), .I2(VCC_net), 
            .I3(n29614), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4540), .I3(n29358), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_9 (.CI(n29614), .I0(n1852), .I1(VCC_net), 
            .CO(n29615));
    SB_CARRY div_46_unary_minus_4_add_3_4 (.CI(n29358), .I0(GND_net), .I1(n23_adj_4540), 
            .CO(n29359));
    SB_CARRY add_2294_16 (.CI(n29071), .I0(n2540), .I1(n86), .CO(n29072));
    SB_LUT4 rem_4_add_1251_8_lut (.I0(GND_net), .I1(n1853), .I2(VCC_net), 
            .I3(n29613), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4541), .I3(n29357), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2294_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n29070), 
            .O(n6113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_4950), .I3(n30471), .O(n32_adj_4413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_8 (.CI(n29613), .I0(n1853), .I1(VCC_net), 
            .CO(n29614));
    SB_CARRY div_46_unary_minus_4_add_3_3 (.CI(n29357), .I0(GND_net), .I1(n24_adj_4541), 
            .CO(n29358));
    SB_CARRY add_2294_15 (.CI(n29070), .I0(n2541), .I1(n87), .CO(n29071));
    SB_LUT4 add_577_3_lut (.I0(duty[1]), .I1(n44224), .I2(n24), .I3(n28662), 
            .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2294_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n29069), 
            .O(n6114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_14 (.CI(n29069), .I0(n2542), .I1(n88), .CO(n29070));
    SB_LUT4 rem_4_add_1251_7_lut (.I0(GND_net), .I1(n1854), .I2(GND_net), 
            .I3(n29612), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4542), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_8 (.CI(n28546), .I0(n1352), .I1(VCC_net), .CO(n28547));
    SB_LUT4 add_2294_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n29068), 
            .O(n6115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_13 (.CI(n29068), .I0(n2543), .I1(n89), .CO(n29069));
    SB_LUT4 add_2294_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n29067), 
            .O(n6116)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_7 (.CI(n29612), .I0(n1854), .I1(GND_net), 
            .CO(n29613));
    SB_CARRY div_46_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4542), 
            .CO(n29357));
    SB_CARRY add_2294_12 (.CI(n29067), .I0(n2544), .I1(n90), .CO(n29068));
    SB_LUT4 add_2294_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n29066), 
            .O(n6117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_11 (.CI(n29066), .I0(n2545), .I1(n91), .CO(n29067));
    SB_LUT4 rem_4_add_1251_6_lut (.I0(GND_net), .I1(n1855), .I2(GND_net), 
            .I3(n29611), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_28_lut (.I0(n2933), .I1(n2933), .I2(n2966_adj_4400), 
            .I3(n29356), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n28545), .O(n1420_adj_4496)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_577_3 (.CI(n28662), .I0(n44224), .I1(n24), .CO(n28663));
    SB_LUT4 add_577_2_lut (.I0(duty[0]), .I1(n44224), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_577_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2294_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n29065), 
            .O(n6118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_10 (.CI(n29065), .I0(n2546), .I1(n92), .CO(n29066));
    SB_LUT4 add_2294_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n29064), 
            .O(n6119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_9 (.CI(n29064), .I0(n2547), .I1(n93), .CO(n29065));
    SB_LUT4 add_2294_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n29063), 
            .O(n6120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_8 (.CI(n29063), .I0(n2548), .I1(n94), .CO(n29064));
    SB_CARRY rem_4_add_1251_6 (.CI(n29611), .I0(n1855), .I1(GND_net), 
            .CO(n29612));
    SB_LUT4 rem_4_add_1988_27_lut (.I0(n2934), .I1(n2934), .I2(n2966_adj_4400), 
            .I3(n29355), .O(n3033)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_577_2 (.CI(VCC_net), .I0(n44224), .I1(n25), .CO(n28662));
    SB_LUT4 rem_4_add_1251_5_lut (.I0(GND_net), .I1(n1856), .I2(VCC_net), 
            .I3(n29610), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_27 (.CI(n29355), .I0(n2934), .I1(n2966_adj_4400), 
            .CO(n29356));
    SB_CARRY rem_4_add_916_7 (.CI(n28545), .I0(n1353), .I1(VCC_net), .CO(n28546));
    SB_LUT4 add_2294_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n29062), 
            .O(n6121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_7 (.CI(n29062), .I0(n2549), .I1(n95), .CO(n29063));
    SB_CARRY rem_4_add_1251_5 (.CI(n29610), .I0(n1856), .I1(VCC_net), 
            .CO(n29611));
    SB_LUT4 rem_4_add_1988_26_lut (.I0(n2935), .I1(n2935), .I2(n2966_adj_4400), 
            .I3(n29354), .O(n3034)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n30471), .I0(GND_net), .I1(n32_adj_4950), 
            .CO(n30472));
    SB_LUT4 rem_4_add_1251_4_lut (.I0(GND_net), .I1(n1857), .I2(VCC_net), 
            .I3(n29609), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_26 (.CI(n29354), .I0(n2935), .I1(n2966_adj_4400), 
            .CO(n29355));
    SB_LUT4 rem_4_add_1988_25_lut (.I0(n2936), .I1(n2936), .I2(n2966_adj_4400), 
            .I3(n29353), .O(n3035)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_4951), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_4 (.CI(n29609), .I0(n1857), .I1(VCC_net), 
            .CO(n29610));
    SB_CARRY rem_4_add_1988_25 (.CI(n29353), .I0(n2936), .I1(n2966_adj_4400), 
            .CO(n29354));
    SB_LUT4 i36279_3_lut (.I0(n43132), .I1(n89), .I2(n27_adj_4809), .I3(GND_net), 
            .O(n43133));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36279_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n28544), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1684 (.I0(n36403), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));
    defparam i3_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1251_3_lut (.I0(GND_net), .I1(n1858), .I2(GND_net), 
            .I3(n29608), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_24_lut (.I0(n2937), .I1(n2937), .I2(n2966_adj_4400), 
            .I3(n29352), .O(n3036)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_916_6 (.CI(n28544), .I0(n1354), .I1(GND_net), .CO(n28545));
    SB_CARRY rem_4_add_1251_3 (.CI(n29608), .I0(n1858), .I1(GND_net), 
            .CO(n29609));
    SB_CARRY rem_4_add_1988_24 (.CI(n29352), .I0(n2937), .I1(n2966_adj_4400), 
            .CO(n29353));
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1958), .I1(VCC_net), 
            .CO(n29608));
    SB_LUT4 rem_4_add_1318_18_lut (.I0(n1976_adj_4628), .I1(n1943), .I2(VCC_net), 
            .I3(n29607), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_23_lut (.I0(n2938), .I1(n2938), .I2(n2966_adj_4400), 
            .I3(n29351), .O(n3037)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1988_23 (.CI(n29351), .I0(n2938), .I1(n2966_adj_4400), 
            .CO(n29352));
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_4951), 
            .CO(n30471));
    SB_LUT4 rem_4_add_1318_17_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n29606), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_22_lut (.I0(n2939), .I1(n2939), .I2(n2966_adj_4400), 
            .I3(n29350), .O(n3038)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2294_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n29061), 
            .O(n6122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_6 (.CI(n29061), .I0(n2550), .I1(n96), .CO(n29062));
    SB_LUT4 add_2294_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n29060), 
            .O(n6123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_5 (.CI(n29060), .I0(n2551), .I1(n97), .CO(n29061));
    SB_LUT4 add_2294_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n29059), 
            .O(n6124)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_4 (.CI(n29059), .I0(n2552), .I1(n98), .CO(n29060));
    SB_LUT4 add_2294_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n29058), 
            .O(n6125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_3 (.CI(n29058), .I0(n2553), .I1(n99), .CO(n29059));
    SB_LUT4 add_2294_2_lut (.I0(GND_net), .I1(n529), .I2(n558), .I3(VCC_net), 
            .O(n6126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2294_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2294_2 (.CI(VCC_net), .I0(n529), .I1(n558), .CO(n29058));
    SB_LUT4 add_2293_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n29057), 
            .O(n6084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2293_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n29056), 
            .O(n6085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_20 (.CI(n29056), .I0(n2448), .I1(n82), .CO(n29057));
    SB_LUT4 add_2293_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n29055), 
            .O(n6086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_19 (.CI(n29055), .I0(n2449), .I1(n83), .CO(n29056));
    SB_LUT4 add_2293_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n29054), 
            .O(n6087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_18 (.CI(n29054), .I0(n2450), .I1(n84), .CO(n29055));
    SB_LUT4 add_2293_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n29053), 
            .O(n6088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_17 (.CI(n29053), .I0(n2451), .I1(n85), .CO(n29054));
    SB_LUT4 add_2293_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n29052), 
            .O(n6089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_16 (.CI(n29052), .I0(n2452), .I1(n86), .CO(n29053));
    SB_LUT4 add_2293_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n29051), 
            .O(n6090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_15 (.CI(n29051), .I0(n2453), .I1(n87), .CO(n29052));
    SB_LUT4 add_2293_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n29050), 
            .O(n6091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_14 (.CI(n29050), .I0(n2454), .I1(n88), .CO(n29051));
    SB_LUT4 add_2293_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n29049), 
            .O(n6092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_13 (.CI(n29049), .I0(n2455), .I1(n89), .CO(n29050));
    SB_LUT4 add_2293_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n29048), 
            .O(n6093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_12 (.CI(n29048), .I0(n2456), .I1(n90), .CO(n29049));
    SB_LUT4 add_2293_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n29047), 
            .O(n6094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_17 (.CI(n29606), .I0(n1944), .I1(VCC_net), 
            .CO(n29607));
    SB_CARRY rem_4_add_1988_22 (.CI(n29350), .I0(n2939), .I1(n2966_adj_4400), 
            .CO(n29351));
    SB_LUT4 rem_4_add_1988_21_lut (.I0(n2940), .I1(n2940), .I2(n2966_adj_4400), 
            .I3(n29349), .O(n3039)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n29605), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n29605), .I0(n1945), .I1(VCC_net), 
            .CO(n29606));
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n29604), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_21 (.CI(n29349), .I0(n2940), .I1(n2966_adj_4400), 
            .CO(n29350));
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n28543), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1685 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n36401));
    defparam i1_3_lut_adj_1685.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n1254), .I1(n1250), .I2(n36401), .I3(n1255), 
            .O(n6_adj_4900));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1687 (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4900), 
            .O(n1283));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i4_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1688 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n36397));
    defparam i1_3_lut_adj_1688.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1689 (.I0(n1351), .I1(n1354), .I2(n36397), .I3(n1355), 
            .O(n8_adj_4397));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i2_4_lut_adj_1689.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1690 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4398));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i1_2_lut_adj_1690.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1691 (.I0(n1352), .I1(n7_adj_4398), .I2(n1353), 
            .I3(n8_adj_4397), .O(n1382));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1692 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n38647));
    defparam i1_2_lut_adj_1692.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1693 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16_adj_4393));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i6_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1694 (.I0(n1756_adj_4456), .I1(n1757_adj_4457), 
            .I2(n1758_adj_4458), .I3(GND_net), .O(n36450));
    defparam i1_3_lut_adj_1694.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1751), .I1(n16_adj_4393), .I2(n1753), .I3(GND_net), 
            .O(n18_adj_4392));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_2293_11 (.CI(n29047), .I0(n2457), .I1(n91), .CO(n29048));
    SB_LUT4 i35219_4_lut (.I0(n27_adj_4809), .I1(n25_adj_4808), .I2(n23_adj_4807), 
            .I3(n41363), .O(n42073));
    defparam i35219_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1722_i20_3_lut (.I0(n12_adj_4798), .I1(n91), 
            .I2(n23_adj_4807), .I3(GND_net), .O(n20_adj_4805));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36168_3_lut (.I0(n43133), .I1(n88), .I2(n29_adj_4810), .I3(GND_net), 
            .O(n43022));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36168_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2293_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n29046), 
            .O(n6095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_10 (.CI(n29046), .I0(n2458), .I1(n92), .CO(n29047));
    SB_CARRY rem_4_add_1318_15 (.CI(n29604), .I0(n1946), .I1(VCC_net), 
            .CO(n29605));
    SB_LUT4 rem_4_add_1988_20_lut (.I0(n2941), .I1(n2941), .I2(n2966_adj_4400), 
            .I3(n29348), .O(n3040)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36044_4_lut (.I0(n37_adj_4816), .I1(n35_adj_4815), .I2(n33_adj_4813), 
            .I3(n41347), .O(n42898));
    defparam i36044_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n29603), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36516_4_lut (.I0(n32_adj_4812), .I1(n43322), .I2(n39_adj_4817), 
            .I3(n41327), .O(n43370));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36516_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36171_4_lut (.I0(n43022), .I1(n20_adj_4805), .I2(n29_adj_4810), 
            .I3(n42073), .O(n43025));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36171_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36608_4_lut (.I0(n43025), .I1(n43370), .I2(n39_adj_4817), 
            .I3(n42898), .O(n43462));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36608_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36609_3_lut (.I0(n43462), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n43463));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36609_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY rem_4_add_916_5 (.CI(n28543), .I0(n1355), .I1(GND_net), .CO(n28544));
    SB_LUT4 add_2293_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n29045), 
            .O(n6096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36275_3_lut (.I0(n43463), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n43129));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36275_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY add_2293_9 (.CI(n29045), .I0(n2459), .I1(n93), .CO(n29046));
    SB_CARRY rem_4_add_1318_14 (.CI(n29603), .I0(n1947), .I1(VCC_net), 
            .CO(n29604));
    SB_CARRY rem_4_add_1988_20 (.CI(n29348), .I0(n2941), .I1(n2966_adj_4400), 
            .CO(n29349));
    SB_LUT4 i36173_3_lut (.I0(n43129), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n43027));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36173_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n43027), .I1(n15962), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4543));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2293_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n29044), 
            .O(n6097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_8 (.CI(n29044), .I0(n2460), .I1(n94), .CO(n29045));
    SB_LUT4 add_2293_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n29043), 
            .O(n6098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_19_lut (.I0(n2942), .I1(n2942), .I2(n2966_adj_4400), 
            .I3(n29347), .O(n3041)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n28542), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_7 (.CI(n29043), .I0(n2461), .I1(n95), .CO(n29044));
    SB_LUT4 add_2293_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n29042), 
            .O(n6099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_6 (.CI(n29042), .I0(n2462), .I1(n96), .CO(n29043));
    SB_LUT4 add_2293_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n29041), 
            .O(n6100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_5 (.CI(n29041), .I0(n2463), .I1(n97), .CO(n29042));
    SB_LUT4 add_2293_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n29040), 
            .O(n6101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_4 (.CI(n29040), .I0(n2464), .I1(n98), .CO(n29041));
    SB_LUT4 add_2293_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n29039), 
            .O(n6102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_3 (.CI(n29039), .I0(n2465), .I1(n99), .CO(n29040));
    SB_LUT4 add_2293_2_lut (.I0(GND_net), .I1(n528), .I2(n558), .I3(VCC_net), 
            .O(n6103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2293_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2293_2 (.CI(VCC_net), .I0(n528), .I1(n558), .CO(n29039));
    SB_LUT4 add_2292_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n29038), 
            .O(n6063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2292_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n29037), 
            .O(n6064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_19 (.CI(n29037), .I0(n2358), .I1(n83), .CO(n29038));
    SB_LUT4 add_2292_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n29036), 
            .O(n6065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_18 (.CI(n29036), .I0(n2359), .I1(n84), .CO(n29037));
    SB_LUT4 add_2292_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n29035), 
            .O(n6066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_17 (.CI(n29035), .I0(n2360), .I1(n85), .CO(n29036));
    SB_LUT4 add_2292_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n29034), 
            .O(n6067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_16 (.CI(n29034), .I0(n2361), .I1(n86), .CO(n29035));
    SB_LUT4 add_2292_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n29033), 
            .O(n6068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_15 (.CI(n29033), .I0(n2362), .I1(n87), .CO(n29034));
    SB_LUT4 add_2292_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n29032), 
            .O(n6069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1696 (.I0(n1754_adj_4454), .I1(n1749), .I2(n36450), 
            .I3(n1755_adj_4455), .O(n13_adj_4394));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i3_4_lut_adj_1696.LUT_INIT = 16'heccc;
    SB_CARRY add_2292_14 (.CI(n29032), .I0(n2363), .I1(n88), .CO(n29033));
    SB_CARRY rem_4_add_916_4 (.CI(n28542), .I0(n1356), .I1(VCC_net), .CO(n28543));
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n29602), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2292_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n29031), 
            .O(n6070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_13 (.CI(n29031), .I0(n2364), .I1(n89), .CO(n29032));
    SB_LUT4 add_2292_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n29030), 
            .O(n6071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_12 (.CI(n29030), .I0(n2365), .I1(n90), .CO(n29031));
    SB_LUT4 add_2292_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n29029), 
            .O(n6072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_11 (.CI(n29029), .I0(n2366), .I1(n91), .CO(n29030));
    SB_LUT4 add_2292_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n29028), 
            .O(n6073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_10 (.CI(n29028), .I0(n2367), .I1(n92), .CO(n29029));
    SB_LUT4 add_2292_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n29027), 
            .O(n6074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1199__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_CARRY add_2292_9 (.CI(n29027), .I0(n2368), .I1(n93), .CO(n29028));
    SB_LUT4 add_2292_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n29026), 
            .O(n6075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_8 (.CI(n29026), .I0(n2369), .I1(n94), .CO(n29027));
    SB_LUT4 add_2292_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n29025), 
            .O(n6076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_7 (.CI(n29025), .I0(n2370), .I1(n95), .CO(n29026));
    SB_LUT4 add_2292_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n29024), 
            .O(n6077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_6 (.CI(n29024), .I0(n2371), .I1(n96), .CO(n29025));
    SB_CARRY rem_4_add_1318_13 (.CI(n29602), .I0(n1948), .I1(VCC_net), 
            .CO(n29603));
    SB_CARRY rem_4_add_1988_19 (.CI(n29347), .I0(n2942), .I1(n2966_adj_4400), 
            .CO(n29348));
    SB_LUT4 add_2292_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n29023), 
            .O(n6078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_5 (.CI(n29023), .I0(n2372), .I1(n97), .CO(n29024));
    SB_LUT4 rem_4_add_1988_18_lut (.I0(n2943), .I1(n2943), .I2(n2966_adj_4400), 
            .I3(n29346), .O(n3042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2292_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n29022), 
            .O(n6079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4792));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4794));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2292_4 (.CI(n29022), .I0(n2373), .I1(n98), .CO(n29023));
    SB_CARRY rem_4_add_1988_18 (.CI(n29346), .I0(n2943), .I1(n2966_adj_4400), 
            .CO(n29347));
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n29601), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n28541), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_12 (.CI(n29601), .I0(n1949), .I1(VCC_net), 
            .CO(n29602));
    SB_LUT4 div_46_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4790));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4337), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n529));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2292_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n29021), 
            .O(n6080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2292_3 (.CI(n29021), .I0(n2374), .I1(n99), .CO(n29022));
    SB_LUT4 rem_4_add_1988_17_lut (.I0(n2944), .I1(n2944), .I2(n2966_adj_4400), 
            .I3(n29345), .O(n3043)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n29600), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1697 (.I0(n13_adj_4394), .I1(n18_adj_4392), .I2(n1752), 
            .I3(n1750), .O(n1778_adj_4818));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i9_4_lut_adj_1697.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4793));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4787));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4788));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4775));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2292_2_lut (.I0(GND_net), .I1(n527), .I2(n558), .I3(VCC_net), 
            .O(n6081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2292_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_11 (.CI(n29600), .I0(n1950), .I1(VCC_net), 
            .CO(n29601));
    SB_CARRY add_2292_2 (.CI(VCC_net), .I0(n527), .I1(n558), .CO(n29021));
    SB_LUT4 div_46_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4777));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n29599), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_10 (.CI(n29599), .I0(n1951), .I1(VCC_net), 
            .CO(n29600));
    SB_LUT4 add_5547_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n29020), 
            .O(n10218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5547_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n29019), 
            .O(n10219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5547_6 (.CI(n29019), .I0(n3354), .I1(GND_net), .CO(n29020));
    SB_LUT4 add_5547_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n29018), 
            .O(n10220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5547_5 (.CI(n29018), .I0(n3355), .I1(GND_net), .CO(n29019));
    SB_LUT4 add_5547_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n29017), 
            .O(n10221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5547_4 (.CI(n29017), .I0(n3356), .I1(VCC_net), .CO(n29018));
    SB_LUT4 add_5547_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n29016), 
            .O(n10222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5547_3 (.CI(n29016), .I0(n3357), .I1(VCC_net), .CO(n29017));
    SB_LUT4 add_5547_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5547_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5547_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n29016));
    SB_LUT4 add_2291_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n29015), 
            .O(n6043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2291_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n29014), 
            .O(n6044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_18 (.CI(n29014), .I0(n2265), .I1(n84), .CO(n29015));
    SB_LUT4 add_2291_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n29013), 
            .O(n6045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_17 (.CI(n29013), .I0(n2266), .I1(n85), .CO(n29014));
    SB_LUT4 add_2291_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n29012), 
            .O(n6046)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_16 (.CI(n29012), .I0(n2267), .I1(n86), .CO(n29013));
    SB_LUT4 add_2291_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n29011), 
            .O(n6047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_15 (.CI(n29011), .I0(n2268), .I1(n87), .CO(n29012));
    SB_LUT4 add_2291_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n29010), 
            .O(n6048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_14 (.CI(n29010), .I0(n2269), .I1(n88), .CO(n29011));
    SB_LUT4 add_2291_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n29009), 
            .O(n6049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_13 (.CI(n29009), .I0(n2270), .I1(n89), .CO(n29010));
    SB_LUT4 add_2291_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n29008), 
            .O(n6050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_12 (.CI(n29008), .I0(n2271), .I1(n90), .CO(n29009));
    SB_LUT4 add_2291_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n29007), 
            .O(n6051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_11 (.CI(n29007), .I0(n2272), .I1(n91), .CO(n29008));
    SB_LUT4 add_2291_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n29006), 
            .O(n6052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_10 (.CI(n29006), .I0(n2273), .I1(n92), .CO(n29007));
    SB_LUT4 add_2291_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n29005), 
            .O(n6053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_9 (.CI(n29005), .I0(n2274), .I1(n93), .CO(n29006));
    SB_LUT4 add_2291_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n29004), 
            .O(n6054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_8 (.CI(n29004), .I0(n2275), .I1(n94), .CO(n29005));
    SB_LUT4 add_2291_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n29003), 
            .O(n6055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_7 (.CI(n29003), .I0(n2276), .I1(n95), .CO(n29004));
    SB_LUT4 add_2291_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n29002), 
            .O(n6056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_6 (.CI(n29002), .I0(n2277), .I1(n96), .CO(n29003));
    SB_LUT4 add_2291_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n29001), 
            .O(n6057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_5 (.CI(n29001), .I0(n2278), .I1(n97), .CO(n29002));
    SB_LUT4 add_2291_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n29000), 
            .O(n6058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_4 (.CI(n29000), .I0(n2279), .I1(n98), .CO(n29001));
    SB_LUT4 add_2291_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n28999), 
            .O(n6059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_3 (.CI(n28999), .I0(n2280), .I1(n99), .CO(n29000));
    SB_LUT4 add_2291_2_lut (.I0(GND_net), .I1(n526), .I2(n558), .I3(VCC_net), 
            .O(n6060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2291_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2291_2 (.CI(VCC_net), .I0(n526), .I1(n558), .CO(n28999));
    SB_LUT4 add_2290_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n28998), 
            .O(n6024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2290_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n28997), 
            .O(n6025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_17 (.CI(n28997), .I0(n2169), .I1(n85), .CO(n28998));
    SB_LUT4 add_2290_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n28996), 
            .O(n6026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_16 (.CI(n28996), .I0(n2170), .I1(n86), .CO(n28997));
    SB_LUT4 add_2290_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n28995), 
            .O(n6027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_15 (.CI(n28995), .I0(n2171), .I1(n87), .CO(n28996));
    SB_LUT4 add_2290_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n28994), 
            .O(n6028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_14 (.CI(n28994), .I0(n2172), .I1(n88), .CO(n28995));
    SB_LUT4 add_2290_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n28993), 
            .O(n6029)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_13 (.CI(n28993), .I0(n2173), .I1(n89), .CO(n28994));
    SB_LUT4 add_2290_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n28992), 
            .O(n6030)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_12 (.CI(n28992), .I0(n2174), .I1(n90), .CO(n28993));
    SB_LUT4 add_2290_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n28991), 
            .O(n6031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_11 (.CI(n28991), .I0(n2175), .I1(n91), .CO(n28992));
    SB_LUT4 add_2290_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n28990), 
            .O(n6032)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_10 (.CI(n28990), .I0(n2176), .I1(n92), .CO(n28991));
    SB_LUT4 add_2290_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n28989), 
            .O(n6033)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_9 (.CI(n28989), .I0(n2177), .I1(n93), .CO(n28990));
    SB_LUT4 add_2290_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n28988), 
            .O(n6034)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_8 (.CI(n28988), .I0(n2178), .I1(n94), .CO(n28989));
    SB_LUT4 add_2290_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n28987), 
            .O(n6035)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_7 (.CI(n28987), .I0(n2179), .I1(n95), .CO(n28988));
    SB_LUT4 add_2290_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n28986), 
            .O(n6036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_6 (.CI(n28986), .I0(n2180), .I1(n96), .CO(n28987));
    SB_LUT4 add_2290_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n28985), 
            .O(n6037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_5 (.CI(n28985), .I0(n2181), .I1(n97), .CO(n28986));
    SB_LUT4 add_2290_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n28984), 
            .O(n6038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_4 (.CI(n28984), .I0(n2182), .I1(n98), .CO(n28985));
    SB_LUT4 add_2290_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n28983), 
            .O(n6039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_3 (.CI(n28983), .I0(n2183), .I1(n99), .CO(n28984));
    SB_LUT4 add_2290_2_lut (.I0(GND_net), .I1(n525), .I2(n558), .I3(VCC_net), 
            .O(n6040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2290_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2290_2 (.CI(VCC_net), .I0(n525), .I1(n558), .CO(n28983));
    SB_LUT4 add_2289_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n28982), 
            .O(n6006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2289_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n28981), 
            .O(n6007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_16 (.CI(n28981), .I0(n2070), .I1(n86), .CO(n28982));
    SB_LUT4 add_2289_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n28980), 
            .O(n6008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_15 (.CI(n28980), .I0(n2071), .I1(n87), .CO(n28981));
    SB_LUT4 add_2289_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n28979), 
            .O(n6009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_14 (.CI(n28979), .I0(n2072), .I1(n88), .CO(n28980));
    SB_LUT4 add_2289_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n28978), 
            .O(n6010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_13 (.CI(n28978), .I0(n2073), .I1(n89), .CO(n28979));
    SB_LUT4 add_2289_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n28977), 
            .O(n6011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_12 (.CI(n28977), .I0(n2074), .I1(n90), .CO(n28978));
    SB_LUT4 add_2289_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n28976), 
            .O(n6012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_11 (.CI(n28976), .I0(n2075), .I1(n91), .CO(n28977));
    SB_LUT4 add_2289_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n28975), 
            .O(n6013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_17 (.CI(n29345), .I0(n2944), .I1(n2966_adj_4400), 
            .CO(n29346));
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n29598), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_10 (.CI(n28975), .I0(n2076), .I1(n92), .CO(n28976));
    SB_LUT4 rem_4_add_1988_16_lut (.I0(n2945), .I1(n2945), .I2(n2966_adj_4400), 
            .I3(n29344), .O(n3044)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1988_16 (.CI(n29344), .I0(n2945), .I1(n2966_adj_4400), 
            .CO(n29345));
    SB_LUT4 add_2289_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n28974), 
            .O(n6014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_9 (.CI(n28974), .I0(n2077), .I1(n93), .CO(n28975));
    SB_LUT4 add_2289_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n28973), 
            .O(n6015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_15_lut (.I0(n2946), .I1(n2946), .I2(n2966_adj_4400), 
            .I3(n29343), .O(n3045)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_9 (.CI(n29598), .I0(n1952), .I1(VCC_net), 
            .CO(n29599));
    SB_CARRY add_2289_8 (.CI(n28973), .I0(n2078), .I1(n94), .CO(n28974));
    SB_LUT4 add_2289_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n28972), 
            .O(n6016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_7 (.CI(n28972), .I0(n2079), .I1(n95), .CO(n28973));
    SB_LUT4 add_2289_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n28971), 
            .O(n6017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_6 (.CI(n28971), .I0(n2080), .I1(n96), .CO(n28972));
    SB_CARRY rem_4_add_1988_15 (.CI(n29343), .I0(n2946), .I1(n2966_adj_4400), 
            .CO(n29344));
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n29597), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2289_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n28970), 
            .O(n6018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_3 (.CI(n28541), .I0(n1357), .I1(VCC_net), .CO(n28542));
    SB_CARRY add_2289_5 (.CI(n28970), .I0(n2081), .I1(n97), .CO(n28971));
    SB_LUT4 add_2289_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n28969), 
            .O(n6019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_4 (.CI(n28969), .I0(n2082), .I1(n98), .CO(n28970));
    SB_LUT4 rem_4_add_1988_14_lut (.I0(n2947), .I1(n2947), .I2(n2966_adj_4400), 
            .I3(n29342), .O(n3046)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_8 (.CI(n29597), .I0(n1953), .I1(VCC_net), 
            .CO(n29598));
    SB_LUT4 add_2289_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n28968), 
            .O(n6020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_3 (.CI(n28968), .I0(n2083), .I1(n99), .CO(n28969));
    SB_LUT4 add_2289_2_lut (.I0(GND_net), .I1(n524), .I2(n558), .I3(VCC_net), 
            .O(n6021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2289_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2289_2 (.CI(VCC_net), .I0(n524), .I1(n558), .CO(n28968));
    SB_CARRY rem_4_add_1988_14 (.CI(n29342), .I0(n2947), .I1(n2966_adj_4400), 
            .CO(n29343));
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n29596), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2288_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n28967), 
            .O(n5989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2288_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n28966), 
            .O(n5990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_13_lut (.I0(n2948), .I1(n2948), .I2(n2966_adj_4400), 
            .I3(n29341), .O(n3047)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_7 (.CI(n29596), .I0(n1954), .I1(GND_net), 
            .CO(n29597));
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n29595), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_13 (.CI(n29341), .I0(n2948), .I1(n2966_adj_4400), 
            .CO(n29342));
    SB_LUT4 rem_4_add_1988_12_lut (.I0(n2949_adj_4410), .I1(n2949_adj_4410), 
            .I2(n2966_adj_4400), .I3(n29340), .O(n3048)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_6 (.CI(n29595), .I0(n1955), .I1(GND_net), 
            .CO(n29596));
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n29594), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_15 (.CI(n28966), .I0(n1968), .I1(n87), .CO(n28967));
    SB_CARRY rem_4_add_1988_12 (.CI(n29340), .I0(n2949_adj_4410), .I1(n2966_adj_4400), 
            .CO(n29341));
    SB_LUT4 add_2288_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n28965), 
            .O(n5991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_11_lut (.I0(n2950_adj_4409), .I1(n2950_adj_4409), 
            .I2(n2966_adj_4400), .I3(n29339), .O(n3049)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_5 (.CI(n29594), .I0(n1956), .I1(VCC_net), 
            .CO(n29595));
    SB_CARRY add_2288_14 (.CI(n28965), .I0(n1969), .I1(n88), .CO(n28966));
    SB_LUT4 add_2288_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n28964), 
            .O(n5992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_13 (.CI(n28964), .I0(n1970), .I1(n89), .CO(n28965));
    SB_CARRY rem_4_add_1988_11 (.CI(n29339), .I0(n2950_adj_4409), .I1(n2966_adj_4400), 
            .CO(n29340));
    SB_LUT4 add_2288_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n28963), 
            .O(n5993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_12 (.CI(n28963), .I0(n1971), .I1(n90), .CO(n28964));
    SB_LUT4 add_2288_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n28962), 
            .O(n5994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_10_lut (.I0(n2951_adj_4408), .I1(n2951_adj_4408), 
            .I2(n2966_adj_4400), .I3(n29338), .O(n3050)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n29593), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_10 (.CI(n29338), .I0(n2951_adj_4408), .I1(n2966_adj_4400), 
            .CO(n29339));
    SB_CARRY rem_4_add_1318_4 (.CI(n29593), .I0(n1957), .I1(VCC_net), 
            .CO(n29594));
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(n29592), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_9_lut (.I0(n2952_adj_4407), .I1(n2952_adj_4407), 
            .I2(n2966_adj_4400), .I3(n29337), .O(n3051)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1318_3 (.CI(n29592), .I0(n1958), .I1(GND_net), 
            .CO(n29593));
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n2058), .I1(VCC_net), 
            .CO(n29592));
    SB_CARRY rem_4_add_1988_9 (.CI(n29337), .I0(n2952_adj_4407), .I1(n2966_adj_4400), 
            .CO(n29338));
    SB_LUT4 rem_4_add_1385_19_lut (.I0(n2075_adj_4599), .I1(n2042), .I2(VCC_net), 
            .I3(n29591), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_8_lut (.I0(n2953_adj_4406), .I1(n2953_adj_4406), 
            .I2(n2966_adj_4400), .I3(n29336), .O(n3052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1988_8 (.CI(n29336), .I0(n2953_adj_4406), .I1(n2966_adj_4400), 
            .CO(n29337));
    SB_LUT4 rem_4_add_1385_18_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n29590), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_7_lut (.I0(n2954_adj_4405), .I1(n2954_adj_4405), 
            .I2(n44233), .I3(n29335), .O(n3053)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_2288_11 (.CI(n28962), .I0(n1972), .I1(n91), .CO(n28963));
    SB_CARRY rem_4_add_1385_18 (.CI(n29590), .I0(n2043), .I1(VCC_net), 
            .CO(n29591));
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n29589), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_17 (.CI(n29589), .I0(n2044), .I1(VCC_net), 
            .CO(n29590));
    SB_CARRY rem_4_add_1988_7 (.CI(n29335), .I0(n2954_adj_4405), .I1(n44233), 
            .CO(n29336));
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n29588), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_6_lut (.I0(n2955_adj_4404), .I1(n2955_adj_4404), 
            .I2(n44233), .I3(n29334), .O(n3054)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_2288_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n28961), 
            .O(n5995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_10 (.CI(n28961), .I0(n1973), .I1(n92), .CO(n28962));
    SB_LUT4 i13180_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n35429), 
            .I3(GND_net), .O(n17925));   // verilog/coms.v(126[12] 289[6])
    defparam i13180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2288_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n28960), 
            .O(n5996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4784));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4785));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4786));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4789));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4779));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4781));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4782));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2288_9 (.CI(n28960), .I0(n1974), .I1(n93), .CO(n28961));
    SB_LUT4 add_2288_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n28959), 
            .O(n5997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_6 (.CI(n29334), .I0(n2955_adj_4404), .I1(n44233), 
            .CO(n29335));
    SB_CARRY add_2288_8 (.CI(n28959), .I0(n1975), .I1(n94), .CO(n28960));
    SB_LUT4 add_2288_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n28958), 
            .O(n5998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_7 (.CI(n28958), .I0(n1976), .I1(n95), .CO(n28959));
    SB_LUT4 add_2288_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n28957), 
            .O(n5999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_6 (.CI(n28957), .I0(n1977), .I1(n96), .CO(n28958));
    SB_LUT4 add_2288_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n28956), 
            .O(n6000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_5 (.CI(n28956), .I0(n1978), .I1(n97), .CO(n28957));
    SB_LUT4 add_2288_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n28955), 
            .O(n6001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_4 (.CI(n28955), .I0(n1979), .I1(n98), .CO(n28956));
    SB_LUT4 add_2288_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n28954), 
            .O(n6002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_3 (.CI(n28954), .I0(n1980), .I1(n99), .CO(n28955));
    SB_LUT4 add_2288_2_lut (.I0(GND_net), .I1(n523), .I2(n558), .I3(VCC_net), 
            .O(n6003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2288_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2288_2 (.CI(VCC_net), .I0(n523), .I1(n558), .CO(n28954));
    SB_LUT4 add_2287_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n28953), 
            .O(n5973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2287_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n28952), 
            .O(n5974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_14 (.CI(n28952), .I0(n1863), .I1(n88), .CO(n28953));
    SB_LUT4 add_2287_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n28951), 
            .O(n5975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_13 (.CI(n28951), .I0(n1864), .I1(n89), .CO(n28952));
    SB_LUT4 add_2287_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n28950), 
            .O(n5976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_12 (.CI(n28950), .I0(n1865), .I1(n90), .CO(n28951));
    SB_LUT4 add_2287_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n28949), 
            .O(n5977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_11 (.CI(n28949), .I0(n1866), .I1(n91), .CO(n28950));
    SB_LUT4 add_2287_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n28948), 
            .O(n5978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_10 (.CI(n28948), .I0(n1867), .I1(n92), .CO(n28949));
    SB_LUT4 add_2287_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n28947), 
            .O(n5979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_9 (.CI(n28947), .I0(n1868), .I1(n93), .CO(n28948));
    SB_LUT4 add_2287_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n28946), 
            .O(n5980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_8 (.CI(n28946), .I0(n1869), .I1(n94), .CO(n28947));
    SB_LUT4 add_2287_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n28945), 
            .O(n5981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_7 (.CI(n28945), .I0(n1870), .I1(n95), .CO(n28946));
    SB_LUT4 add_2287_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n28944), 
            .O(n5982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_6 (.CI(n28944), .I0(n1871), .I1(n96), .CO(n28945));
    SB_LUT4 add_2287_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n28943), 
            .O(n5983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_5 (.CI(n28943), .I0(n1872), .I1(n97), .CO(n28944));
    SB_LUT4 add_2287_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n28942), 
            .O(n5984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_4 (.CI(n28942), .I0(n1873), .I1(n98), .CO(n28943));
    SB_LUT4 add_2287_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n28941), 
            .O(n5985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_3 (.CI(n28941), .I0(n1874), .I1(n99), .CO(n28942));
    SB_LUT4 add_2287_2_lut (.I0(GND_net), .I1(n522), .I2(n558), .I3(VCC_net), 
            .O(n5986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2287_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2287_2 (.CI(VCC_net), .I0(n522), .I1(n558), .CO(n28941));
    SB_LUT4 add_2286_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n28940), 
            .O(n5958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2286_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n28939), 
            .O(n5959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_13 (.CI(n28939), .I0(n1755), .I1(n89), .CO(n28940));
    SB_LUT4 add_2286_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n28938), 
            .O(n5960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_12 (.CI(n28938), .I0(n1756), .I1(n90), .CO(n28939));
    SB_LUT4 add_2286_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n28937), 
            .O(n5961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_11 (.CI(n28937), .I0(n1757), .I1(n91), .CO(n28938));
    SB_LUT4 add_2286_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n28936), 
            .O(n5962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_10 (.CI(n28936), .I0(n1758), .I1(n92), .CO(n28937));
    SB_LUT4 add_2286_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n28935), 
            .O(n5963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_9 (.CI(n28935), .I0(n1759), .I1(n93), .CO(n28936));
    SB_LUT4 add_2286_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n28934), 
            .O(n5964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_8 (.CI(n28934), .I0(n1760), .I1(n94), .CO(n28935));
    SB_LUT4 add_2286_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n28933), 
            .O(n5965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_7 (.CI(n28933), .I0(n1761), .I1(n95), .CO(n28934));
    SB_LUT4 add_2286_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n28932), 
            .O(n5966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_6 (.CI(n28932), .I0(n1762), .I1(n96), .CO(n28933));
    SB_LUT4 add_2286_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n28931), 
            .O(n5967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_5 (.CI(n28931), .I0(n1763), .I1(n97), .CO(n28932));
    SB_LUT4 add_2286_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n28930), 
            .O(n5968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_4 (.CI(n28930), .I0(n1764), .I1(n98), .CO(n28931));
    SB_LUT4 add_2286_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n28929), 
            .O(n5969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_3 (.CI(n28929), .I0(n1765), .I1(n99), .CO(n28930));
    SB_LUT4 add_2286_2_lut (.I0(GND_net), .I1(n521), .I2(n558), .I3(VCC_net), 
            .O(n5970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2286_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2286_2 (.CI(VCC_net), .I0(n521), .I1(n558), .CO(n28929));
    SB_LUT4 add_2285_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n28928), 
            .O(n5944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2285_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n28927), 
            .O(n5945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_12 (.CI(n28927), .I0(n1644), .I1(n90), .CO(n28928));
    SB_LUT4 add_2285_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n28926), 
            .O(n5946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_11 (.CI(n28926), .I0(n1645), .I1(n91), .CO(n28927));
    SB_LUT4 add_2285_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n28925), 
            .O(n5947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_10 (.CI(n28925), .I0(n1646), .I1(n92), .CO(n28926));
    SB_LUT4 add_2285_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n28924), 
            .O(n5948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_9 (.CI(n28924), .I0(n1647), .I1(n93), .CO(n28925));
    SB_LUT4 add_2285_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n28923), 
            .O(n5949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_8 (.CI(n28923), .I0(n1648), .I1(n94), .CO(n28924));
    SB_LUT4 add_2285_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n28922), 
            .O(n5950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_7 (.CI(n28922), .I0(n1649), .I1(n95), .CO(n28923));
    SB_LUT4 add_2285_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n28921), 
            .O(n5951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_6 (.CI(n28921), .I0(n1650), .I1(n96), .CO(n28922));
    SB_LUT4 add_2285_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n28920), 
            .O(n5952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_5 (.CI(n28920), .I0(n1651), .I1(n97), .CO(n28921));
    SB_LUT4 add_2285_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n28919), 
            .O(n5953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_4 (.CI(n28919), .I0(n1652), .I1(n98), .CO(n28920));
    SB_LUT4 add_2285_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n28918), 
            .O(n5954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_3 (.CI(n28918), .I0(n1653), .I1(n99), .CO(n28919));
    SB_LUT4 add_2285_2_lut (.I0(GND_net), .I1(n520), .I2(n558), .I3(VCC_net), 
            .O(n5955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2285_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2285_2 (.CI(VCC_net), .I0(n520), .I1(n558), .CO(n28918));
    SB_LUT4 add_2284_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n28917), 
            .O(n5931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2284_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n28916), 
            .O(n5932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_11 (.CI(n28916), .I0(n1530), .I1(n91), .CO(n28917));
    SB_LUT4 add_2284_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n28915), 
            .O(n5933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_10 (.CI(n28915), .I0(n1531), .I1(n92), .CO(n28916));
    SB_LUT4 add_2284_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n28914), 
            .O(n5934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_9 (.CI(n28914), .I0(n1532), .I1(n93), .CO(n28915));
    SB_LUT4 add_2284_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n28913), 
            .O(n5935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_8 (.CI(n28913), .I0(n1533), .I1(n94), .CO(n28914));
    SB_LUT4 add_2284_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n28912), 
            .O(n5936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_7 (.CI(n28912), .I0(n1534), .I1(n95), .CO(n28913));
    SB_LUT4 add_2284_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n28911), 
            .O(n5937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_6 (.CI(n28911), .I0(n1535), .I1(n96), .CO(n28912));
    SB_LUT4 add_2284_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n28910), 
            .O(n5938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_5 (.CI(n28910), .I0(n1536), .I1(n97), .CO(n28911));
    SB_LUT4 add_2284_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n28909), 
            .O(n5939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35383_3_lut (.I0(n2253), .I1(n2320), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35384_3_lut (.I0(n2352), .I1(n2419), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2451_adj_4571));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35384_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2284_4 (.CI(n28909), .I0(n1537), .I1(n98), .CO(n28910));
    SB_LUT4 add_2284_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n28908), 
            .O(n5940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_3 (.CI(n28908), .I0(n1538), .I1(n99), .CO(n28909));
    SB_LUT4 add_2284_2_lut (.I0(GND_net), .I1(n519), .I2(n558), .I3(VCC_net), 
            .O(n5941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2284_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2284_2 (.CI(VCC_net), .I0(n519), .I1(n558), .CO(n28908));
    SB_LUT4 add_2283_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n28907), 
            .O(n5919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2283_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n28906), 
            .O(n5920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_10 (.CI(n28906), .I0(n1413), .I1(n92), .CO(n28907));
    SB_LUT4 add_2283_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n28905), 
            .O(n5921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_9 (.CI(n28905), .I0(n1414), .I1(n93), .CO(n28906));
    SB_LUT4 add_2283_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n28904), 
            .O(n5922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_8 (.CI(n28904), .I0(n1415), .I1(n94), .CO(n28905));
    SB_LUT4 add_2283_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n28903), 
            .O(n5923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_7 (.CI(n28903), .I0(n1416), .I1(n95), .CO(n28904));
    SB_LUT4 add_2283_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n28902), 
            .O(n5924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_6 (.CI(n28902), .I0(n1417), .I1(n96), .CO(n28903));
    SB_LUT4 add_2283_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n28901), 
            .O(n5925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_5 (.CI(n28901), .I0(n1418), .I1(n97), .CO(n28902));
    SB_LUT4 add_2283_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n28900), 
            .O(n5926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_4 (.CI(n28900), .I0(n1419), .I1(n98), .CO(n28901));
    SB_LUT4 add_2283_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n28899), 
            .O(n5927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_3 (.CI(n28899), .I0(n1420), .I1(n99), .CO(n28900));
    SB_LUT4 add_2283_2_lut (.I0(GND_net), .I1(n518), .I2(n558), .I3(VCC_net), 
            .O(n5928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2283_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2283_2 (.CI(VCC_net), .I0(n518), .I1(n558), .CO(n28899));
    SB_LUT4 add_2282_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n28898), 
            .O(n5908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2282_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n28897), 
            .O(n5909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2282_9 (.CI(n28897), .I0(n1293), .I1(n93), .CO(n28898));
    SB_LUT4 add_2282_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n28896), 
            .O(n5910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2282_8 (.CI(n28896), .I0(n1294), .I1(n94), .CO(n28897));
    SB_LUT4 add_2282_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n28895), 
            .O(n5911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2282_7 (.CI(n28895), .I0(n1295), .I1(n95), .CO(n28896));
    SB_LUT4 i34552_4_lut (.I0(n33_adj_4789), .I1(n21_adj_4782), .I2(n19_adj_4781), 
            .I3(n17_adj_4779), .O(n41405));
    defparam i34552_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35291_4_lut (.I0(n15_adj_4777), .I1(n13_adj_4775), .I2(n2552), 
            .I3(n98), .O(n42145));
    defparam i35291_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i35832_4_lut (.I0(n21_adj_4782), .I1(n19_adj_4781), .I2(n17_adj_4779), 
            .I3(n42145), .O(n42686));
    defparam i35832_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35830_4_lut (.I0(n27_adj_4786), .I1(n25_adj_4785), .I2(n23_adj_4784), 
            .I3(n42686), .O(n42684));
    defparam i35830_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34556_4_lut (.I0(n33_adj_4789), .I1(n31_adj_4788), .I2(n29_adj_4787), 
            .I3(n42684), .O(n41409));
    defparam i34556_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2282_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n28894), 
            .O(n5912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_5_lut (.I0(n2956_adj_4403), .I1(n2956_adj_4403), 
            .I2(n2966_adj_4400), .I3(n29333), .O(n3055)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2282_6 (.CI(n28894), .I0(n1296), .I1(n96), .CO(n28895));
    SB_LUT4 div_46_LessThan_1665_i10_4_lut (.I0(n529), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4773));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540_adj_4511), .I1(n2607), .I2(n2570), 
            .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36282_3_lut (.I0(n10_adj_4773), .I1(n87), .I2(n33_adj_4789), 
            .I3(GND_net), .O(n43136));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36282_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36283_3_lut (.I0(n43136), .I1(n86), .I2(n35_adj_4790), .I3(GND_net), 
            .O(n43137));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36283_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2282_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n28893), 
            .O(n5913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_16 (.CI(n29588), .I0(n2045), .I1(VCC_net), 
            .CO(n29589));
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n29587), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n29333), .I0(n2956_adj_4403), .I1(n2966_adj_4400), 
            .CO(n29334));
    SB_CARRY add_2282_5 (.CI(n28893), .I0(n1297), .I1(n97), .CO(n28894));
    SB_CARRY rem_4_add_1385_15 (.CI(n29587), .I0(n2046), .I1(VCC_net), 
            .CO(n29588));
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n29586), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_4_lut (.I0(n2957_adj_4402), .I1(n2957_adj_4402), 
            .I2(n2966_adj_4400), .I3(n29332), .O(n3056)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_1665_i36_3_lut (.I0(n18_adj_4780), .I1(n83), 
            .I2(n41_adj_4794), .I3(GND_net), .O(n36_adj_4791));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34544_4_lut (.I0(n39_adj_4793), .I1(n37_adj_4792), .I2(n35_adj_4790), 
            .I3(n41405), .O(n41397));
    defparam i34544_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36531_4_lut (.I0(n36_adj_4791), .I1(n16_adj_4778), .I2(n41_adj_4794), 
            .I3(n41393), .O(n43385));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36531_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36162_3_lut (.I0(n43137), .I1(n85), .I2(n37_adj_4792), .I3(GND_net), 
            .O(n43016));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36162_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2282_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n28892), 
            .O(n5914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_4 (.CI(n29332), .I0(n2957_adj_4402), .I1(n2966_adj_4400), 
            .CO(n29333));
    SB_CARRY rem_4_add_1385_14 (.CI(n29586), .I0(n2047), .I1(VCC_net), 
            .CO(n29587));
    SB_LUT4 rem_4_add_1988_3_lut (.I0(n2958_adj_4401), .I1(n2958_adj_4401), 
            .I2(n44233), .I3(n29331), .O(n3057)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_2282_4 (.CI(n28892), .I0(n1298), .I1(n98), .CO(n28893));
    SB_LUT4 div_46_LessThan_1665_i22_3_lut (.I0(n14_adj_4776), .I1(n91), 
            .I2(n25_adj_4785), .I3(GND_net), .O(n22_adj_4783));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36529_4_lut (.I0(n22_adj_4783), .I1(n12_adj_4774), .I2(n25_adj_4785), 
            .I3(n41423), .O(n43383));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36529_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36530_3_lut (.I0(n43383), .I1(n90), .I2(n27_adj_4786), .I3(GND_net), 
            .O(n43384));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36530_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36441_3_lut (.I0(n43384), .I1(n89), .I2(n29_adj_4787), .I3(GND_net), 
            .O(n43295));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36441_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36050_4_lut (.I0(n39_adj_4793), .I1(n37_adj_4792), .I2(n35_adj_4790), 
            .I3(n41409), .O(n42904));
    defparam i36050_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36604_4_lut (.I0(n43016), .I1(n43385), .I2(n41_adj_4794), 
            .I3(n41397), .O(n43458));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36604_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36373_3_lut (.I0(n43295), .I1(n88), .I2(n31_adj_4788), .I3(GND_net), 
            .O(n43227));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36373_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36622_4_lut (.I0(n43227), .I1(n43458), .I2(n41_adj_4794), 
            .I3(n42904), .O(n43476));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36622_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36623_3_lut (.I0(n43476), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n43477));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36623_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_2282_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n28891), 
            .O(n5915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2282_3 (.CI(n28891), .I0(n1299), .I1(n99), .CO(n28892));
    SB_LUT4 i36619_3_lut (.I0(n43477), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n43473));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36619_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n43473), .I1(n16001), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4469), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_rep_75_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), 
            .I3(GND_net), .O(n1356));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i858_rep_75_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2282_2_lut (.I0(GND_net), .I1(n517), .I2(n558), .I3(VCC_net), 
            .O(n5916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2282_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n29331), .I0(n2958_adj_4401), .I1(n44233), 
            .CO(n29332));
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647_adj_4463), .I1(n1714), .I2(n1679), 
            .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4769));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2282_2 (.CI(VCC_net), .I0(n517), .I1(n558), .CO(n28891));
    SB_LUT4 add_2281_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n28890), 
            .O(n5898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2281_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n28889), 
            .O(n5899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4767));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4771));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4770));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4336), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n528));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4764));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4765));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1699 (.I0(n24670), .I1(n1766), .I2(GND_net), 
            .I3(GND_net), .O(n38531));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_2_lut_adj_1699.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4752));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4754));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2281_8 (.CI(n28889), .I0(n1170), .I1(n94), .CO(n28890));
    SB_LUT4 div_46_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4761));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4762));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(color_23__N_164[7]), .I1(n11_adj_4490), 
            .I2(color_23__N_164[1]), .I3(n38531), .O(n38537));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4763));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i29528_4_lut (.I0(n38537), .I1(n17240), .I2(color[1]), .I3(n13_adj_4489), 
            .O(n36299));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i29528_4_lut.LUT_INIT = 16'hc0c4;
    SB_LUT4 i13366_3_lut (.I0(n17321), .I1(r_Bit_Index[0]), .I2(n17180), 
            .I3(GND_net), .O(n18111));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13366_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i13181_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n35429), 
            .I3(GND_net), .O(n17926));   // verilog/coms.v(126[12] 289[6])
    defparam i13181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1607_3_lut (.I0(n2358_adj_4578), .I1(n2425), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2457_adj_4517));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2454_adj_4568));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1701 (.I0(n17240), .I1(color[4]), .I2(n36415), 
            .I3(GND_net), .O(n32662));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1701.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_1702 (.I0(n2439), .I1(n2438), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4889));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i1_2_lut_adj_1702.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1703 (.I0(n2456_adj_4518), .I1(n2458_adj_4516), 
            .I2(GND_net), .I3(GND_net), .O(n38945));
    defparam i1_2_lut_adj_1703.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n2454_adj_4568), .I1(n38945), .I2(n2455_adj_4567), 
            .I3(n2457_adj_4517), .O(n36550));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut_adj_1705 (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n38783));
    defparam i1_2_lut_adj_1705.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4766));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1706 (.I0(n17240), .I1(color[3]), .I2(n36415), 
            .I3(GND_net), .O(n32660));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1706.LUT_INIT = 16'ha8a8;
    SB_LUT4 add_2281_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n28888), 
            .O(n5900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13386_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1144), .I3(GND_net), .O(n18131));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1707 (.I0(n2451_adj_4571), .I1(n2453_adj_4569), 
            .I2(n2450_adj_4572), .I3(n18_adj_4889), .O(n30_adj_4885));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1708 (.I0(n2444), .I1(n2445), .I2(n36550), .I3(n2446), 
            .O(n28_adj_4887));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1709 (.I0(n2449_adj_4573), .I1(n2447_adj_4575), 
            .I2(n2448_adj_4574), .I3(n2452_adj_4570), .O(n29_adj_4886));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1710 (.I0(n2440), .I1(n2442), .I2(n2441), .I3(n2443), 
            .O(n27_adj_4888));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n1854), .I1(n38783), .I2(n1855), .I3(n1857), 
            .O(n36480));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'ha080;
    SB_LUT4 i16_4_lut_adj_1712 (.I0(n27_adj_4888), .I1(n29_adj_4886), .I2(n28_adj_4887), 
            .I3(n30_adj_4885), .O(n2471_adj_4515));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i16_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372_adj_4577), 
            .I3(GND_net), .O(n2455_adj_4567));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1713 (.I0(n1846), .I1(n36480), .I2(n1847), .I3(n1848), 
            .O(n18_adj_4331));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i7_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_CARRY add_2281_7 (.CI(n28888), .I0(n1171), .I1(n95), .CO(n28889));
    SB_LUT4 rem_4_i1672_3_lut (.I0(n2455_adj_4567), .I1(n2522), .I2(n2471_adj_4515), 
            .I3(GND_net), .O(n2554));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_2_lut (.I0(n1851), .I1(n1853), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4332));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4756));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4758));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1714 (.I0(n17240), .I1(color[20]), .I2(n36429), 
            .I3(GND_net), .O(n32680));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1714.LUT_INIT = 16'h8a8a;
    SB_LUT4 i9_4_lut_adj_1715 (.I0(n1852), .I1(n18_adj_4331), .I2(n1845), 
            .I3(n1844), .O(n20_adj_4330));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i9_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2281_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n28887), 
            .O(n5901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n3058), .I1(VCC_net), 
            .CO(n29331));
    SB_LUT4 div_46_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4759));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10_4_lut_adj_1716 (.I0(n1849), .I1(n20_adj_4330), .I2(n16_adj_4332), 
            .I3(n1850), .O(n1877));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i13312_3_lut (.I0(encoder0_position[8]), .I1(n3014), .I2(count_enable), 
            .I3(GND_net), .O(n18057));   // quad.v(35[10] 41[6])
    defparam i13312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13311_3_lut (.I0(encoder0_position[7]), .I1(n3015), .I2(count_enable), 
            .I3(GND_net), .O(n18056));   // quad.v(35[10] 41[6])
    defparam i13311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34622_4_lut (.I0(n35_adj_4766), .I1(n23_adj_4759), .I2(n21_adj_4758), 
            .I3(n19_adj_4756), .O(n41475));
    defparam i34622_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2281_6 (.CI(n28887), .I0(n1172), .I1(n96), .CO(n28888));
    SB_LUT4 i35367_4_lut (.I0(n17_adj_4754), .I1(n15_adj_4752), .I2(n2464), 
            .I3(n98), .O(n42221));
    defparam i35367_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 add_2281_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n28886), 
            .O(n5902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2281_5 (.CI(n28886), .I0(n1173), .I1(n97), .CO(n28887));
    SB_LUT4 add_2281_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n28885), 
            .O(n5903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1717 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n36465));
    defparam i1_3_lut_adj_1717.LUT_INIT = 16'hfefe;
    SB_CARRY add_2281_4 (.CI(n28885), .I0(n1174), .I1(n98), .CO(n28886));
    SB_LUT4 i35850_4_lut (.I0(n23_adj_4759), .I1(n21_adj_4758), .I2(n19_adj_4756), 
            .I3(n42221), .O(n42704));
    defparam i35850_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35848_4_lut (.I0(n29_adj_4763), .I1(n27_adj_4762), .I2(n25_adj_4761), 
            .I3(n42704), .O(n42702));
    defparam i35848_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34624_4_lut (.I0(n35_adj_4766), .I1(n33_adj_4765), .I2(n31_adj_4764), 
            .I3(n42702), .O(n41477));
    defparam i34624_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1606_i12_4_lut (.I0(n528), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4750));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36290_3_lut (.I0(n12_adj_4750), .I1(n87), .I2(n35_adj_4766), 
            .I3(GND_net), .O(n43144));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36290_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2281_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n28884), 
            .O(n5904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2281_3 (.CI(n28884), .I0(n1175), .I1(n99), .CO(n28885));
    SB_LUT4 rem_4_add_916_2_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(VCC_net), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2281_2_lut (.I0(GND_net), .I1(n516), .I2(n558), .I3(VCC_net), 
            .O(n5905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2281_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2281_2 (.CI(VCC_net), .I0(n516), .I1(n558), .CO(n28884));
    SB_LUT4 div_46_LessThan_1606_i38_3_lut (.I0(n20_adj_4757), .I1(n83), 
            .I2(n43_adj_4771), .I3(GND_net), .O(n38_adj_4768));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36291_3_lut (.I0(n43144), .I1(n86), .I2(n37_adj_4767), .I3(GND_net), 
            .O(n43145));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36291_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34617_4_lut (.I0(n41_adj_4770), .I1(n39_adj_4769), .I2(n37_adj_4767), 
            .I3(n41475), .O(n41470));
    defparam i34617_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36288_4_lut (.I0(n38_adj_4768), .I1(n18_adj_4755), .I2(n43_adj_4771), 
            .I3(n41466), .O(n43142));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36288_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2280_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n28883), 
            .O(n5889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2280_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n28882), 
            .O(n5890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_7 (.CI(n28882), .I0(n1044), .I1(n95), .CO(n28883));
    SB_LUT4 i36156_3_lut (.I0(n43145), .I1(n85), .I2(n39_adj_4769), .I3(GND_net), 
            .O(n43010));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36156_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1606_i24_3_lut (.I0(n16_adj_4753), .I1(n91), 
            .I2(n27_adj_4762), .I3(GND_net), .O(n24_adj_4760));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36525_4_lut (.I0(n24_adj_4760), .I1(n14_adj_4751), .I2(n27_adj_4762), 
            .I3(n41493), .O(n43379));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36525_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36526_3_lut (.I0(n43379), .I1(n90), .I2(n29_adj_4763), .I3(GND_net), 
            .O(n43380));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36526_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36443_3_lut (.I0(n43380), .I1(n89), .I2(n31_adj_4764), .I3(GND_net), 
            .O(n43297));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36443_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2280_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n28881), 
            .O(n5891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n29585), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_6 (.CI(n28881), .I0(n1045), .I1(n96), .CO(n28882));
    SB_LUT4 rem_4_add_2055_29_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n29330), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1385_13 (.CI(n29585), .I0(n2048), .I1(VCC_net), 
            .CO(n29586));
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n29584), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_28_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n29329), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_12 (.CI(n29584), .I0(n2049), .I1(VCC_net), 
            .CO(n29585));
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n29583), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_11 (.CI(n29583), .I0(n2050), .I1(VCC_net), 
            .CO(n29584));
    SB_LUT4 add_2280_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n28880), 
            .O(n5892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_5 (.CI(n28880), .I0(n1046), .I1(n97), .CO(n28881));
    SB_LUT4 add_2280_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n28879), 
            .O(n5893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_4 (.CI(n28879), .I0(n1047), .I1(n98), .CO(n28880));
    SB_LUT4 i36070_4_lut (.I0(n41_adj_4770), .I1(n39_adj_4769), .I2(n37_adj_4767), 
            .I3(n41477), .O(n42924));
    defparam i36070_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2280_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n28878), 
            .O(n5894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_3 (.CI(n28878), .I0(n1048), .I1(n99), .CO(n28879));
    SB_LUT4 i36508_4_lut (.I0(n43010), .I1(n43142), .I2(n43_adj_4771), 
            .I3(n41470), .O(n43362));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36508_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1358), .I1(GND_net), 
            .CO(n28541));
    SB_LUT4 add_2280_2_lut (.I0(GND_net), .I1(n515), .I2(n558), .I3(VCC_net), 
            .O(n5895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2280_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2280_2 (.CI(VCC_net), .I0(n515), .I1(n558), .CO(n28878));
    SB_LUT4 i36371_3_lut (.I0(n43297), .I1(n88), .I2(n33_adj_4765), .I3(GND_net), 
            .O(n43225));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36371_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2279_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n28877), 
            .O(n5881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2279_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n28876), 
            .O(n5882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2279_6 (.CI(n28876), .I0(n915), .I1(n96), .CO(n28877));
    SB_LUT4 add_2279_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n28875), 
            .O(n5883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2279_5 (.CI(n28875), .I0(n916), .I1(n97), .CO(n28876));
    SB_LUT4 i36610_4_lut (.I0(n43225), .I1(n43362), .I2(n43_adj_4771), 
            .I3(n42924), .O(n43464));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36610_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36611_3_lut (.I0(n43464), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n43465));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36611_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n29582), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_28 (.CI(n29329), .I0(n3033), .I1(VCC_net), 
            .CO(n29330));
    SB_LUT4 add_2279_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n28874), 
            .O(n5884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2279_4 (.CI(n28874), .I0(n917), .I1(n98), .CO(n28875));
    SB_LUT4 add_2279_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n28873), 
            .O(n5885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_10 (.CI(n29582), .I0(n2051), .I1(VCC_net), 
            .CO(n29583));
    SB_CARRY add_2279_3 (.CI(n28873), .I0(n918), .I1(n99), .CO(n28874));
    SB_LUT4 add_2279_2_lut (.I0(GND_net), .I1(n514), .I2(n558), .I3(VCC_net), 
            .O(n5886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2279_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13388_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1144), .I3(GND_net), .O(n18133));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n43465), .I1(n15998), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n29328), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2279_2 (.CI(VCC_net), .I0(n514), .I1(n558), .CO(n28873));
    SB_LUT4 rem_4_add_648_7_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n28872), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2055_27 (.CI(n29328), .I0(n3034), .I1(VCC_net), 
            .CO(n29329));
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n29581), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_9 (.CI(n29581), .I0(n2052), .I1(VCC_net), 
            .CO(n29582));
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n29327), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n28871), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_26 (.CI(n29327), .I0(n3035), .I1(VCC_net), 
            .CO(n29328));
    SB_CARRY rem_4_add_648_6 (.CI(n28871), .I0(n954), .I1(GND_net), .CO(n28872));
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n29580), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_8 (.CI(n29580), .I0(n2053), .I1(VCC_net), 
            .CO(n29581));
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n29579), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n29326), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958_adj_4401));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_25 (.CI(n29326), .I0(n3036), .I1(VCC_net), 
            .CO(n29327));
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n28870), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_7 (.CI(n29579), .I0(n2054), .I1(GND_net), 
            .CO(n29580));
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n29325), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_5 (.CI(n28870), .I0(n955), .I1(GND_net), .CO(n28871));
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n28869), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_4 (.CI(n28869), .I0(n956), .I1(VCC_net), .CO(n28870));
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n28868), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n29578), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_3 (.CI(n28868), .I0(n957), .I1(VCC_net), .CO(n28869));
    SB_LUT4 rem_4_add_782_9_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n28540), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2055_24 (.CI(n29325), .I0(n3037), .I1(VCC_net), 
            .CO(n29326));
    SB_LUT4 rem_4_add_648_2_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(VCC_net), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n29324), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n958), .I1(GND_net), .CO(n28868));
    SB_CARRY rem_4_add_1385_6 (.CI(n29578), .I0(n2055), .I1(GND_net), 
            .CO(n29579));
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n29577), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_5 (.CI(n29577), .I0(n2056), .I1(VCC_net), 
            .CO(n29578));
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n29576), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_4 (.CI(n29576), .I0(n2057), .I1(VCC_net), 
            .CO(n29577));
    SB_CARRY rem_4_add_2055_23 (.CI(n29324), .I0(n3038), .I1(VCC_net), 
            .CO(n29325));
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n29323), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_22 (.CI(n29323), .I0(n3039), .I1(VCC_net), 
            .CO(n29324));
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(n29575), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n29322), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n28539), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4747));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1385_3 (.CI(n29575), .I0(n2058), .I1(GND_net), 
            .CO(n29576));
    SB_CARRY rem_4_add_2055_21 (.CI(n29322), .I0(n3040), .I1(VCC_net), 
            .CO(n29323));
    SB_LUT4 i13387_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1144), .I3(GND_net), .O(n18132));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13387_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2158), .I1(VCC_net), 
            .CO(n29575));
    SB_CARRY rem_4_add_782_8 (.CI(n28539), .I0(n1152), .I1(VCC_net), .CO(n28540));
    SB_LUT4 i13390_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1144), .I3(GND_net), .O(n18135));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n29321), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_20_lut (.I0(n2174_adj_4589), .I1(n2141), .I2(VCC_net), 
            .I3(n29574), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2055_20 (.CI(n29321), .I0(n3041), .I1(VCC_net), 
            .CO(n29322));
    SB_LUT4 rem_4_add_1452_19_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n29573), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_19 (.CI(n29573), .I0(n2142), .I1(VCC_net), 
            .CO(n29574));
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n29320), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1199__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_LUT4 div_46_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4749));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2055_19 (.CI(n29320), .I0(n3042), .I1(VCC_net), 
            .CO(n29321));
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n29572), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n29319), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_18 (.CI(n29572), .I0(n2143), .I1(VCC_net), 
            .CO(n29573));
    SB_LUT4 div_46_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4745));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n29571), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_18 (.CI(n29319), .I0(n3043), .I1(VCC_net), 
            .CO(n29320));
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n29318), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_17 (.CI(n29571), .I0(n2144), .I1(VCC_net), 
            .CO(n29572));
    SB_CARRY rem_4_add_2055_17 (.CI(n29318), .I0(n3044), .I1(VCC_net), 
            .CO(n29319));
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n28538), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n29317), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n29570), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_16 (.CI(n29570), .I0(n2145), .I1(VCC_net), 
            .CO(n29571));
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n29569), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_15 (.CI(n29569), .I0(n2146), .I1(VCC_net), 
            .CO(n29570));
    SB_CARRY rem_4_add_2055_16 (.CI(n29317), .I0(n3045), .I1(VCC_net), 
            .CO(n29318));
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n29568), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4335), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n527));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n29316), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_14 (.CI(n29568), .I0(n2147), .I1(VCC_net), 
            .CO(n29569));
    SB_CARRY rem_4_add_2055_15 (.CI(n29316), .I0(n3046), .I1(VCC_net), 
            .CO(n29317));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n29315), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_7 (.CI(n28538), .I0(n1153), .I1(VCC_net), .CO(n28539));
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n29567), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_13 (.CI(n29567), .I0(n2148), .I1(VCC_net), 
            .CO(n29568));
    SB_CARRY rem_4_add_2055_14 (.CI(n29315), .I0(n3047), .I1(VCC_net), 
            .CO(n29316));
    SB_DFF communication_counter_1199__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_DFF communication_counter_1199__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(76[28:51])
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n29566), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n29314), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_12 (.CI(n29566), .I0(n2149), .I1(VCC_net), 
            .CO(n29567));
    SB_LUT4 div_46_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4739));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2055_13 (.CI(n29314), .I0(n3048), .I1(VCC_net), 
            .CO(n29315));
    SB_LUT4 i13389_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1144), .I3(GND_net), .O(n18134));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n29565), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4740));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n29313), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_11 (.CI(n29565), .I0(n2150), .I1(VCC_net), 
            .CO(n29566));
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n29564), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_12 (.CI(n29313), .I0(n3049), .I1(VCC_net), 
            .CO(n29314));
    SB_CARRY rem_4_add_1452_10 (.CI(n29564), .I0(n2151), .I1(VCC_net), 
            .CO(n29565));
    SB_LUT4 div_46_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4741));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n29312), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n29563), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_11 (.CI(n29312), .I0(n3050), .I1(VCC_net), 
            .CO(n29313));
    SB_LUT4 i13392_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1144), .I3(GND_net), .O(n18137));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13392_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_9 (.CI(n29563), .I0(n2152), .I1(VCC_net), 
            .CO(n29564));
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n29311), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4748));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n29562), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1719 (.I0(n1947), .I1(n1954), .I2(n36465), .I3(n1955), 
            .O(n15_adj_4985));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i3_4_lut_adj_1719.LUT_INIT = 16'heaaa;
    SB_CARRY rem_4_add_1452_8 (.CI(n29562), .I0(n2153), .I1(VCC_net), 
            .CO(n29563));
    SB_CARRY rem_4_add_2055_10 (.CI(n29311), .I0(n3051), .I1(VCC_net), 
            .CO(n29312));
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n29561), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n29310), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n28537), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_7 (.CI(n29561), .I0(n2154), .I1(GND_net), 
            .CO(n29562));
    SB_CARRY rem_4_add_2055_9 (.CI(n29310), .I0(n3052), .I1(VCC_net), 
            .CO(n29311));
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n29560), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_6 (.CI(n29560), .I0(n2155), .I1(GND_net), 
            .CO(n29561));
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n29309), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n29559), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_5 (.CI(n29559), .I0(n2156), .I1(VCC_net), 
            .CO(n29560));
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n29558), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_4 (.CI(n29558), .I0(n2157), .I1(VCC_net), 
            .CO(n29559));
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(n29557), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_3 (.CI(n29557), .I0(n2158), .I1(GND_net), 
            .CO(n29558));
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2258), .I1(VCC_net), 
            .CO(n29557));
    SB_LUT4 rem_4_add_1519_21_lut (.I0(n2273_adj_4581), .I1(n2240), .I2(VCC_net), 
            .I3(n29556), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1519_20_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n29555), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_20 (.CI(n29555), .I0(n2241), .I1(VCC_net), 
            .CO(n29556));
    SB_CARRY rem_4_add_2055_8 (.CI(n29309), .I0(n3053), .I1(VCC_net), 
            .CO(n29310));
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n29554), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n29308), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4730));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_782_6 (.CI(n28537), .I0(n1154), .I1(GND_net), .CO(n28538));
    SB_CARRY rem_4_add_2055_7 (.CI(n29308), .I0(n3054), .I1(GND_net), 
            .CO(n29309));
    SB_CARRY rem_4_add_1519_19 (.CI(n29554), .I0(n2242), .I1(VCC_net), 
            .CO(n29555));
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n29553), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n29307), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_18 (.CI(n29553), .I0(n2243), .I1(VCC_net), 
            .CO(n29554));
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n29552), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_17 (.CI(n29552), .I0(n2244), .I1(VCC_net), 
            .CO(n29553));
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n29551), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n28536), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_16 (.CI(n29551), .I0(n2245), .I1(VCC_net), 
            .CO(n29552));
    SB_CARRY rem_4_add_2055_6 (.CI(n29307), .I0(n3055), .I1(GND_net), 
            .CO(n29308));
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n29550), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_15 (.CI(n29550), .I0(n2246), .I1(VCC_net), 
            .CO(n29551));
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n29306), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_5 (.CI(n29306), .I0(n3056), .I1(VCC_net), 
            .CO(n29307));
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n29549), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_14 (.CI(n29549), .I0(n2247), .I1(VCC_net), 
            .CO(n29550));
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n29305), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n29548), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_13 (.CI(n29548), .I0(n2248), .I1(VCC_net), 
            .CO(n29549));
    SB_CARRY rem_4_add_2055_4 (.CI(n29305), .I0(n3057), .I1(VCC_net), 
            .CO(n29306));
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n29547), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_12 (.CI(n29547), .I0(n2249), .I1(VCC_net), 
            .CO(n29548));
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n29546), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_11 (.CI(n29546), .I0(n2250), .I1(VCC_net), 
            .CO(n29547));
    SB_LUT4 div_46_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4732));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(n29304), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4734));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_782_5 (.CI(n28536), .I0(n1155), .I1(GND_net), .CO(n28537));
    SB_LUT4 div_46_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4736));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n29545), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4737));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2055_3 (.CI(n29304), .I0(n3058), .I1(GND_net), 
            .CO(n29305));
    SB_LUT4 div_46_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4742));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3158), .I1(VCC_net), 
            .CO(n29304));
    SB_CARRY rem_4_add_1519_10 (.CI(n29545), .I0(n2251), .I1(VCC_net), 
            .CO(n29546));
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n29544), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4743));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4744));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1519_9 (.CI(n29544), .I0(n2252), .I1(VCC_net), 
            .CO(n29545));
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n29543), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_8 (.CI(n29543), .I0(n2253), .I1(VCC_net), 
            .CO(n29544));
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n29542), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34708_4_lut (.I0(n37_adj_4744), .I1(n25_adj_4737), .I2(n23_adj_4736), 
            .I3(n21_adj_4734), .O(n41561));
    defparam i34708_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1519_7 (.CI(n29542), .I0(n2254), .I1(GND_net), 
            .CO(n29543));
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n29541), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_6 (.CI(n29541), .I0(n2255), .I1(GND_net), 
            .CO(n29542));
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n29540), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_5 (.CI(n29540), .I0(n2256), .I1(VCC_net), 
            .CO(n29541));
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n29539), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_4 (.CI(n29539), .I0(n2257), .I1(VCC_net), 
            .CO(n29540));
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(n29538), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13391_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1144), .I3(GND_net), .O(n18136));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13391_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_3 (.CI(n29538), .I0(n2258), .I1(GND_net), 
            .CO(n29539));
    SB_LUT4 rem_4_add_715_8_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n28813), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4578), .I1(VCC_net), 
            .CO(n29538));
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n28812), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_22_lut (.I0(n2372_adj_4577), .I1(n2339), .I2(VCC_net), 
            .I3(n29537), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1586_21_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n29536), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35503_4_lut (.I0(n19_adj_4732), .I1(n17_adj_4730), .I2(n2373), 
            .I3(n98), .O(n42357));
    defparam i35503_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY rem_4_add_715_7 (.CI(n28812), .I0(n1053), .I1(VCC_net), .CO(n28813));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n28811), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_6 (.CI(n28811), .I0(n1054), .I1(GND_net), .CO(n28812));
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n28535), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35902_4_lut (.I0(n25_adj_4737), .I1(n23_adj_4736), .I2(n21_adj_4734), 
            .I3(n42357), .O(n42756));
    defparam i35902_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY rem_4_add_1586_21 (.CI(n29536), .I0(n2340), .I1(VCC_net), 
            .CO(n29537));
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n29535), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35898_4_lut (.I0(n31_adj_4741), .I1(n29_adj_4740), .I2(n27_adj_4739), 
            .I3(n42756), .O(n42752));
    defparam i35898_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n28810), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_20 (.CI(n29535), .I0(n2341), .I1(VCC_net), 
            .CO(n29536));
    SB_CARRY rem_4_add_715_5 (.CI(n28810), .I0(n1055), .I1(GND_net), .CO(n28811));
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n28809), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_4 (.CI(n28809), .I0(n1056), .I1(VCC_net), .CO(n28810));
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n28808), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n29534), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_3 (.CI(n28808), .I0(n1057), .I1(VCC_net), .CO(n28809));
    SB_LUT4 rem_4_add_715_2_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(VCC_net), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_19 (.CI(n29534), .I0(n2342), .I1(VCC_net), 
            .CO(n29535));
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n29533), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1058), .I1(GND_net), 
            .CO(n28808));
    SB_CARRY rem_4_add_1586_18 (.CI(n29533), .I0(n2343), .I1(VCC_net), 
            .CO(n29534));
    SB_LUT4 i34718_4_lut (.I0(n37_adj_4744), .I1(n35_adj_4743), .I2(n33_adj_4742), 
            .I3(n42752), .O(n41571));
    defparam i34718_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n29532), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_17 (.CI(n29532), .I0(n2344), .I1(VCC_net), 
            .CO(n29533));
    SB_LUT4 div_46_LessThan_1545_i14_4_lut (.I0(n527), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4728));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n29531), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n29531), .I0(n2345), .I1(VCC_net), 
            .CO(n29532));
    SB_LUT4 i36294_3_lut (.I0(n14_adj_4728), .I1(n87), .I2(n37_adj_4744), 
            .I3(GND_net), .O(n43148));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36294_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_849_10_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n28800), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n28799), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_9 (.CI(n28799), .I0(n1251), .I1(VCC_net), .CO(n28800));
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n29530), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36295_3_lut (.I0(n43148), .I1(n86), .I2(n39_adj_4745), .I3(GND_net), 
            .O(n43149));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36295_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1586_15 (.CI(n29530), .I0(n2346), .I1(VCC_net), 
            .CO(n29531));
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n28798), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n29529), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_14 (.CI(n29529), .I0(n2347), .I1(VCC_net), 
            .CO(n29530));
    SB_LUT4 div_46_LessThan_1545_i40_3_lut (.I0(n22_adj_4735), .I1(n83), 
            .I2(n45_adj_4749), .I3(GND_net), .O(n40_adj_4746));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_849_8 (.CI(n28798), .I0(n1252), .I1(VCC_net), .CO(n28799));
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n28797), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_7 (.CI(n28797), .I0(n1253), .I1(VCC_net), .CO(n28798));
    SB_LUT4 i34692_4_lut (.I0(n43_adj_4748), .I1(n41_adj_4747), .I2(n39_adj_4745), 
            .I3(n41561), .O(n41545));
    defparam i34692_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n29528), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n28796), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35882_4_lut (.I0(n40_adj_4746), .I1(n20_adj_4733), .I2(n45_adj_4749), 
            .I3(n41542), .O(n42736));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35882_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_849_6 (.CI(n28796), .I0(n1254), .I1(GND_net), .CO(n28797));
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n28795), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36152_3_lut (.I0(n43149), .I1(n85), .I2(n41_adj_4747), .I3(GND_net), 
            .O(n43006));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36152_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1586_13 (.CI(n29528), .I0(n2348), .I1(VCC_net), 
            .CO(n29529));
    SB_CARRY rem_4_add_849_5 (.CI(n28795), .I0(n1255), .I1(GND_net), .CO(n28796));
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n29527), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n28794), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_4 (.CI(n28794), .I0(n1256), .I1(VCC_net), .CO(n28795));
    SB_LUT4 i13394_3_lut (.I0(setpoint[2]), .I1(n4380), .I2(n38059), .I3(GND_net), 
            .O(n18139));   // verilog/coms.v(126[12] 289[6])
    defparam i13394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n28793), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_12 (.CI(n29527), .I0(n2349), .I1(VCC_net), 
            .CO(n29528));
    SB_CARRY rem_4_add_849_3 (.CI(n28793), .I0(n1257), .I1(VCC_net), .CO(n28794));
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n29526), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_2_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(VCC_net), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i26_3_lut (.I0(n18_adj_4731), .I1(n91), 
            .I2(n29_adj_4740), .I3(GND_net), .O(n26_adj_4738));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1258), .I1(GND_net), 
            .CO(n28793));
    SB_CARRY rem_4_add_1586_11 (.CI(n29526), .I0(n2350), .I1(VCC_net), 
            .CO(n29527));
    SB_LUT4 i36466_4_lut (.I0(n26_adj_4738), .I1(n16_adj_4729), .I2(n29_adj_4740), 
            .I3(n41591), .O(n43320));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36466_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_782_4 (.CI(n28535), .I0(n1156), .I1(VCC_net), .CO(n28536));
    SB_LUT4 i36467_3_lut (.I0(n43320), .I1(n90), .I2(n31_adj_4741), .I3(GND_net), 
            .O(n43321));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36467_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13393_3_lut (.I0(setpoint[1]), .I1(n4379), .I2(n38059), .I3(GND_net), 
            .O(n18138));   // verilog/coms.v(126[12] 289[6])
    defparam i13393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n29525), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36320_3_lut (.I0(n43321), .I1(n89), .I2(n33_adj_4742), .I3(GND_net), 
            .O(n43174));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36320_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36118_4_lut (.I0(n43_adj_4748), .I1(n41_adj_4747), .I2(n39_adj_4745), 
            .I3(n41571), .O(n42972));
    defparam i36118_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1586_10 (.CI(n29525), .I0(n2351), .I1(VCC_net), 
            .CO(n29526));
    SB_LUT4 i13396_3_lut (.I0(setpoint[4]), .I1(n4382), .I2(n38059), .I3(GND_net), 
            .O(n18141));   // verilog/coms.v(126[12] 289[6])
    defparam i13396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n29524), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36367_4_lut (.I0(n43006), .I1(n42736), .I2(n45_adj_4749), 
            .I3(n41545), .O(n43221));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36367_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY rem_4_add_1586_9 (.CI(n29524), .I0(n2352), .I1(VCC_net), 
            .CO(n29525));
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n29523), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35444_3_lut (.I0(n43174), .I1(n88), .I2(n35_adj_4743), .I3(GND_net), 
            .O(n42298));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35444_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1586_8 (.CI(n29523), .I0(n2353), .I1(VCC_net), 
            .CO(n29524));
    SB_LUT4 i36369_4_lut (.I0(n42298), .I1(n43221), .I2(n45_adj_4749), 
            .I3(n42972), .O(n43223));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36369_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n43223), .I1(n15992), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n28534), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n29522), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_7 (.CI(n29522), .I0(n2354), .I1(GND_net), 
            .CO(n29523));
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n29521), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1721 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4983));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i7_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_782_3 (.CI(n28534), .I0(n1157), .I1(VCC_net), .CO(n28535));
    SB_CARRY rem_4_add_1586_6 (.CI(n29521), .I0(n2355), .I1(GND_net), 
            .CO(n29522));
    SB_LUT4 div_46_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4724));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_229[23]), 
            .I2(n3_adj_4351), .I3(n28775), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_229[22]), 
            .I2(n3_adj_4351), .I3(n28774), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n28774), .I0(displacement_23__N_229[22]), 
            .I1(n3_adj_4351), .CO(n28775));
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n29520), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_229[21]), 
            .I2(n3_adj_4351), .I3(n28773), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_5 (.CI(n29520), .I0(n2356), .I1(VCC_net), 
            .CO(n29521));
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n28773), .I0(displacement_23__N_229[21]), 
            .I1(n3_adj_4351), .CO(n28774));
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4579), .I2(VCC_net), 
            .I3(n29519), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_229[20]), 
            .I2(n3_adj_4351), .I3(n28772), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n28772), .I0(displacement_23__N_229[20]), 
            .I1(n3_adj_4351), .CO(n28773));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_229[19]), 
            .I2(n6_adj_4347), .I3(n28771), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n28771), .I0(displacement_23__N_229[19]), 
            .I1(n6_adj_4347), .CO(n28772));
    SB_LUT4 div_46_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4727));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_229[18]), 
            .I2(n7), .I3(n28770), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n28770), .I0(displacement_23__N_229[18]), 
            .I1(n7), .CO(n28771));
    SB_CARRY rem_4_add_1586_4 (.CI(n29519), .I0(n2357_adj_4579), .I1(VCC_net), 
            .CO(n29520));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_229[17]), 
            .I2(n8_adj_4373), .I3(n28769), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n28769), .I0(displacement_23__N_229[17]), 
            .I1(n8_adj_4373), .CO(n28770));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_229[16]), 
            .I2(n9_adj_4374), .I3(n28768), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4578), .I2(GND_net), 
            .I3(n29518), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_3 (.CI(n29518), .I0(n2358_adj_4578), .I1(GND_net), 
            .CO(n29519));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4516), .I1(VCC_net), 
            .CO(n29518));
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n28768), .I0(displacement_23__N_229[16]), 
            .I1(n9_adj_4374), .CO(n28769));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_229[15]), 
            .I2(n10_adj_4375), .I3(n28767), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4726));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n28767), .I0(displacement_23__N_229[15]), 
            .I1(n10_adj_4375), .CO(n28768));
    SB_LUT4 i13395_3_lut (.I0(setpoint[3]), .I1(n4381), .I2(n38059), .I3(GND_net), 
            .O(n18140));   // verilog/coms.v(126[12] 289[6])
    defparam i13395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1653_23_lut (.I0(n2471_adj_4515), .I1(n2438), .I2(VCC_net), 
            .I3(n29517), .O(n2537_adj_4514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_229[14]), 
            .I2(n11_adj_4376), .I3(n28766), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_30_lut (.I0(n3164), .I1(n3131), .I2(VCC_net), 
            .I3(n29280), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n28766), .I0(displacement_23__N_229[14]), 
            .I1(n11_adj_4376), .CO(n28767));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_229[13]), 
            .I2(n12_adj_4377), .I3(n28765), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13327_3_lut (.I0(encoder0_position[23]), .I1(n2999), .I2(count_enable), 
            .I3(GND_net), .O(n18072));   // quad.v(35[10] 41[6])
    defparam i13327_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n28765), .I0(displacement_23__N_229[13]), 
            .I1(n12_adj_4377), .CO(n28766));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_229[12]), 
            .I2(n13_adj_4378), .I3(n28764), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n28764), .I0(displacement_23__N_229[12]), 
            .I1(n13_adj_4378), .CO(n28765));
    SB_LUT4 div_46_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4725));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n29279), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(GND_net), .I1(n2439), .I2(VCC_net), 
            .I3(n29516), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_229[11]), 
            .I2(n14_adj_4379), .I3(n28763), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n28763), .I0(displacement_23__N_229[11]), 
            .I1(n14_adj_4379), .CO(n28764));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_229[10]), 
            .I2(n15_adj_4380), .I3(n28762), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n28762), .I0(displacement_23__N_229[10]), 
            .I1(n15_adj_4380), .CO(n28763));
    SB_CARRY rem_4_add_1653_22 (.CI(n29516), .I0(n2439), .I1(VCC_net), 
            .CO(n29517));
    SB_LUT4 div_46_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n526));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_229[9]), 
            .I2(n16_adj_4381), .I3(n28761), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n28761), .I0(displacement_23__N_229[9]), 
            .I1(n16_adj_4381), .CO(n28762));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_229[8]), 
            .I2(n17_adj_4382), .I3(n28760), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13326_3_lut (.I0(encoder0_position[22]), .I1(n3000), .I2(count_enable), 
            .I3(GND_net), .O(n18071));   // quad.v(35[10] 41[6])
    defparam i13326_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n28760), .I0(displacement_23__N_229[8]), 
            .I1(n17_adj_4382), .CO(n28761));
    SB_LUT4 i13325_3_lut (.I0(encoder0_position[21]), .I1(n3001), .I2(count_enable), 
            .I3(GND_net), .O(n18070));   // quad.v(35[10] 41[6])
    defparam i13325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_229[7]), 
            .I2(n18_adj_4383), .I3(n28759), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_29 (.CI(n29279), .I0(n3132), .I1(VCC_net), 
            .CO(n29280));
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n28759), .I0(displacement_23__N_229[7]), 
            .I1(n18_adj_4383), .CO(n28760));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_229[6]), 
            .I2(n19_adj_4384), .I3(n28758), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_21_lut (.I0(GND_net), .I1(n2440), .I2(VCC_net), 
            .I3(n29515), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n29278), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_21 (.CI(n29515), .I0(n2440), .I1(VCC_net), 
            .CO(n29516));
    SB_LUT4 rem_4_add_1653_20_lut (.I0(GND_net), .I1(n2441), .I2(VCC_net), 
            .I3(n29514), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_28 (.CI(n29278), .I0(n3133), .I1(VCC_net), 
            .CO(n29279));
    SB_CARRY rem_4_add_1653_20 (.CI(n29514), .I0(n2441), .I1(VCC_net), 
            .CO(n29515));
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n29277), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n28758), .I0(displacement_23__N_229[6]), 
            .I1(n19_adj_4384), .CO(n28759));
    SB_LUT4 rem_4_add_1653_19_lut (.I0(GND_net), .I1(n2442), .I2(VCC_net), 
            .I3(n29513), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_27 (.CI(n29277), .I0(n3134), .I1(VCC_net), 
            .CO(n29278));
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n29276), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_229[5]), 
            .I2(n20_adj_4385), .I3(n28757), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n28757), .I0(displacement_23__N_229[5]), 
            .I1(n20_adj_4385), .CO(n28758));
    SB_CARRY rem_4_add_1653_19 (.CI(n29513), .I0(n2442), .I1(VCC_net), 
            .CO(n29514));
    SB_CARRY rem_4_add_2122_26 (.CI(n29276), .I0(n3135), .I1(VCC_net), 
            .CO(n29277));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_229[4]), 
            .I2(n21_adj_4386), .I3(n28756), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n28756), .I0(displacement_23__N_229[4]), 
            .I1(n21_adj_4386), .CO(n28757));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_229[3]), 
            .I2(n22_adj_4387), .I3(n28755), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_18_lut (.I0(GND_net), .I1(n2443), .I2(VCC_net), 
            .I3(n29512), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n28755), .I0(displacement_23__N_229[3]), 
            .I1(n22_adj_4387), .CO(n28756));
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n29275), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_2_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(VCC_net), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_229[2]), 
            .I2(n23_adj_4388), .I3(n28754), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n28754), .I0(displacement_23__N_229[2]), 
            .I1(n23_adj_4388), .CO(n28755));
    SB_LUT4 div_46_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4721));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_229[1]), 
            .I2(n24_adj_4389), .I3(n28753), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n28753), .I0(displacement_23__N_229[1]), 
            .I1(n24_adj_4389), .CO(n28754));
    SB_CARRY rem_4_add_1653_18 (.CI(n29512), .I0(n2443), .I1(VCC_net), 
            .CO(n29513));
    SB_CARRY rem_4_add_2122_25 (.CI(n29275), .I0(n3136), .I1(VCC_net), 
            .CO(n29276));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_229[0]), 
            .I2(n25_adj_4390), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_17_lut (.I0(GND_net), .I1(n2444), .I2(VCC_net), 
            .I3(n29511), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n29274), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4722));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4723));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_229[0]), 
            .I1(n25_adj_4390), .CO(n28753));
    SB_CARRY rem_4_add_1653_17 (.CI(n29511), .I0(n2444), .I1(VCC_net), 
            .CO(n29512));
    SB_LUT4 rem_4_add_1653_16_lut (.I0(GND_net), .I1(n2445), .I2(VCC_net), 
            .I3(n29510), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_24 (.CI(n29274), .I0(n3137), .I1(VCC_net), 
            .CO(n29275));
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1158), .I1(GND_net), 
            .CO(n28534));
    SB_CARRY rem_4_add_1653_16 (.CI(n29510), .I0(n2445), .I1(VCC_net), 
            .CO(n29511));
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n29273), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_15_lut (.I0(GND_net), .I1(n2446), .I2(VCC_net), 
            .I3(n29509), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_23 (.CI(n29273), .I0(n3138), .I1(VCC_net), 
            .CO(n29274));
    SB_CARRY rem_4_add_1653_15 (.CI(n29509), .I0(n2446), .I1(VCC_net), 
            .CO(n29510));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(GND_net), .I1(n2447_adj_4575), .I2(VCC_net), 
            .I3(n29508), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n29272), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_22 (.CI(n29272), .I0(n3139), .I1(VCC_net), 
            .CO(n29273));
    SB_CARRY rem_4_add_1653_14 (.CI(n29508), .I0(n2447_adj_4575), .I1(VCC_net), 
            .CO(n29509));
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n29271), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_21 (.CI(n29271), .I0(n3140), .I1(VCC_net), 
            .CO(n29272));
    SB_LUT4 rem_4_add_1653_13_lut (.I0(GND_net), .I1(n2448_adj_4574), .I2(VCC_net), 
            .I3(n29507), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n29270), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4718));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1653_13 (.CI(n29507), .I0(n2448_adj_4574), .I1(VCC_net), 
            .CO(n29508));
    SB_LUT4 rem_4_add_1653_12_lut (.I0(GND_net), .I1(n2449_adj_4573), .I2(VCC_net), 
            .I3(n29506), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_12 (.CI(n29506), .I0(n2449_adj_4573), .I1(VCC_net), 
            .CO(n29507));
    SB_CARRY rem_4_add_2122_20 (.CI(n29270), .I0(n3141), .I1(VCC_net), 
            .CO(n29271));
    SB_LUT4 rem_4_add_1653_11_lut (.I0(GND_net), .I1(n2450_adj_4572), .I2(VCC_net), 
            .I3(n29505), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n29269), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_11 (.CI(n29505), .I0(n2450_adj_4572), .I1(VCC_net), 
            .CO(n29506));
    SB_CARRY rem_4_add_2122_19 (.CI(n29269), .I0(n3142), .I1(VCC_net), 
            .CO(n29270));
    SB_LUT4 rem_4_add_1653_10_lut (.I0(GND_net), .I1(n2451_adj_4571), .I2(VCC_net), 
            .I3(n29504), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n29268), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_10 (.CI(n29504), .I0(n2451_adj_4571), .I1(VCC_net), 
            .CO(n29505));
    SB_CARRY rem_4_add_2122_18 (.CI(n29268), .I0(n3143), .I1(VCC_net), 
            .CO(n29269));
    SB_LUT4 rem_4_add_1653_9_lut (.I0(GND_net), .I1(n2452_adj_4570), .I2(VCC_net), 
            .I3(n29503), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n29267), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4720));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2122_17 (.CI(n29267), .I0(n3144), .I1(VCC_net), 
            .CO(n29268));
    SB_CARRY rem_4_add_1653_9 (.CI(n29503), .I0(n2452_adj_4570), .I1(VCC_net), 
            .CO(n29504));
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n29266), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n29266), .I0(n3145), .I1(VCC_net), 
            .CO(n29267));
    SB_LUT4 rem_4_add_1653_8_lut (.I0(GND_net), .I1(n2453_adj_4569), .I2(VCC_net), 
            .I3(n29502), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n29265), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_8 (.CI(n29502), .I0(n2453_adj_4569), .I1(VCC_net), 
            .CO(n29503));
    SB_CARRY rem_4_add_2122_15 (.CI(n29265), .I0(n3146), .I1(VCC_net), 
            .CO(n29266));
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n29264), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_7_lut (.I0(GND_net), .I1(n2454_adj_4568), .I2(GND_net), 
            .I3(n29501), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_14 (.CI(n29264), .I0(n3147), .I1(VCC_net), 
            .CO(n29265));
    SB_DFF blink_53 (.Q(blink), .C(LED_c), .D(blink_N_255));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    SB_CARRY rem_4_add_1653_7 (.CI(n29501), .I0(n2454_adj_4568), .I1(GND_net), 
            .CO(n29502));
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n29263), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4712));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1653_6_lut (.I0(GND_net), .I1(n2455_adj_4567), .I2(GND_net), 
            .I3(n29500), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_13 (.CI(n29263), .I0(n3148), .I1(VCC_net), 
            .CO(n29264));
    SB_CARRY rem_4_add_1653_6 (.CI(n29500), .I0(n2455_adj_4567), .I1(GND_net), 
            .CO(n29501));
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n29262), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_5_lut (.I0(GND_net), .I1(n2456_adj_4518), .I2(VCC_net), 
            .I3(n29499), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_12 (.CI(n29262), .I0(n3149), .I1(VCC_net), 
            .CO(n29263));
    SB_LUT4 div_46_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4714));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13324_3_lut (.I0(encoder0_position[20]), .I1(n3002), .I2(count_enable), 
            .I3(GND_net), .O(n18069));   // quad.v(35[10] 41[6])
    defparam i13324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13323_3_lut (.I0(encoder0_position[19]), .I1(n3003), .I2(count_enable), 
            .I3(GND_net), .O(n18068));   // quad.v(35[10] 41[6])
    defparam i13323_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_5 (.CI(n29499), .I0(n2456_adj_4518), .I1(VCC_net), 
            .CO(n29500));
    SB_LUT4 rem_4_add_1653_4_lut (.I0(GND_net), .I1(n2457_adj_4517), .I2(VCC_net), 
            .I3(n29498), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n29261), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_4 (.CI(n29498), .I0(n2457_adj_4517), .I1(VCC_net), 
            .CO(n29499));
    SB_CARRY rem_4_add_2122_11 (.CI(n29261), .I0(n3150), .I1(VCC_net), 
            .CO(n29262));
    SB_LUT4 rem_4_add_1653_3_lut (.I0(GND_net), .I1(n2458_adj_4516), .I2(GND_net), 
            .I3(n29497), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n29260), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4716));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1653_3 (.CI(n29497), .I0(n2458_adj_4516), .I1(GND_net), 
            .CO(n29498));
    SB_CARRY rem_4_add_2122_10 (.CI(n29260), .I0(n3151), .I1(VCC_net), 
            .CO(n29261));
    SB_LUT4 div_46_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4717));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4497), .I1(VCC_net), 
            .CO(n29497));
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n29259), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4514), .I2(VCC_net), 
            .I3(n29496), .O(n2636_adj_4480)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2122_9 (.CI(n29259), .I0(n3152), .I1(VCC_net), 
            .CO(n29260));
    SB_LUT4 rem_4_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4513), .I2(VCC_net), 
            .I3(n29495), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n29258), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4710));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13322_3_lut (.I0(encoder0_position[18]), .I1(n3004), .I2(count_enable), 
            .I3(GND_net), .O(n18067));   // quad.v(35[10] 41[6])
    defparam i13322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34840_4_lut (.I0(n23_adj_4716), .I1(n21_adj_4714), .I2(n19_adj_4712), 
            .I3(n17_adj_4710), .O(n41694));
    defparam i34840_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1720_23 (.CI(n29495), .I0(n2538_adj_4513), .I1(VCC_net), 
            .CO(n29496));
    SB_CARRY rem_4_add_2122_8 (.CI(n29258), .I0(n3153), .I1(VCC_net), 
            .CO(n29259));
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4512), .I2(VCC_net), 
            .I3(n29494), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_22 (.CI(n29494), .I0(n2539_adj_4512), .I1(VCC_net), 
            .CO(n29495));
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541_adj_4510), .I1(n2608), .I2(n2570), 
            .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n29257), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_7 (.CI(n29257), .I0(n3154), .I1(GND_net), 
            .CO(n29258));
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4511), .I2(VCC_net), 
            .I3(n29493), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34801_4_lut (.I0(n29_adj_4720), .I1(n27_adj_4718), .I2(n25_adj_4717), 
            .I3(n41694), .O(n41654));
    defparam i34801_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n29256), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13336_3_lut (.I0(encoder1_position[7]), .I1(n2965), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18081));   // quad.v(35[10] 41[6])
    defparam i13336_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_21 (.CI(n29493), .I0(n2540_adj_4511), .I1(VCC_net), 
            .CO(n29494));
    SB_CARRY rem_4_add_2122_6 (.CI(n29256), .I0(n3155), .I1(GND_net), 
            .CO(n29257));
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4510), .I2(VCC_net), 
            .I3(n29492), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n29255), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_20 (.CI(n29492), .I0(n2541_adj_4510), .I1(VCC_net), 
            .CO(n29493));
    SB_CARRY rem_4_add_2122_5 (.CI(n29255), .I0(n3156), .I1(VCC_net), 
            .CO(n29256));
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4509), .I2(VCC_net), 
            .I3(n29491), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_19 (.CI(n29491), .I0(n2542_adj_4509), .I1(VCC_net), 
            .CO(n29492));
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n29254), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_4 (.CI(n29254), .I0(n3157), .I1(VCC_net), 
            .CO(n29255));
    SB_LUT4 i36213_4_lut (.I0(n35_adj_4723), .I1(n33_adj_4722), .I2(n31_adj_4721), 
            .I3(n41654), .O(n43067));
    defparam i36213_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4508), .I2(VCC_net), 
            .I3(n29490), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(n29253), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_18 (.CI(n29490), .I0(n2543_adj_4508), .I1(VCC_net), 
            .CO(n29491));
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4507), .I2(VCC_net), 
            .I3(n29489), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_3 (.CI(n29253), .I0(n3158), .I1(GND_net), 
            .CO(n29254));
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3258), .I1(VCC_net), 
            .CO(n29253));
    SB_CARRY rem_4_add_1720_17 (.CI(n29489), .I0(n2544_adj_4507), .I1(VCC_net), 
            .CO(n29490));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4506), .I2(VCC_net), 
            .I3(n29488), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i16_4_lut (.I0(n526), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4709));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_1720_16 (.CI(n29488), .I0(n2545_adj_4506), .I1(VCC_net), 
            .CO(n29489));
    SB_LUT4 i36088_3_lut (.I0(n16_adj_4709), .I1(n87), .I2(n39_adj_4725), 
            .I3(GND_net), .O(n42942));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36088_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4505), .I2(VCC_net), 
            .I3(n29487), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_15 (.CI(n29487), .I0(n2546_adj_4505), .I1(VCC_net), 
            .CO(n29488));
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4504), .I2(VCC_net), 
            .I3(n29486), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_14 (.CI(n29486), .I0(n2547_adj_4504), .I1(VCC_net), 
            .CO(n29487));
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539_adj_4512), .I1(n2606), .I2(n2570), 
            .I3(GND_net), .O(n2638_adj_4478));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4503), .I2(VCC_net), 
            .I3(n29485), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36089_3_lut (.I0(n42942), .I1(n86), .I2(n41_adj_4726), .I3(GND_net), 
            .O(n42943));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36089_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1720_13 (.CI(n29485), .I0(n2548_adj_4503), .I1(VCC_net), 
            .CO(n29486));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4502), .I2(VCC_net), 
            .I3(n29484), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_12 (.CI(n29484), .I0(n2549_adj_4502), .I1(VCC_net), 
            .CO(n29485));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4501), .I2(VCC_net), 
            .I3(n29483), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_11 (.CI(n29483), .I0(n2550_adj_4501), .I1(VCC_net), 
            .CO(n29484));
    GND i1 (.Y(GND_net));
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4500), .I2(VCC_net), 
            .I3(n29482), .O(n2618_adj_4491)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut_adj_1722 (.I0(n2638_adj_4478), .I1(n2640), .I2(n2639), 
            .I3(n2641), .O(n30_adj_4897));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1720_10 (.CI(n29482), .I0(n2551_adj_4500), .I1(VCC_net), 
            .CO(n29483));
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4499), .I2(VCC_net), 
            .I3(n29481), .O(n2619_adj_4492)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13335_3_lut (.I0(encoder1_position[6]), .I1(n2966), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18080));   // quad.v(35[10] 41[6])
    defparam i13335_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_9 (.CI(n29481), .I0(n2552_adj_4499), .I1(VCC_net), 
            .CO(n29482));
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4498), .I2(VCC_net), 
            .I3(n29480), .O(n2620_adj_4486)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35521_4_lut (.I0(n41_adj_4726), .I1(n39_adj_4725), .I2(n27_adj_4718), 
            .I3(n41690), .O(n42375));
    defparam i35521_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY rem_4_add_1720_8 (.CI(n29480), .I0(n2553_adj_4498), .I1(VCC_net), 
            .CO(n29481));
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n29479), .O(n2621_adj_4485)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36149_3_lut (.I0(n22_adj_4715), .I1(n93), .I2(n27_adj_4718), 
            .I3(GND_net), .O(n43003));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36149_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35434_3_lut (.I0(n42943), .I1(n85), .I2(n43_adj_4727), .I3(GND_net), 
            .O(n42288));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35434_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1482_i28_3_lut (.I0(n20_adj_4713), .I1(n91), 
            .I2(n31_adj_4721), .I3(GND_net), .O(n28_adj_4719));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36462_4_lut (.I0(n28_adj_4719), .I1(n18_adj_4711), .I2(n31_adj_4721), 
            .I3(n41650), .O(n43316));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36462_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36463_3_lut (.I0(n43316), .I1(n90), .I2(n33_adj_4722), .I3(GND_net), 
            .O(n43317));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36463_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36336_3_lut (.I0(n43317), .I1(n89), .I2(n35_adj_4723), .I3(GND_net), 
            .O(n43190));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36336_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35523_4_lut (.I0(n41_adj_4726), .I1(n39_adj_4725), .I2(n37_adj_4724), 
            .I3(n43067), .O(n42377));
    defparam i35523_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36333_4_lut (.I0(n42288), .I1(n43003), .I2(n43_adj_4727), 
            .I3(n42375), .O(n43187));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36333_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35432_3_lut (.I0(n43190), .I1(n88), .I2(n37_adj_4724), .I3(GND_net), 
            .O(n42286));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35432_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36549_4_lut (.I0(n42286), .I1(n43187), .I2(n43_adj_4727), 
            .I3(n42377), .O(n43403));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36549_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36550_3_lut (.I0(n43403), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n43404));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36550_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n43404), .I1(n16007), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4705));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4708));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4707));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4702));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4703));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4704));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4706));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n525));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4692));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4694));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4696));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4698));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4699));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4701));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4690));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13334_3_lut (.I0(encoder1_position[5]), .I1(n2967), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18079));   // quad.v(35[10] 41[6])
    defparam i13334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13333_3_lut (.I0(encoder1_position[4]), .I1(n2968), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18078));   // quad.v(35[10] 41[6])
    defparam i13333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34952_4_lut (.I0(n25_adj_4696), .I1(n23_adj_4694), .I2(n21_adj_4692), 
            .I3(n19_adj_4690), .O(n41806));
    defparam i34952_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34944_4_lut (.I0(n31_adj_4701), .I1(n29_adj_4699), .I2(n27_adj_4698), 
            .I3(n41806), .O(n41798));
    defparam i34944_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36227_4_lut (.I0(n37_adj_4704), .I1(n35_adj_4703), .I2(n33_adj_4702), 
            .I3(n41798), .O(n43081));
    defparam i36227_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1417_i18_4_lut (.I0(n525), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4689));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i13332_3_lut (.I0(encoder1_position[3]), .I1(n2969), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18077));   // quad.v(35[10] 41[6])
    defparam i13332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13331_3_lut (.I0(encoder1_position[2]), .I1(n2970), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18076));   // quad.v(35[10] 41[6])
    defparam i13331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36096_3_lut (.I0(n18_adj_4689), .I1(n87), .I2(n41_adj_4706), 
            .I3(GND_net), .O(n42950));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36096_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36097_3_lut (.I0(n42950), .I1(n86), .I2(n43_adj_4707), .I3(GND_net), 
            .O(n42951));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36097_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13330_3_lut (.I0(encoder1_position[1]), .I1(n2971), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n18075));   // quad.v(35[10] 41[6])
    defparam i13330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35557_4_lut (.I0(n43_adj_4707), .I1(n41_adj_4706), .I2(n29_adj_4699), 
            .I3(n41804), .O(n42411));
    defparam i35557_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1417_i26_3_lut (.I0(n24_adj_4695), .I1(n93), 
            .I2(n29_adj_4699), .I3(GND_net), .O(n26_adj_4697));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35426_3_lut (.I0(n42951), .I1(n85), .I2(n45_adj_4708), .I3(GND_net), 
            .O(n42280));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35426_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1417_i30_3_lut (.I0(n22_adj_4693), .I1(n91), 
            .I2(n33_adj_4702), .I3(GND_net), .O(n30_adj_4700));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36460_4_lut (.I0(n30_adj_4700), .I1(n20_adj_4691), .I2(n33_adj_4702), 
            .I3(n41796), .O(n43314));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36460_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36461_3_lut (.I0(n43314), .I1(n90), .I2(n35_adj_4703), .I3(GND_net), 
            .O(n43315));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36461_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36338_3_lut (.I0(n43315), .I1(n89), .I2(n37_adj_4704), .I3(GND_net), 
            .O(n43192));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36338_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35561_4_lut (.I0(n43_adj_4707), .I1(n41_adj_4706), .I2(n39_adj_4705), 
            .I3(n43081), .O(n42415));
    defparam i35561_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36144_4_lut (.I0(n42280), .I1(n26_adj_4697), .I2(n45_adj_4708), 
            .I3(n42411), .O(n42998));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36144_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35424_3_lut (.I0(n43192), .I1(n88), .I2(n39_adj_4705), .I3(GND_net), 
            .O(n42278));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35424_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36146_4_lut (.I0(n42278), .I1(n42998), .I2(n45_adj_4708), 
            .I3(n42415), .O(n43000));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36146_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n43000), .I1(n16011), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4688));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4687));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4686));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4685));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4675));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4677));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13407_3_lut (.I0(setpoint[15]), .I1(n4393), .I2(n38059), 
            .I3(GND_net), .O(n18152));   // verilog/coms.v(126[12] 289[6])
    defparam i13407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4679));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4681));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4682));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4684));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4673));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34998_4_lut (.I0(n27_adj_4679), .I1(n25_adj_4677), .I2(n23_adj_4675), 
            .I3(n21_adj_4673), .O(n41852));
    defparam i34998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34992_4_lut (.I0(n33_adj_4684), .I1(n31_adj_4682), .I2(n29_adj_4681), 
            .I3(n41852), .O(n41846));
    defparam i34992_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1350_i20_4_lut (.I0(n524), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4672));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1350_i28_3_lut (.I0(n26_adj_4678), .I1(n93), 
            .I2(n31_adj_4682), .I3(GND_net), .O(n28_adj_4680));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1350_i32_3_lut (.I0(n24_adj_4676), .I1(n91), 
            .I2(n35_adj_4685), .I3(GND_net), .O(n32_adj_4683));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36456_4_lut (.I0(n32_adj_4683), .I1(n22_adj_4674), .I2(n35_adj_4685), 
            .I3(n41842), .O(n43310));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36456_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36457_3_lut (.I0(n43310), .I1(n90), .I2(n37_adj_4686), .I3(GND_net), 
            .O(n43311));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36457_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36344_3_lut (.I0(n43311), .I1(n89), .I2(n39_adj_4687), .I3(GND_net), 
            .O(n43198));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36344_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13406_3_lut (.I0(setpoint[14]), .I1(n4392), .I2(n38059), 
            .I3(GND_net), .O(n18151));   // verilog/coms.v(126[12] 289[6])
    defparam i13406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36235_4_lut (.I0(n39_adj_4687), .I1(n37_adj_4686), .I2(n35_adj_4685), 
            .I3(n41846), .O(n43089));
    defparam i36235_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36458_4_lut (.I0(n28_adj_4680), .I1(n20_adj_4672), .I2(n31_adj_4682), 
            .I3(n41850), .O(n43312));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36458_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35412_3_lut (.I0(n43198), .I1(n88), .I2(n41_adj_4688), .I3(GND_net), 
            .O(n42266));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35412_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36512_4_lut (.I0(n42266), .I1(n43312), .I2(n41_adj_4688), 
            .I3(n43089), .O(n43366));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36512_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36513_3_lut (.I0(n43366), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n43367));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36513_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36496_3_lut (.I0(n43367), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n43350));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36496_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n43350), .I1(n16004), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4670));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4669));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4671));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4668));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4664));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4665));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4667));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13405_3_lut (.I0(setpoint[13]), .I1(n4391), .I2(n38059), 
            .I3(GND_net), .O(n18150));   // verilog/coms.v(126[12] 289[6])
    defparam i13405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4658));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4660));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4662));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13404_3_lut (.I0(setpoint[12]), .I1(n4390), .I2(n38059), 
            .I3(GND_net), .O(n18149));   // verilog/coms.v(126[12] 289[6])
    defparam i13404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4656));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35053_4_lut (.I0(n29_adj_4662), .I1(n27_adj_4660), .I2(n25_adj_4658), 
            .I3(n23_adj_4656), .O(n41907));
    defparam i35053_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35043_4_lut (.I0(n35_adj_4667), .I1(n33_adj_4665), .I2(n31_adj_4664), 
            .I3(n41907), .O(n41897));
    defparam i35043_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1281_i22_4_lut (.I0(n523), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4655));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1281_i30_3_lut (.I0(n28_adj_4661), .I1(n93), 
            .I2(n33_adj_4665), .I3(GND_net), .O(n30_adj_4663));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1281_i34_3_lut (.I0(n26_adj_4659), .I1(n91), 
            .I2(n37_adj_4668), .I3(GND_net), .O(n34_adj_4666));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36454_4_lut (.I0(n34_adj_4666), .I1(n24_adj_4657), .I2(n37_adj_4668), 
            .I3(n41891), .O(n43308));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36454_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36455_3_lut (.I0(n43308), .I1(n90), .I2(n39_adj_4669), .I3(GND_net), 
            .O(n43309));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36455_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36346_3_lut (.I0(n43309), .I1(n89), .I2(n41_adj_4670), .I3(GND_net), 
            .O(n43200));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36346_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36243_4_lut (.I0(n41_adj_4670), .I1(n39_adj_4669), .I2(n37_adj_4668), 
            .I3(n41897), .O(n43097));
    defparam i36243_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36444_4_lut (.I0(n30_adj_4663), .I1(n22_adj_4655), .I2(n33_adj_4665), 
            .I3(n41903), .O(n43298));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36444_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35408_3_lut (.I0(n43200), .I1(n88), .I2(n43_adj_4671), .I3(GND_net), 
            .O(n42262));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35408_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36535_4_lut (.I0(n42262), .I1(n43298), .I2(n43_adj_4671), 
            .I3(n43097), .O(n43389));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36535_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36536_3_lut (.I0(n43389), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n43390));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36536_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n43390), .I1(n15959), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4651));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4361), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4650));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4654));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4653));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13403_3_lut (.I0(setpoint[11]), .I1(n4389), .I2(n38059), 
            .I3(GND_net), .O(n18148));   // verilog/coms.v(126[12] 289[6])
    defparam i13403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4644));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4646));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4648));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4642));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35108_4_lut (.I0(n31_adj_4648), .I1(n29_adj_4646), .I2(n27_adj_4644), 
            .I3(n25_adj_4642), .O(n41962));
    defparam i35108_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1210_i36_3_lut (.I0(n28_adj_4645), .I1(n91), 
            .I2(n39_adj_4654), .I3(GND_net), .O(n36_adj_4652));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1210_i24_4_lut (.I0(n522), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4641));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1210_i32_3_lut (.I0(n30_adj_4647), .I1(n93), 
            .I2(n35_adj_4651), .I3(GND_net), .O(n32_adj_4649));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35091_4_lut (.I0(n37_adj_4653), .I1(n35_adj_4651), .I2(n33_adj_4650), 
            .I3(n41962), .O(n41945));
    defparam i35091_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36452_4_lut (.I0(n36_adj_4652), .I1(n26_adj_4643), .I2(n39_adj_4654), 
            .I3(n41937), .O(n43306));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36452_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36134_4_lut (.I0(n32_adj_4649), .I1(n24_adj_4641), .I2(n35_adj_4651), 
            .I3(n41956), .O(n42988));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36134_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36584_4_lut (.I0(n42988), .I1(n43306), .I2(n39_adj_4654), 
            .I3(n41945), .O(n43438));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36584_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36585_3_lut (.I0(n43438), .I1(n90), .I2(n1865), .I3(GND_net), 
            .O(n43439));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36585_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36538_3_lut (.I0(n43439), .I1(n89), .I2(n1864), .I3(GND_net), 
            .O(n43392));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36538_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36136_3_lut (.I0(n43392), .I1(n88), .I2(n1863), .I3(GND_net), 
            .O(n42990));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36136_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n42990), .I1(n15953), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'hceef;
    SB_LUT4 i13010_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13293), .I3(GND_net), .O(n17755));   // verilog/coms.v(126[12] 289[6])
    defparam i13010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13402_3_lut (.I0(setpoint[10]), .I1(n4388), .I2(n38059), 
            .I3(GND_net), .O(n18147));   // verilog/coms.v(126[12] 289[6])
    defparam i13402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13401_3_lut (.I0(setpoint[9]), .I1(n4387), .I2(n38059), .I3(GND_net), 
            .O(n18146));   // verilog/coms.v(126[12] 289[6])
    defparam i13401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4637));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4636));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4334), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4640));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4632));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4635));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4634));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4639));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4630));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35145_4_lut (.I0(n33_adj_4635), .I1(n31_adj_4634), .I2(n29_adj_4632), 
            .I3(n27_adj_4630), .O(n41999));
    defparam i35145_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1137_i38_3_lut (.I0(n30_adj_4633), .I1(n91), 
            .I2(n41_adj_4640), .I3(GND_net), .O(n38_adj_4638));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1137_i26_4_lut (.I0(n521), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_4629));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36138_3_lut (.I0(n26_adj_4629), .I1(n95), .I2(n33_adj_4635), 
            .I3(GND_net), .O(n42992));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36138_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36139_3_lut (.I0(n42992), .I1(n94), .I2(n35_adj_4636), .I3(GND_net), 
            .O(n42993));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36139_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35132_4_lut (.I0(n39_adj_4639), .I1(n37_adj_4637), .I2(n35_adj_4636), 
            .I3(n41999), .O(n41986));
    defparam i35132_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36448_4_lut (.I0(n38_adj_4638), .I1(n28_adj_4631), .I2(n41_adj_4640), 
            .I3(n41980), .O(n43302));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36448_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35392_3_lut (.I0(n42993), .I1(n93), .I2(n37_adj_4637), .I3(GND_net), 
            .O(n42246));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35392_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36576_4_lut (.I0(n42246), .I1(n43302), .I2(n41_adj_4640), 
            .I3(n41986), .O(n43430));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36576_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36577_3_lut (.I0(n43430), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n43431));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36577_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36556_3_lut (.I0(n43431), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n43410));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36556_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n43410), .I1(n15989), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hceef;
    SB_LUT4 i13400_3_lut (.I0(setpoint[8]), .I1(n4386), .I2(n38059), .I3(GND_net), 
            .O(n18145));   // verilog/coms.v(126[12] 289[6])
    defparam i13400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4623));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4624));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4344), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4627));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4626));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4619));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4621));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4622));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4617));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34476_4_lut (.I0(n35_adj_4622), .I1(n33_adj_4621), .I2(n31_adj_4619), 
            .I3(n29_adj_4617), .O(n41329));
    defparam i34476_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1062_i40_3_lut (.I0(n32_adj_4620), .I1(n91), 
            .I2(n43_adj_4627), .I3(GND_net), .O(n40_adj_4625));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1062_i28_4_lut (.I0(n520), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4616));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36301_3_lut (.I0(n28_adj_4616), .I1(n95), .I2(n35_adj_4622), 
            .I3(GND_net), .O(n43155));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36301_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36302_3_lut (.I0(n43155), .I1(n94), .I2(n37_adj_4623), .I3(GND_net), 
            .O(n43156));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36302_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13399_3_lut (.I0(setpoint[7]), .I1(n4385), .I2(n38059), .I3(GND_net), 
            .O(n18144));   // verilog/coms.v(126[12] 289[6])
    defparam i13399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34468_4_lut (.I0(n41_adj_4626), .I1(n39_adj_4624), .I2(n37_adj_4623), 
            .I3(n41329), .O(n41321));
    defparam i34468_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36446_4_lut (.I0(n40_adj_4625), .I1(n30_adj_4618), .I2(n43_adj_4627), 
            .I3(n42040), .O(n43300));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36446_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36129_3_lut (.I0(n43156), .I1(n93), .I2(n39_adj_4624), .I3(GND_net), 
            .O(n42983));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36129_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36553_4_lut (.I0(n42983), .I1(n43300), .I2(n43_adj_4627), 
            .I3(n41321), .O(n43407));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36553_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36554_3_lut (.I0(n43407), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n43408));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36554_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n43408), .I1(n15986), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4470), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4612));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13415_3_lut (.I0(setpoint[23]), .I1(n4401), .I2(n38059), 
            .I3(GND_net), .O(n18160));   // verilog/coms.v(126[12] 289[6])
    defparam i13415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4342), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4611));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4615));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13414_3_lut (.I0(setpoint[22]), .I1(n4400), .I2(n38059), 
            .I3(GND_net), .O(n18159));   // verilog/coms.v(126[12] 289[6])
    defparam i13414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4614));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut (.I0(bit_ctr[30]), .I1(n41273), .I2(n4472), .I3(GND_net), 
            .O(n34096));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1730 (.I0(bit_ctr[0]), .I1(n41272), .I2(n4472), 
            .I3(GND_net), .O(n34094));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1730.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4608));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4610));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1731 (.I0(n35274), .I1(r_Clock_Count[0]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n35004));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1731.LUT_INIT = 16'heaea;
    SB_LUT4 div_46_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4606));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34502_4_lut (.I0(n37_adj_4610), .I1(n35), .I2(n33_adj_4608), 
            .I3(n31_adj_4606), .O(n41355));
    defparam i34502_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_985_i42_3_lut (.I0(n34_adj_4609), .I1(n91), 
            .I2(n45_adj_4615), .I3(GND_net), .O(n42_adj_4613));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_985_i30_4_lut (.I0(n519), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4605));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36303_3_lut (.I0(n30_adj_4605), .I1(n95), .I2(n37_adj_4610), 
            .I3(GND_net), .O(n43157));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36303_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36304_3_lut (.I0(n43157), .I1(n94), .I2(n39_adj_4611), .I3(GND_net), 
            .O(n43158));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36304_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34492_4_lut (.I0(n43_adj_4614), .I1(n41_adj_4612), .I2(n39_adj_4611), 
            .I3(n41355), .O(n41345));
    defparam i34492_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35876_4_lut (.I0(n42_adj_4613), .I1(n32_adj_4607), .I2(n45_adj_4615), 
            .I3(n41339), .O(n42730));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35876_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36127_3_lut (.I0(n43158), .I1(n93), .I2(n41_adj_4612), .I3(GND_net), 
            .O(n42981));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36127_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36357_4_lut (.I0(n42981), .I1(n42730), .I2(n45_adj_4615), 
            .I3(n41345), .O(n43211));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36357_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n43211), .I1(n15983), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4604));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12824_4_lut (.I0(n17321), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n17180), .O(n17569));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12824_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i22_3_lut_adj_1733 (.I0(bit_ctr[31]), .I1(n41274), .I2(n4472), 
            .I3(GND_net), .O(n34098));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1733.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4603));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4602));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n1454), .I1(n38647), .I2(n1455), .I3(n1457), 
            .O(n36444));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'ha080;
    SB_LUT4 i6_2_lut (.I0(n1952), .I1(n1953), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4984));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4365), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12818_2_lut (.I0(n38107), .I1(n17561), .I2(GND_net), .I3(GND_net), 
            .O(n17563));   // verilog/coms.v(126[12] 289[6])
    defparam i12818_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_46_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_906_i32_4_lut (.I0(n518), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32_adj_4600));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36309_3_lut (.I0(n32_adj_4600), .I1(n95), .I2(n39_adj_4602), 
            .I3(GND_net), .O(n43163));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36309_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36310_3_lut (.I0(n43163), .I1(n94), .I2(n41_adj_4603), .I3(GND_net), 
            .O(n43164));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36310_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35243_4_lut (.I0(n41_adj_4603), .I1(n39_adj_4602), .I2(n37), 
            .I3(n41389), .O(n42097));
    defparam i35243_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35870_3_lut (.I0(n34_adj_4601), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n42724));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35870_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36121_3_lut (.I0(n43164), .I1(n93), .I2(n43_adj_4604), .I3(GND_net), 
            .O(n42975));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36121_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36305_4_lut (.I0(n42975), .I1(n42724), .I2(n43_adj_4604), 
            .I3(n42097), .O(n43159));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36305_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36306_3_lut (.I0(n43159), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n43160));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36306_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n43160), .I1(n15950), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hceef;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4319));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4598));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4594));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4596));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4595));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_825_i34_4_lut (.I0(n517), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36311_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4595), .I3(GND_net), 
            .O(n43165));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36311_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36312_3_lut (.I0(n43165), .I1(n94), .I2(n43_adj_4596), .I3(GND_net), 
            .O(n43166));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36312_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12821_4_lut (.I0(n17321), .I1(r_Bit_Index[2]), .I2(n4661), 
            .I3(n17180), .O(n17566));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12821_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i35259_4_lut (.I0(n43_adj_4596), .I1(n41_adj_4595), .I2(n39_adj_4594), 
            .I3(n41407), .O(n42113));
    defparam i35259_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_825_i38_3_lut (.I0(n36_adj_4592), .I1(n96), 
            .I2(n39_adj_4594), .I3(GND_net), .O(n38_adj_4593));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36117_3_lut (.I0(n43166), .I1(n93), .I2(n45_adj_4598), .I3(GND_net), 
            .O(n44_adj_4597));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36117_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35868_4_lut (.I0(n44_adj_4597), .I1(n38_adj_4593), .I2(n45_adj_4598), 
            .I3(n42113), .O(n42722));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35868_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n42722), .I1(n15946), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_742_i36_4_lut (.I0(n516), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_742_i40_3_lut (.I0(n38_adj_4590), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4591));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36521_4_lut (.I0(n40_adj_4591), .I1(n36), .I2(n41), .I3(n41417), 
            .O(n43375));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36521_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36522_3_lut (.I0(n43375), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n43376));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36522_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36451_3_lut (.I0(n43376), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n43305));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36451_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n43305), .I1(n15980), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hceef;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13011_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13293), .I3(GND_net), .O(n17756));   // verilog/coms.v(126[12] 289[6])
    defparam i13011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13012_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13293), .I3(GND_net), .O(n17757));   // verilog/coms.v(126[12] 289[6])
    defparam i13012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13013_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13293), .I3(GND_net), .O(n17758));   // verilog/coms.v(126[12] 289[6])
    defparam i13013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13014_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13293), .I3(GND_net), .O(n17759));   // verilog/coms.v(126[12] 289[6])
    defparam i13014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13015_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13293), .I3(GND_net), .O(n17760));   // verilog/coms.v(126[12] 289[6])
    defparam i13015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13016_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13293), .I3(GND_net), .O(n17761));   // verilog/coms.v(126[12] 289[6])
    defparam i13016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13017_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13293), .I3(GND_net), .O(n17762));   // verilog/coms.v(126[12] 289[6])
    defparam i13017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13018_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13293), .I3(GND_net), .O(n17763));   // verilog/coms.v(126[12] 289[6])
    defparam i13018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13019_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13293), .I3(GND_net), .O(n17764));   // verilog/coms.v(126[12] 289[6])
    defparam i13019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13020_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13293), .I3(GND_net), .O(n17765));   // verilog/coms.v(126[12] 289[6])
    defparam i13020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13021_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13293), .I3(GND_net), .O(n17766));   // verilog/coms.v(126[12] 289[6])
    defparam i13021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13022_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13293), .I3(GND_net), .O(n17767));   // verilog/coms.v(126[12] 289[6])
    defparam i13022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13023_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13293), .I3(GND_net), .O(n17768));   // verilog/coms.v(126[12] 289[6])
    defparam i13023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13024_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13293), .I3(GND_net), .O(n17769));   // verilog/coms.v(126[12] 289[6])
    defparam i13024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13025_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13293), .I3(GND_net), .O(n17770));   // verilog/coms.v(126[12] 289[6])
    defparam i13025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13026_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13293), .I3(GND_net), .O(n17771));   // verilog/coms.v(126[12] 289[6])
    defparam i13026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13027_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13293), .I3(GND_net), .O(n17772));   // verilog/coms.v(126[12] 289[6])
    defparam i13027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13028_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13293), .I3(GND_net), .O(n17773));   // verilog/coms.v(126[12] 289[6])
    defparam i13028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13029_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13293), .I3(GND_net), .O(n17774));   // verilog/coms.v(126[12] 289[6])
    defparam i13029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419_adj_4495), .I2(n1382), 
            .I3(GND_net), .O(n1451));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13030_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13293), .I3(GND_net), .O(n17775));   // verilog/coms.v(126[12] 289[6])
    defparam i13030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13031_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13293), .I3(GND_net), .O(n17776));   // verilog/coms.v(126[12] 289[6])
    defparam i13031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13032_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13293), .I3(GND_net), .O(n17777));   // verilog/coms.v(126[12] 289[6])
    defparam i13032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13033_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13293), .I3(GND_net), .O(n17778));   // verilog/coms.v(126[12] 289[6])
    defparam i13033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13034_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13293), .I3(GND_net), .O(n17779));   // verilog/coms.v(126[12] 289[6])
    defparam i13034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13035_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13293), .I3(GND_net), .O(n17780));   // verilog/coms.v(126[12] 289[6])
    defparam i13035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13036_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13293), .I3(GND_net), .O(n17781));   // verilog/coms.v(126[12] 289[6])
    defparam i13036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4473), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4474), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12812_2_lut (.I0(n38107), .I1(n17555), .I2(GND_net), .I3(GND_net), 
            .O(n17557));   // verilog/coms.v(126[12] 289[6])
    defparam i12812_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12815_2_lut (.I0(n38107), .I1(n17558), .I2(GND_net), .I3(GND_net), 
            .O(n17560));   // verilog/coms.v(126[12] 289[6])
    defparam i12815_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418_adj_4494), .I2(n1382), 
            .I3(GND_net), .O(n1450));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12806_2_lut (.I0(n38107), .I1(n17549), .I2(GND_net), .I3(GND_net), 
            .O(n17551));   // verilog/coms.v(126[12] 289[6])
    defparam i12806_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12809_2_lut (.I0(n38107), .I1(n17552), .I2(GND_net), .I3(GND_net), 
            .O(n17554));   // verilog/coms.v(126[12] 289[6])
    defparam i12809_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_46_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4588));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23493_2_lut_4_lut (.I0(communication_counter[30]), .I1(n3_adj_4475), 
            .I2(communication_counter[31]), .I3(n6_adj_4343), .O(n28152));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i23493_2_lut_4_lut.LUT_INIT = 16'hca00;
    SB_LUT4 i34799_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n12_adj_4907), .I3(start), .O(n41299));
    defparam i34799_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 div_46_LessThan_657_i38_4_lut (.I0(n515), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4585));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n12_adj_4907), .I3(state[1]), .O(n36850));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 div_46_LessThan_657_i42_3_lut (.I0(n40_adj_4586), .I1(n96), 
            .I2(n43_adj_4588), .I3(GND_net), .O(n42_adj_4587));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36315_4_lut (.I0(n42_adj_4587), .I1(n38_adj_4585), .I2(n43_adj_4588), 
            .I3(n41429), .O(n43169));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36315_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36316_3_lut (.I0(n43169), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n43170));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36316_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n43170), .I1(n15943), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hceef;
    SB_LUT4 i13037_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13293), .I3(GND_net), .O(n17782));   // verilog/coms.v(126[12] 289[6])
    defparam i13037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23381_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4461), .I3(GND_net), 
            .O(n6_adj_4395));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23381_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i23389_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4395), .I3(GND_net), 
            .O(n8_adj_4391));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23389_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4312), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n514));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1739 (.I0(blink), .I1(n15_adj_4372), .I2(GND_net), 
            .I3(GND_net), .O(blink_N_255));
    defparam i1_2_lut_adj_1739.LUT_INIT = 16'h9999;
    SB_LUT4 i23365_2_lut (.I0(n513), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4919));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23365_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(n85), .I1(n84), .I2(n16011), .I3(GND_net), 
            .O(n15959));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut (.I0(n83), .I1(n82), .I2(n81), .I3(n15998), 
            .O(n16011));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_570_i40_4_lut (.I0(n514), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4582));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_570_i44_3_lut (.I0(n42_adj_4583), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4584));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35862_4_lut (.I0(n44_adj_4584), .I1(n40_adj_4582), .I2(n45), 
            .I3(n41435), .O(n42716));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35862_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n42716), .I1(n15940), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hceef;
    SB_LUT4 i13038_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13293), .I3(GND_net), .O(n17783));   // verilog/coms.v(126[12] 289[6])
    defparam i13038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13231_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n35435), .I3(GND_net), .O(n17976));   // verilog/coms.v(126[12] 289[6])
    defparam i13231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13232_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n35435), .I3(GND_net), .O(n17977));   // verilog/coms.v(126[12] 289[6])
    defparam i13232_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13039_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13293), .I3(GND_net), .O(n17784));   // verilog/coms.v(126[12] 289[6])
    defparam i13039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13040_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13293), .I3(GND_net), .O(n17785));   // verilog/coms.v(126[12] 289[6])
    defparam i13040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13041_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13293), .I3(GND_net), .O(n17786));   // verilog/coms.v(126[12] 289[6])
    defparam i13041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13233_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n35435), .I3(GND_net), .O(n17978));   // verilog/coms.v(126[12] 289[6])
    defparam i13233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1741 (.I0(n82), .I1(n81), .I2(n15998), 
            .I3(GND_net), .O(n16007));
    defparam i1_2_lut_3_lut_adj_1741.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13042_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13293), .I3(GND_net), .O(n17787));   // verilog/coms.v(126[12] 289[6])
    defparam i13042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13043_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13293), .I3(GND_net), .O(n17788));   // verilog/coms.v(126[12] 289[6])
    defparam i13043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13044_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13293), .I3(GND_net), .O(n17789));   // verilog/coms.v(126[12] 289[6])
    defparam i13044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_106[0]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13045_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13293), .I3(GND_net), .O(n17790));   // verilog/coms.v(126[12] 289[6])
    defparam i13045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13046_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13293), .I3(GND_net), .O(n17791));   // verilog/coms.v(126[12] 289[6])
    defparam i13046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13047_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13293), .I3(GND_net), .O(n17792));   // verilog/coms.v(126[12] 289[6])
    defparam i13047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_106[1]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13048_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13293), .I3(GND_net), .O(n17793));   // verilog/coms.v(126[12] 289[6])
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13049_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13293), .I3(GND_net), .O(n17794));   // verilog/coms.v(126[12] 289[6])
    defparam i13049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13050_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13293), .I3(GND_net), .O(n17795));   // verilog/coms.v(126[12] 289[6])
    defparam i13050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13051_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13293), .I3(GND_net), .O(n17796));   // verilog/coms.v(126[12] 289[6])
    defparam i13051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29534_2_lut_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n4_adj_4906), .I3(one_wire_N_513[11]), .O(n36306));
    defparam i29534_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i23349_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_4325), .I3(GND_net), 
            .O(n6_adj_4324));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23349_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i10_4_lut_adj_1742 (.I0(n19_adj_4983), .I1(n15_adj_4985), .I2(n1948), 
            .I3(n1951), .O(n22_adj_4982));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_71_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_106[2]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1743 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n15998));
    defparam i1_2_lut_4_lut_adj_1743.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1744 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n16001));
    defparam i1_2_lut_3_lut_adj_1744.LUT_INIT = 16'hf7f7;
    SB_LUT4 i23333_2_lut (.I0(n512), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23333_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23317_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n511), .I3(n558), 
            .O(n4_adj_4333));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23317_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i11_4_lut_adj_1745 (.I0(n1949), .I1(n22_adj_4982), .I2(n18_adj_4984), 
            .I3(n1950), .O(n1976_adj_4628));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1745.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1254_3_lut (.I0(n1845), .I1(n1912), .I2(n1877), .I3(GND_net), 
            .O(n1944));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_106[3]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23341_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n512), .I3(n558), 
            .O(n4_adj_4325));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23341_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 mux_71_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_106[4]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1746 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n36512));
    defparam i1_3_lut_adj_1746.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1747 (.I0(n2046), .I1(n2054), .I2(n36512), .I3(n2055), 
            .O(n16_adj_4977));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i3_4_lut_adj_1747.LUT_INIT = 16'heaaa;
    SB_LUT4 i9_4_lut_adj_1748 (.I0(n2047), .I1(n2051), .I2(n2048), .I3(n2050), 
            .O(n22_adj_4975));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i9_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n2053), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_4976));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i22_3_lut_adj_1749 (.I0(bit_ctr[22]), .I1(n41275), .I2(n4472), 
            .I3(GND_net), .O(n34104));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1749.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_1750 (.I0(n2044), .I1(n22_adj_4975), .I2(n16_adj_4977), 
            .I3(n2045), .O(n24_adj_4974));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 i12803_2_lut (.I0(n38107), .I1(n17546), .I2(GND_net), .I3(GND_net), 
            .O(n17548));   // verilog/coms.v(126[12] 289[6])
    defparam i12803_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23373_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n513), .I3(n558), 
            .O(n4_adj_4461));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23373_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i12_4_lut_adj_1751 (.I0(n2049), .I1(n24_adj_4974), .I2(n20_adj_4976), 
            .I3(n2052), .O(n2075_adj_4599));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1752 (.I0(color_23__N_164[1]), .I1(n24670), .I2(n1766), 
            .I3(GND_net), .O(n38509));
    defparam i1_3_lut_adj_1752.LUT_INIT = 16'h0404;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(color_23__N_164[7]), .I1(n13_adj_4489), 
            .I2(n11_adj_4490), .I3(n38509), .O(n36415));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_adj_1754 (.I0(n17240), .I1(color[2]), .I2(n36415), 
            .I3(GND_net), .O(n32658));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1754.LUT_INIT = 16'ha8a8;
    SB_LUT4 i24_3_lut (.I0(n41267), .I1(bit_ctr[28]), .I2(n4472), .I3(GND_net), 
            .O(n34082));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_481_i42_4_lut (.I0(n513), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4580));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i36347_3_lut (.I0(n42_adj_4580), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n43201));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36347_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36348_3_lut (.I0(n43201), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n43202));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i36348_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 mux_71_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_106[5]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n43202), .I1(n15937), .I2(n96), .I3(n36150), 
            .O(n806));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'hefce;
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24_3_lut_adj_1756 (.I0(n41266), .I1(bit_ctr[29]), .I2(n4472), 
            .I3(GND_net), .O(n34080));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1756.LUT_INIT = 16'hcaca;
    SB_LUT4 i13052_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13293), 
            .I3(GND_net), .O(n17797));   // verilog/coms.v(126[12] 289[6])
    defparam i13052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13053_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13293), 
            .I3(GND_net), .O(n17798));   // verilog/coms.v(126[12] 289[6])
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_106[6]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13054_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13293), 
            .I3(GND_net), .O(n17799));   // verilog/coms.v(126[12] 289[6])
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13055_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13293), 
            .I3(GND_net), .O(n17800));   // verilog/coms.v(126[12] 289[6])
    defparam i13055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13056_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13293), 
            .I3(GND_net), .O(n17801));   // verilog/coms.v(126[12] 289[6])
    defparam i13056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13057_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13293), 
            .I3(GND_net), .O(n17802));   // verilog/coms.v(126[12] 289[6])
    defparam i13057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13058_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13293), 
            .I3(GND_net), .O(n17803));   // verilog/coms.v(126[12] 289[6])
    defparam i13058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13059_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13293), 
            .I3(GND_net), .O(n17804));   // verilog/coms.v(126[12] 289[6])
    defparam i13059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13060_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13293), 
            .I3(GND_net), .O(n17805));   // verilog/coms.v(126[12] 289[6])
    defparam i13060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_106[7]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13061_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13293), 
            .I3(GND_net), .O(n17806));   // verilog/coms.v(126[12] 289[6])
    defparam i13061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13293), 
            .I3(GND_net), .O(n17808));   // verilog/coms.v(126[12] 289[6])
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13064_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13293), 
            .I3(GND_net), .O(n17809));   // verilog/coms.v(126[12] 289[6])
    defparam i13064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_106[8]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13065_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13293), 
            .I3(GND_net), .O(n17810));   // verilog/coms.v(126[12] 289[6])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13066_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13293), 
            .I3(GND_net), .O(n17811));   // verilog/coms.v(126[12] 289[6])
    defparam i13066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_106[9]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13067_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13293), 
            .I3(GND_net), .O(n17812));   // verilog/coms.v(126[12] 289[6])
    defparam i13067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_106[10]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_106[11]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13068_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13293), 
            .I3(GND_net), .O(n17813));   // verilog/coms.v(126[12] 289[6])
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13069_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13293), 
            .I3(GND_net), .O(n17814));   // verilog/coms.v(126[12] 289[6])
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23480_2_lut_4_lut (.I0(communication_counter[28]), .I1(n5_adj_4473), 
            .I2(communication_counter[31]), .I3(n855), .O(n4_adj_4396));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i23480_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 mux_71_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13070_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13293), 
            .I3(GND_net), .O(n17815));   // verilog/coms.v(126[12] 289[6])
    defparam i13070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13071_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13293), 
            .I3(GND_net), .O(n17816));   // verilog/coms.v(126[12] 289[6])
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_106[12]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13072_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13293), 
            .I3(GND_net), .O(n17817));   // verilog/coms.v(126[12] 289[6])
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13073_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13293), 
            .I3(GND_net), .O(n17818));   // verilog/coms.v(126[12] 289[6])
    defparam i13073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_106[13]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13074_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13293), 
            .I3(GND_net), .O(n17819));   // verilog/coms.v(126[12] 289[6])
    defparam i13074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13075_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13293), 
            .I3(GND_net), .O(n17820));   // verilog/coms.v(126[12] 289[6])
    defparam i13075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13076_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13293), .I3(GND_net), .O(n17821));   // verilog/coms.v(126[12] 289[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13077_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13293), .I3(GND_net), .O(n17822));   // verilog/coms.v(126[12] 289[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_106[14]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13078_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13293), .I3(GND_net), .O(n17823));   // verilog/coms.v(126[12] 289[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13079_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13293), .I3(GND_net), .O(n17824));   // verilog/coms.v(126[12] 289[6])
    defparam i13079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_106[15]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13080_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13293), .I3(GND_net), .O(n17825));   // verilog/coms.v(126[12] 289[6])
    defparam i13080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_106[16]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_106[17]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13081_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13293), .I3(GND_net), .O(n17826));   // verilog/coms.v(126[12] 289[6])
    defparam i13081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13082_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13293), .I3(GND_net), .O(n17827));   // verilog/coms.v(126[12] 289[6])
    defparam i13082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i23309_2_lut (.I0(n511), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4911));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23309_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_70_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_106[18]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_106[19]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4369), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n512));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_46_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_70_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_106[20]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_390_i44_4_lut (.I0(n512), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35858_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n42712));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35858_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_3_lut_adj_1757 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n36470));
    defparam i1_3_lut_adj_1757.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_71_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_106[21]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n42712), .I1(n15933), .I2(n97), .I3(n36148), 
            .O(n671));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hefce;
    SB_LUT4 i4_4_lut_adj_1759 (.I0(n2154), .I1(n2147), .I2(n36470), .I3(n2155), 
            .O(n18_adj_4918));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i4_4_lut_adj_1759.LUT_INIT = 16'heccc;
    SB_LUT4 mux_71_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13083_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13293), .I3(GND_net), .O(n17828));   // verilog/coms.v(126[12] 289[6])
    defparam i13083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_106[22]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1760 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4971));   // verilog/TinyFPGA_B.v(231[5:22])
    defparam i4_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4971), .I2(control_mode[2]), 
            .I3(GND_net), .O(n15922));   // verilog/TinyFPGA_B.v(231[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i23293_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4329));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i23293_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4607));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34486_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n41339));
    defparam i34486_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i2_3_lut_adj_1761 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n15922), .I3(GND_net), .O(n15_adj_4367));   // verilog/TinyFPGA_B.v(231[5:22])
    defparam i2_3_lut_adj_1761.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_46_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4609));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4370), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4367), .I3(n15), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(231[5] 234[10])
    defparam mux_71_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_106[23]), 
            .I2(n15_adj_4313), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(230[5] 234[10])
    defparam mux_70_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_297_i46_4_lut (.I0(n511), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46_adj_4576));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4390));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4389));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4388));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4387));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n46_adj_4576), .I1(n15977), .I2(n98), 
            .I3(n36146), .O(n533));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hefce;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4386));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4385));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n224), .I1(n99), .I2(n15930), .I3(n558), 
            .O(n5_adj_4892));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'h555d;
    SB_LUT4 div_46_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4371), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34665_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n41204));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34665_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n41204), .I1(n15930), .I2(n99), .I3(n5_adj_4892), 
            .O(n392));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hefce;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1765 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n15962));
    defparam i1_2_lut_adj_1765.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1766 (.I0(n81), .I1(n15998), .I2(GND_net), .I3(GND_net), 
            .O(n15992));
    defparam i1_2_lut_adj_1766.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12771_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[19] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17516));   // verilog/coms.v(126[12] 289[6])
    defparam i12771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12772_3_lut (.I0(Kp[0]), .I1(\data_in_frame[2] [0]), .I2(n17068), 
            .I3(GND_net), .O(n17517));   // verilog/coms.v(126[12] 289[6])
    defparam i12772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12773_3_lut (.I0(Ki[0]), .I1(\data_in_frame[3] [0]), .I2(n17068), 
            .I3(GND_net), .O(n17518));   // verilog/coms.v(126[12] 289[6])
    defparam i12773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12774_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17519));   // verilog/coms.v(126[12] 289[6])
    defparam i12774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12775_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17520));   // verilog/coms.v(126[12] 289[6])
    defparam i12775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12776_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n35419), 
            .I3(GND_net), .O(n17521));   // verilog/coms.v(126[12] 289[6])
    defparam i12776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12770_2_lut (.I0(n38107), .I1(n17513), .I2(GND_net), .I3(GND_net), 
            .O(n17515));   // verilog/coms.v(126[12] 289[6])
    defparam i12770_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i22_3_lut_adj_1767 (.I0(bit_ctr[25]), .I1(n41278), .I2(n4472), 
            .I3(GND_net), .O(n34110));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1767.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1768 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n38949));
    defparam i1_2_lut_adj_1768.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12777_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[7] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17522));   // verilog/coms.v(126[12] 289[6])
    defparam i12777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1769 (.I0(n84), .I1(n16011), .I2(GND_net), .I3(GND_net), 
            .O(n16004));
    defparam i1_2_lut_adj_1769.LUT_INIT = 16'hdddd;
    SB_LUT4 i12778_3_lut (.I0(encoder0_position[0]), .I1(n3022), .I2(count_enable), 
            .I3(GND_net), .O(n17523));   // quad.v(35[10] 41[6])
    defparam i12778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i29450_2_lut (.I0(n97_adj_4328), .I1(n737), .I2(GND_net), 
            .I3(GND_net), .O(n36217));
    defparam i29450_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1770 (.I0(n5_adj_4326), .I1(n36217), .I2(\FRAME_MATCHER.i_31__N_2390 ), 
            .I3(n2855), .O(n37799));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1770.LUT_INIT = 16'hbbfb;
    SB_LUT4 div_46_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(\FRAME_MATCHER.i_31__N_2388 ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n37799), .I3(n10454), .O(n34728));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'heafa;
    SB_LUT4 i22_3_lut_adj_1772 (.I0(bit_ctr[24]), .I1(n41277), .I2(n4472), 
            .I3(GND_net), .O(n34108));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1772.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1773 (.I0(bit_ctr[23]), .I1(n41276), .I2(n4472), 
            .I3(GND_net), .O(n34106));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1773.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4384));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12780_3_lut (.I0(encoder1_position[0]), .I1(n2972), .I2(count_enable_adj_4350), 
            .I3(GND_net), .O(n17525));   // quad.v(35[10] 41[6])
    defparam i12780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12781_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n37457), 
            .I3(GND_net), .O(n17526));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1774 (.I0(n17240), .I1(color[19]), .I2(n36429), 
            .I3(GND_net), .O(n32678));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1774.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1_3_lut_adj_1775 (.I0(n17240), .I1(color[18]), .I2(n36429), 
            .I3(GND_net), .O(n32676));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i1_3_lut_adj_1775.LUT_INIT = 16'h8a8a;
    SB_LUT4 i12782_4_lut (.I0(r_SM_Main[2]), .I1(n1), .I2(n25555), .I3(r_SM_Main[1]), 
            .O(n17527));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12782_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i18183_3_lut (.I0(r_SM_Main_adj_5026[0]), .I1(o_Tx_Serial_N_3351), 
            .I2(r_SM_Main_adj_5026[1]), .I3(GND_net), .O(n22916));   // verilog/uart_tx.v(31[16:25])
    defparam i18183_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i18184_3_lut (.I0(tx_o), .I1(n22916), .I2(r_SM_Main_adj_5026[2]), 
            .I3(GND_net), .O(n17528));
    defparam i18184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4383));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n2654), .I1(n38949), .I2(n2655), .I3(n2657), 
            .O(n36563));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'ha080;
    SB_LUT4 i18188_3_lut (.I0(n17108), .I1(r_SM_Main_adj_5026[1]), .I2(tx_active), 
            .I3(GND_net), .O(n17529));   // verilog/uart_tx.v(31[16:25])
    defparam i18188_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i12786_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1144), .I3(GND_net), .O(n17531));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12793_3_lut (.I0(setpoint[0]), .I1(n4378), .I2(n38059), .I3(GND_net), 
            .O(n17538));   // verilog/coms.v(126[12] 289[6])
    defparam i12793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4382));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4381));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4380));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1777 (.I0(color_23__N_164[1]), .I1(n24670), .I2(n1766), 
            .I3(GND_net), .O(n38525));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_3_lut_adj_1777.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4618));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(color_23__N_164[7]), .I1(n13_adj_4489), 
            .I2(n11_adj_4490), .I3(n38525), .O(n36429));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i29551_3_lut (.I0(n36429), .I1(n17240), .I2(color[17]), .I3(GND_net), 
            .O(n36325));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i29551_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i13380_3_lut (.I0(color[12]), .I1(n17240), .I2(n17159), .I3(GND_net), 
            .O(n18125));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i13380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35186_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n42040));
    defparam i35186_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4620));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4631));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13379_3_lut (.I0(color[11]), .I1(n17240), .I2(n17159), .I3(GND_net), 
            .O(n18124));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i13379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35126_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n41980));
    defparam i35126_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13378_3_lut (.I0(color[10]), .I1(n17240), .I2(n17159), .I3(GND_net), 
            .O(n18123));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i13378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4633));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35102_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n41956));
    defparam i35102_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4647));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4643));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(color_23__N_164[4]), .I1(color_23__N_164[6]), 
            .I2(color_23__N_164[2]), .I3(color_23__N_164[0]), .O(n13_adj_4489));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(color_23__N_164[7]), .I1(n13_adj_4489), 
            .I2(n11_adj_4490), .I3(color_23__N_164[1]), .O(n15_adj_4372));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i35083_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n41937));
    defparam i35083_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4645));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4657));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35037_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n41891));
    defparam i35037_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4659));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35049_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n41903));
    defparam i35049_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4661));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i3_2_lut (.I0(color_23__N_164[3]), .I1(color_23__N_164[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4490));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(color_23__N_164[7]), .I1(n11_adj_4490), 
            .I2(color_23__N_164[1]), .I3(n1766), .O(n38485));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n38485), .I1(n15_adj_4372), .I2(n13_adj_4489), 
            .I3(blink), .O(n17159));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'h0a3b;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4379));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4378));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4377));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4376));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1783 (.I0(color_23__N_164[1]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n38565));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_2_lut_adj_1783.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(color_23__N_164[7]), .I1(n13_adj_4489), 
            .I2(n11_adj_4490), .I3(n38565), .O(n17240));   // verilog/TinyFPGA_B.v(78[6:36])
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4375));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13377_3_lut (.I0(color[9]), .I1(n17240), .I2(n17159), .I3(GND_net), 
            .O(n18122));   // verilog/TinyFPGA_B.v(75[8] 98[4])
    defparam i13377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4374));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4373));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12794_3_lut (.I0(quadB_debounced_adj_4349), .I1(reg_B_adj_5035[0]), 
            .I2(n37455), .I3(GND_net), .O(n17539));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36626_4_lut_3_lut (.I0(ID1), .I1(ID2), .I2(ID0), .I3(GND_net), 
            .O(n24670));   // verilog/TinyFPGA_B.v(87[9:10])
    defparam i36626_4_lut_3_lut.LUT_INIT = 16'hbdbd;
    SB_LUT4 i12_4_lut_3_lut (.I0(ID1), .I1(ID2), .I2(ID0), .I3(GND_net), 
            .O(n1766));   // verilog/TinyFPGA_B.v(87[9:10])
    defparam i12_4_lut_3_lut.LUT_INIT = 16'h9494;
    SB_LUT4 div_46_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4674));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_3_lut_adj_1785 (.I0(n35270), .I1(r_Clock_Count[7]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n34716));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1785.LUT_INIT = 16'heaea;
    SB_LUT4 i34988_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n41842));
    defparam i34988_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4347));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4676));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4351));   // verilog/TinyFPGA_B.v(252[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1786 (.I0(n35273), .I1(r_Clock_Count[6]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n34804));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1786.LUT_INIT = 16'heaea;
    SB_LUT4 i34996_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n41850));
    defparam i34996_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1787 (.I0(n35269), .I1(r_Clock_Count[5]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n34912));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1787.LUT_INIT = 16'heaea;
    SB_LUT4 rem_4_i1535_3_lut (.I0(n2254), .I1(n2321), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35387_3_lut (.I0(n2153), .I1(n2220), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1788 (.I0(n35272), .I1(r_Clock_Count[4]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n35000));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1788.LUT_INIT = 16'heaea;
    SB_LUT4 i1_3_lut_adj_1789 (.I0(n35275), .I1(r_Clock_Count[3]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n35090));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1789.LUT_INIT = 16'heaea;
    SB_LUT4 i35389_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i35389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1790 (.I0(n35276), .I1(r_Clock_Count[2]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n35088));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1790.LUT_INIT = 16'heaea;
    SB_LUT4 i1_3_lut_adj_1791 (.I0(n35271), .I1(r_Clock_Count[1]), .I2(n40_adj_4978), 
            .I3(GND_net), .O(n35086));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1791.LUT_INIT = 16'heaea;
    SB_LUT4 rem_4_i1530_3_lut (.I0(n2249), .I1(n2316), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12764_4_lut (.I0(n17330), .I1(r_Bit_Index_adj_5028[2]), .I2(n4683), 
            .I3(n17186), .O(n17509));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12764_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 rem_4_i1529_3_lut (.I0(n2248), .I1(n2315), .I2(n2273_adj_4581), 
            .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4678));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12767_4_lut (.I0(n17330), .I1(r_Bit_Index_adj_5028[1]), .I2(r_Bit_Index_adj_5028[0]), 
            .I3(n17186), .O(n17512));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12767_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4422), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358_adj_4578));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4691));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1467_rep_27_3_lut (.I0(n2154), .I1(n2221), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1467_rep_27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1464_rep_23_3_lut (.I0(n2151), .I1(n2218), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1464_rep_23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36140_3_lut (.I0(n39138), .I1(n1853), .I2(n42403), .I3(GND_net), 
            .O(n2150));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12736_4_lut (.I0(n541), .I1(r_Clock_Count_adj_5027[1]), .I2(n320), 
            .I3(r_SM_Main_adj_5026[2]), .O(n17481));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12736_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i36141_3_lut (.I0(n2150), .I1(n2217), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1462_3_lut (.I0(n2149), .I1(n2216), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1792 (.I0(bit_ctr[26]), .I1(n41279), .I2(n4472), 
            .I3(GND_net), .O(n34112));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1792.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174_adj_4589), 
            .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1793 (.I0(bit_ctr[1]), .I1(n41280), .I2(n4472), 
            .I3(GND_net), .O(n34114));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1793.LUT_INIT = 16'hacac;
    SB_LUT4 i34942_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n41796));
    defparam i34942_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13158_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n35418), 
            .I3(GND_net), .O(n17903));   // verilog/coms.v(126[12] 289[6])
    defparam i13158_3_lut.LUT_INIT = 16'hacac;
    coms setpoint_23__I_0 (.n18036(n18036), .PWMLimit({PWMLimit}), .clk32MHz(clk32MHz), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .GND_net(GND_net), 
         .n18035(n18035), .n18034(n18034), .n18033(n18033), .n18032(n18032), 
         .n18031(n18031), .n18030(n18030), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n18029(n18029), 
         .n18028(n18028), .n18027(n18027), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .n17973(n17973), .\data_in_frame[15] ({\data_in_frame[15] }), .n17902(n17902), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n17972(n17972), .\data_out_frame[16] ({\data_out_frame[16] [7:6], 
         Open_0, \data_out_frame[16] [4], Open_1, Open_2, Open_3, 
         Open_4}), .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n17933(n17933), .\data_in_frame[10] ({\data_in_frame[10] }), .n17932(n17932), 
         .n17901(n17901), .n17931(n17931), .n17930(n17930), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n17929(n17929), .n17928(n17928), .n17927(n17927), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .n17900(n17900), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[4][1] (\data_out_frame[4] [1]), .\data_out_frame[4][0] (\data_out_frame[4] [0]), 
         .n18153(n18153), .setpoint({setpoint}), .n18154(n18154), .n18155(n18155), 
         .n18156(n18156), .n18157(n18157), .n18158(n18158), .n18142(n18142), 
         .n18143(n18143), .n17515(n17515), .n17548(n17548), .n17554(n17554), 
         .n17551(n17551), .n17560(n17560), .n17557(n17557), .n17563(n17563), 
         .n18159(n18159), .n18160(n18160), .n18144(n18144), .n18145(n18145), 
         .n18146(n18146), .n18147(n18147), .n18148(n18148), .n18149(n18149), 
         .n18150(n18150), .n18151(n18151), .n18152(n18152), .n18140(n18140), 
         .n18141(n18141), .n18138(n18138), .n18139(n18139), .n17926(n17926), 
         .n17925(n17925), .n18108(n18108), .VCC_net(VCC_net), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .n17899(n17899), .n18037(n18037), .n18038(n18038), .n18039(n18039), 
         .n18040(n18040), .n18041(n18041), .n18042(n18042), .n17898(n17898), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .n17897(n17897), .n17896(n17896), 
         .n17895(n17895), .n44420(n44420), .n44421(n44421), .n17971(n17971), 
         .n17970(n17970), .\data_in_frame[14] ({\data_in_frame[14] }), .n17969(n17969), 
         .n17968(n17968), .n17967(n17967), .n17966(n17966), .n17894(n17894), 
         .n17893(n17893), .n17892(n17892), .n18048(n18048), .n18049(n18049), 
         .n18046(n18046), .n18047(n18047), .n17891(n17891), .n18043(n18043), 
         .n18044(n18044), .n18045(n18045), .n17890(n17890), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n17889(n17889), .n17888(n17888), .n17887(n17887), .n17886(n17886), 
         .n17885(n17885), .n17884(n17884), .n17883(n17883), .n17882(n17882), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .n17881(n17881), .n17880(n17880), 
         .n17879(n17879), .n17965(n17965), .n17878(n17878), .n17877(n17877), 
         .n17876(n17876), .n17875(n17875), .n17964(n17964), .n17874(n17874), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n17873(n17873), .n17872(n17872), 
         .n17871(n17871), .n17870(n17870), .n17924(n17924), .n17869(n17869), 
         .n17923(n17923), .n17868(n17868), .n17867(n17867), .n17866(n17866), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .n17922(n17922), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n17921(n17921), .\data_out_frame[5] ({\data_out_frame[5] }), .n17920(n17920), 
         .\data_out_frame[4][2] (\data_out_frame[4] [2]), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n17919(n17919), .n17918(n17918), .n17917(n17917), .n17916(n17916), 
         .n17915(n17915), .n17914(n17914), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n17913(n17913), .n17912(n17912), .n17911(n17911), .n17910(n17910), 
         .n17909(n17909), .n17908(n17908), .n17907(n17907), .n17906(n17906), 
         .n17905(n17905), .n17904(n17904), .n17865(n17865), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .n17864(n17864), .n17863(n17863), .n17862(n17862), .n17861(n17861), 
         .n17860(n17860), .n17859(n17859), .n17963(n17963), .n17858(n17858), 
         .\data_in_frame[0] ({\data_in_frame[0] }), .n17857(n17857), .n17856(n17856), 
         .n17855(n17855), .n17854(n17854), .n17853(n17853), .n17852(n17852), 
         .n17851(n17851), .control_mode({control_mode}), .n17850(n17850), 
         .n17849(n17849), .n17848(n17848), .n17962(n17962), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .n17847(n17847), .n17846(n17846), .n17845(n17845), .n17844(n17844), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n17843(n17843), 
         .n17842(n17842), .n17841(n17841), .n17840(n17840), .n17839(n17839), 
         .n17838(n17838), .n17837(n17837), .rx_data_ready(rx_data_ready), 
         .n17836(n17836), .n17835(n17835), .n17974(n17974), .n17961(n17961), 
         .\data_out_frame[16][3] (\data_out_frame[16] [3]), .n17834(n17834), 
         .\data_out_frame[16][5] (\data_out_frame[16] [5]), .n17833(n17833), 
         .n17832(n17832), .n17831(n17831), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n17513(n17513), .n17546(n17546), .n17549(n17549), .n17552(n17552), 
         .n17960(n17960), .n17959(n17959), .n17958(n17958), .n17830(n17830), 
         .n17555(n17555), .n17558(n17558), .n17561(n17561), .n7821(n7821), 
         .n17829(n17829), .n17828(n17828), .n17827(n17827), .n17826(n17826), 
         .n17825(n17825), .n17824(n17824), .n17823(n17823), .n17822(n17822), 
         .n17821(n17821), .n17820(n17820), .n17819(n17819), .n13293(n13293), 
         .n17818(n17818), .n17817(n17817), .n17816(n17816), .n17815(n17815), 
         .n17814(n17814), .n17813(n17813), .n17812(n17812), .n17811(n17811), 
         .n17810(n17810), .n17809(n17809), .n17808(n17808), .n17806(n17806), 
         .\data_out_frame[16][1] (\data_out_frame[16] [1]), .n17805(n17805), 
         .\data_out_frame[16][0] (\data_out_frame[16] [0]), .n17804(n17804), 
         .n17803(n17803), .n17802(n17802), .n17801(n17801), .n17800(n17800), 
         .n17799(n17799), .n17798(n17798), .n17797(n17797), .n17796(n17796), 
         .n17795(n17795), .n17794(n17794), .n17793(n17793), .n17792(n17792), 
         .n17791(n17791), .n17790(n17790), .n17789(n17789), .n17788(n17788), 
         .n17787(n17787), .n17978(n17978), .n17786(n17786), .n17785(n17785), 
         .n17784(n17784), .n17977(n17977), .n17976(n17976), .n17783(n17783), 
         .n17782(n17782), .n17781(n17781), .n17780(n17780), .n17779(n17779), 
         .n17778(n17778), .n17777(n17777), .n17776(n17776), .n17775(n17775), 
         .n17774(n17774), .n17773(n17773), .n17772(n17772), .n17771(n17771), 
         .n17770(n17770), .n17769(n17769), .n17768(n17768), .n17767(n17767), 
         .n17766(n17766), .n17765(n17765), .n17764(n17764), .n17763(n17763), 
         .n17762(n17762), .n17761(n17761), .n17760(n17760), .n17759(n17759), 
         .n17758(n17758), .n17757(n17757), .n17756(n17756), .\FRAME_MATCHER.i_31__N_2390 (\FRAME_MATCHER.i_31__N_2390 ), 
         .n17755(n17755), .n17754(n17754), .n17753(n17753), .n17752(n17752), 
         .n17751(n17751), .n17750(n17750), .n17749(n17749), .n17748(n17748), 
         .n17747(n17747), .n17746(n17746), .n17745(n17745), .n17744(n17744), 
         .n17743(n17743), .ID1(ID1), .ID0(ID0), .n17742(n17742), .n17741(n17741), 
         .n17740(n17740), .n17739(n17739), .n17738(n17738), .n17737(n17737), 
         .n17736(n17736), .n17735(n17735), .n17734(n17734), .n17733(n17733), 
         .n17732(n17732), .ID2(ID2), .n17731(n17731), .n17730(n17730), 
         .n17729(n17729), .\data_in_frame[12] ({\data_in_frame[12] }), .n17728(n17728), 
         .n17727(n17727), .n17726(n17726), .n17725(n17725), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n17724(n17724), .n17723(n17723), .n17722(n17722), .n17721(n17721), 
         .n17720(n17720), .n17719(n17719), .n17718(n17718), .n17717(n17717), 
         .n17716(n17716), .n17715(n17715), .n17714(n17714), .n17713(n17713), 
         .\data_in[3] ({\data_in[3] }), .n17712(n17712), .n17711(n17711), 
         .n17710(n17710), .n17709(n17709), .n17708(n17708), .n17707(n17707), 
         .n17706(n17706), .n17705(n17705), .\data_in[2] ({\data_in[2] }), 
         .n17704(n17704), .n17703(n17703), .n17702(n17702), .n17701(n17701), 
         .n17700(n17700), .n17699(n17699), .n17698(n17698), .n17697(n17697), 
         .\data_in[1] ({\data_in[1] }), .n17696(n17696), .n17695(n17695), 
         .n17694(n17694), .n17693(n17693), .n17692(n17692), .n17691(n17691), 
         .n17690(n17690), .n17689(n17689), .\data_in[0] ({\data_in[0] }), 
         .n17688(n17688), .n17687(n17687), .n17686(n17686), .n17685(n17685), 
         .n17684(n17684), .n17683(n17683), .n17682(n17682), .\Ki[7] (Ki[7]), 
         .n17681(n17681), .\Ki[6] (Ki[6]), .n17680(n17680), .\Ki[5] (Ki[5]), 
         .n17679(n17679), .\Ki[4] (Ki[4]), .n17678(n17678), .\Ki[3] (Ki[3]), 
         .n17677(n17677), .\Ki[2] (Ki[2]), .n17676(n17676), .\Ki[1] (Ki[1]), 
         .n122(n122), .n2855(n2855), .n63(n63_adj_4399), .n5(n5_adj_4468), 
         .n3741(n3741), .\FRAME_MATCHER.state_31__N_2586[2] (\FRAME_MATCHER.state_31__N_2586 [2]), 
         .n17675(n17675), .\Kp[7] (Kp[7]), .n17674(n17674), .\Kp[6] (Kp[6]), 
         .n17673(n17673), .\Kp[5] (Kp[5]), .n17672(n17672), .\Kp[4] (Kp[4]), 
         .n17671(n17671), .\Kp[3] (Kp[3]), .n17670(n17670), .\Kp[2] (Kp[2]), 
         .n17669(n17669), .\Kp[1] (Kp[1]), .n17668(n17668), .gearBoxRatio({gearBoxRatio}), 
         .n17667(n17667), .n17666(n17666), .n17665(n17665), .n17664(n17664), 
         .n17663(n17663), .n17662(n17662), .n17661(n17661), .n17660(n17660), 
         .n17659(n17659), .n17658(n17658), .n17657(n17657), .n17656(n17656), 
         .n17655(n17655), .n17654(n17654), .n17653(n17653), .n17652(n17652), 
         .n17651(n17651), .n17650(n17650), .n17649(n17649), .n17648(n17648), 
         .n17647(n17647), .n17646(n17646), .n17645(n17645), .IntegralLimit({IntegralLimit}), 
         .n17644(n17644), .n17643(n17643), .n17642(n17642), .n17641(n17641), 
         .n17640(n17640), .n17639(n17639), .n17638(n17638), .n17637(n17637), 
         .n17636(n17636), .n17635(n17635), .n17634(n17634), .\FRAME_MATCHER.i_31__N_2388 (\FRAME_MATCHER.i_31__N_2388 ), 
         .n2778(n2778), .n17633(n17633), .n17632(n17632), .n17631(n17631), 
         .n17630(n17630), .n17629(n17629), .n17628(n17628), .n17627(n17627), 
         .n17626(n17626), .n17625(n17625), .n17624(n17624), .n17957(n17957), 
         .n737(n737), .\data_in_frame[18] ({\data_in_frame[18] }), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .n17100(n17100), .n17068(n17068), .n17935(n17935), .n17956(n17956), 
         .n17955(n17955), .n17623(n17623), .n17954(n17954), .n123(n123), 
         .n10454(n10454), .n17953(n17953), .n17952(n17952), .n17951(n17951), 
         .n17950(n17950), .n17949(n17949), .n17948(n17948), .n17947(n17947), 
         .n17946(n17946), .n17945(n17945), .n17944(n17944), .n17943(n17943), 
         .n17942(n17942), .n17941(n17941), .n17975(n17975), .LED_c(LED_c), 
         .n97(n97_adj_4328), .n16(n16_adj_4979), .n7(n7_adj_4311), .n17934(n17934), 
         .\FRAME_MATCHER.state_31__N_2458[1] (\FRAME_MATCHER.state_31__N_2458 [1]), 
         .n17940(n17940), .n17939(n17939), .n17938(n17938), .n17937(n17937), 
         .n17936(n17936), .n17390(n17390), .n17903(n17903), .n4380(n4380), 
         .rx_data({rx_data}), .n4379(n4379), .n4382(n4382), .n4381(n4381), 
         .n17538(n17538), .n34728(n34728), .n17522(n17522), .n17521(n17521), 
         .n17520(n17520), .n17519(n17519), .n17518(n17518), .\Ki[0] (Ki[0]), 
         .n17517(n17517), .\Kp[0] (Kp[0]), .n17516(n17516), .n61(n61_adj_4327), 
         .n4393(n4393), .n4392(n4392), .n4391(n4391), .n4390(n4390), 
         .n4389(n4389), .n4388(n4388), .n4387(n4387), .n4386(n4386), 
         .n4385(n4385), .n4401(n4401), .n4400(n4400), .n35431(n35431), 
         .n35432(n35432), .n35433(n35433), .n35430(n35430), .n35434(n35434), 
         .n35429(n35429), .n38107(n38107), .\duty[10] (duty[10]), .n35428(n35428), 
         .n35435(n35435), .n4378(n4378), .n35419(n35419), .n35423(n35423), 
         .n35420(n35420), .n35416(n35416), .n35417(n35417), .n4384(n4384), 
         .n4383(n4383), .n35421(n35421), .n35422(n35422), .n35418(n35418), 
         .n4399(n4399), .n4398(n4398), .n4397(n4397), .n4396(n4396), 
         .n4395(n4395), .n38059(n38059), .n4394(n4394), .tx_active(tx_active), 
         .n17466(n17466), .\r_Clock_Count[6] (r_Clock_Count_adj_5027[6]), 
         .n17463(n17463), .\r_Clock_Count[7] (r_Clock_Count_adj_5027[7]), 
         .n17481(n17481), .\r_Clock_Count[1] (r_Clock_Count_adj_5027[1]), 
         .n17512(n17512), .r_Bit_Index({r_Bit_Index_adj_5028}), .n17509(n17509), 
         .n18130(n18130), .r_SM_Main({r_SM_Main_adj_5026}), .n18105(n18105), 
         .tx_o(tx_o), .tx_enable(tx_enable), .n19634(n19634), .n17529(n17529), 
         .n17528(n17528), .n541(n541), .n314(n314), .n315(n315), .n320(n320), 
         .o_Tx_Serial_N_3351(o_Tx_Serial_N_3351), .n17108(n17108), .n4683(n4683), 
         .n17186(n17186), .n17330(n17330), .n35270(n35270), .r_Clock_Count({r_Clock_Count}), 
         .n35268(n35268), .n35273(n35273), .n18165(n18165), .n35086(n35086), 
         .n35088(n35088), .n35090(n35090), .n35000(n35000), .n34912(n34912), 
         .n34804(n34804), .n34716(n34716), .n17566(n17566), .r_Bit_Index_adj_14({r_Bit_Index}), 
         .n17569(n17569), .n35004(n35004), .n18111(n18111), .n25741(n25741), 
         .r_SM_Main_adj_15({r_SM_Main}), .n35269(n35269), .r_Rx_Data(r_Rx_Data), 
         .n35272(n35272), .PIN_13_N_105(PIN_13_N_105), .n35275(n35275), 
         .n35276(n35276), .n35271(n35271), .n35274(n35274), .n41248(n41248), 
         .n41247(n41247), .n17576(n17576), .n17575(n17575), .n17574(n17574), 
         .n17573(n17573), .n17572(n17572), .n17571(n17571), .n17570(n17570), 
         .n17527(n17527), .n17180(n17180), .n17321(n17321), .n4661(n4661), 
         .n35374(n35374), .n25555(n25555), .n1(n1), .n24764(n24764), 
         .n4(n4_adj_4366), .n4_adj_12(n4_adj_4368), .n15912(n15912), .n15917(n15917), 
         .n4_adj_13(n4_adj_4362), .n6(n6_adj_4908), .n44844(n44844)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(204[8] 225[4])
    SB_LUT4 i12825_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n24764), 
            .I3(n15912), .O(n17570));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12825_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12826_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n24764), 
            .I3(n15917), .O(n17571));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12826_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_46_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4693));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4695));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12827_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4366), 
            .I3(n15912), .O(n17572));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12827_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12828_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4366), 
            .I3(n15917), .O(n17573));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12828_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12829_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4368), 
            .I3(n15912), .O(n17574));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12829_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12830_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4368), 
            .I3(n15917), .O(n17575));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12830_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i22_3_lut_adj_1794 (.I0(bit_ctr[9]), .I1(n41288), .I2(n4472), 
            .I3(GND_net), .O(n34130));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1794.LUT_INIT = 16'hacac;
    SB_LUT4 i12831_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4362), 
            .I3(n15912), .O(n17576));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12831_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35101_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35101_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i12833_4_lut (.I0(n17312), .I1(state[1]), .I2(state_3__N_362[1]), 
            .I3(n17058), .O(n17578));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12833_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i12846_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n36865), .I3(GND_net), .O(n17591));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12847_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n36865), .I3(GND_net), .O(n17592));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1795 (.I0(bit_ctr[8]), .I1(n41287), .I2(n4472), 
            .I3(GND_net), .O(n34128));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1795.LUT_INIT = 16'hacac;
    SB_LUT4 i12848_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n36865), .I3(GND_net), .O(n17593));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12849_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n36865), .I3(GND_net), .O(n17594));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12850_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n36865), .I3(GND_net), .O(n17595));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12851_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n36865), .I3(GND_net), .O(n17596));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1796 (.I0(bit_ctr[7]), .I1(n41286), .I2(n4472), 
            .I3(GND_net), .O(n34126));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1796.LUT_INIT = 16'hacac;
    SB_LUT4 i12852_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n36865), .I3(GND_net), .O(n17597));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12853_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n36865), .I3(GND_net), .O(n17598));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12854_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n36865), .I3(GND_net), .O(n17599));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2_adj_4329), 
            .I3(n5_adj_4892), .O(n36146));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_4911), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i12855_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n36865), .I3(GND_net), .O(n17600));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35096_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n511), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35096_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i12856_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n36865), .I3(GND_net), .O(n17601));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12857_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n36865), .I3(GND_net), .O(n17602));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12644_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n36865), .I3(GND_net), .O(n17389));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_4333), 
            .I3(n36146), .O(n36148));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i13398_3_lut (.I0(setpoint[6]), .I1(n4384), .I2(n38059), .I3(GND_net), 
            .O(n18143));   // verilog/coms.v(126[12] 289[6])
    defparam i13398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12645_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n17068), .I3(GND_net), .O(n17390));   // verilog/coms.v(126[12] 289[6])
    defparam i12645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34950_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n41804));
    defparam i34950_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i35099_2_lut (.I0(start), .I1(n25771), .I2(GND_net), .I3(GND_net), 
            .O(n41301));   // verilog/neopixel.v(35[12] 117[6])
    defparam i35099_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31_4_lut (.I0(n41301), .I1(n41299), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n34150));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1797 (.I0(control_mode[0]), .I1(n15922), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4313));   // verilog/TinyFPGA_B.v(232[5:22])
    defparam i1_2_lut_3_lut_adj_1797.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36147_3_lut (.I0(n1953), .I1(n2020), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36148_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13397_3_lut (.I0(setpoint[5]), .I1(n4383), .I2(n38059), .I3(GND_net), 
            .O(n18142));   // verilog/coms.v(126[12] 289[6])
    defparam i13397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1798 (.I0(bit_ctr[11]), .I1(n41290), .I2(n4472), 
            .I3(GND_net), .O(n34134));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1798.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1799 (.I0(control_mode[0]), .I1(n15922), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(232[5:22])
    defparam i1_2_lut_3_lut_adj_1799.LUT_INIT = 16'hefef;
    SB_LUT4 i35093_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n512), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35093_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i35549_3_lut (.I0(n2075_adj_4599), .I1(n1976_adj_4628), .I2(n1877), 
            .I3(GND_net), .O(n42403));
    defparam i35549_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1262_rep_44_3_lut (.I0(n1920), .I1(n2019), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n39142));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1262_rep_44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1329_rep_40_3_lut (.I0(n39142), .I1(n2118), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n39138));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1329_rep_40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1800 (.I0(bit_ctr[10]), .I1(n41289), .I2(n4472), 
            .I3(GND_net), .O(n34132));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1800.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_4324), 
            .I3(n36148), .O(n36150));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1395_3_lut (.I0(n2050), .I1(n2117), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1801 (.I0(bit_ctr[13]), .I1(n41292), .I2(n4472), 
            .I3(GND_net), .O(n34138));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1801.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1802 (.I0(bit_ctr[12]), .I1(n41291), .I2(n4472), 
            .I3(GND_net), .O(n34136));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1802.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1803 (.I0(bit_ctr[15]), .I1(n41294), .I2(n4472), 
            .I3(GND_net), .O(n34142));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1803.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1804 (.I0(bit_ctr[14]), .I1(n41293), .I2(n4472), 
            .I3(GND_net), .O(n34140));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1804.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_4325), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2), .I3(n649), 
            .O(n784));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4461), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i22_3_lut_adj_1805 (.I0(bit_ctr[17]), .I1(n41296), .I2(n4472), 
            .I3(GND_net), .O(n34146));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1805.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1806 (.I0(bit_ctr[16]), .I1(n41295), .I2(n4472), 
            .I3(GND_net), .O(n34144));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1806.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_4919), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i15_4_lut_adj_1807 (.I0(n2652), .I1(n30_adj_4897), .I2(n2637_adj_4479), 
            .I3(n2636_adj_4480), .O(n34_adj_4893));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i15_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1808 (.I0(n36563), .I1(n2650), .I2(n2649), .I3(n2648), 
            .O(n32_adj_4895));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i35088_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n513), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i35088_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i24_3_lut_adj_1809 (.I0(n41268), .I1(bit_ctr[19]), .I2(n4472), 
            .I3(GND_net), .O(n34084));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1809.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4395), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i22_3_lut_adj_1810 (.I0(bit_ctr[18]), .I1(n41297), .I2(n4472), 
            .I3(GND_net), .O(n34148));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1810.LUT_INIT = 16'hacac;
    SB_LUT4 i13413_3_lut (.I0(setpoint[21]), .I1(n4399), .I2(n38059), 
            .I3(GND_net), .O(n18158));   // verilog/coms.v(126[12] 289[6])
    defparam i13413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_4391), 
            .I3(n36150), .O(n914));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 i25_4_lut (.I0(n25711), .I1(n36199), .I2(state[0]), .I3(n8_adj_4341), 
            .O(n11_adj_4891));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13412_3_lut (.I0(setpoint[20]), .I1(n4398), .I2(n38059), 
            .I3(GND_net), .O(n18157));   // verilog/coms.v(126[12] 289[6])
    defparam i13412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12858_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n36865), .I3(GND_net), .O(n17603));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i638_3_lut_3_lut (.I0(n938), .I1(n5885), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4711));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1334_3_lut (.I0(n1957), .I1(n2024), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i637_3_lut_3_lut (.I0(n938), .I1(n5884), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34797_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n41650));
    defparam i34797_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4713));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4715));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34836_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n41690));
    defparam i34836_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i639_3_lut_3_lut (.I0(n938), .I1(n5886), .I2(n514), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13411_3_lut (.I0(setpoint[19]), .I1(n4397), .I2(n38059), 
            .I3(GND_net), .O(n18156));   // verilog/coms.v(126[12] 289[6])
    defparam i13411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i636_3_lut_3_lut (.I0(n938), .I1(n5883), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4729));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34738_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n41591));
    defparam i34738_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4731));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4733));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i635_3_lut_3_lut (.I0(n938), .I1(n5882), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34689_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n41542));
    defparam i34689_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4735));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i634_3_lut_3_lut (.I0(n938), .I1(n5881), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13410_3_lut (.I0(setpoint[18]), .I1(n4396), .I2(n38059), 
            .I3(GND_net), .O(n18155));   // verilog/coms.v(126[12] 289[6])
    defparam i13410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12859_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n36865), .I3(GND_net), .O(n17604));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13191_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n35428), .I3(GND_net), .O(n17936));   // verilog/coms.v(126[12] 289[6])
    defparam i13191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13409_3_lut (.I0(setpoint[17]), .I1(n4395), .I2(n38059), 
            .I3(GND_net), .O(n18154));   // verilog/coms.v(126[12] 289[6])
    defparam i13409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13192_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n35428), .I3(GND_net), .O(n17937));   // verilog/coms.v(126[12] 289[6])
    defparam i13192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13193_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n35428), .I3(GND_net), .O(n17938));   // verilog/coms.v(126[12] 289[6])
    defparam i13193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29379_2_lut (.I0(n28152), .I1(n746), .I2(GND_net), .I3(GND_net), 
            .O(n953));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i29379_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13194_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n35431), .I3(GND_net), .O(n17939));   // verilog/coms.v(126[12] 289[6])
    defparam i13194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12860_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n36865), .I3(GND_net), .O(n17605));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4583));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12861_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n36865), .I3(GND_net), .O(n17606));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut_adj_1811 (.I0(n2653), .I1(n2646), .I2(n2651), .I3(n2647), 
            .O(n33_adj_4894));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i14_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1812 (.I0(n2644), .I1(n2642_adj_4477), .I2(n2643_adj_4476), 
            .I3(n2645), .O(n31_adj_4896));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1813 (.I0(n31_adj_4896), .I1(n33_adj_4894), .I2(n32_adj_4895), 
            .I3(n34_adj_4893), .O(n2669));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i18_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4419), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36175_3_lut (.I0(n1853), .I1(n1920), .I2(n1877), .I3(GND_net), 
            .O(n1952));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36176_3_lut (.I0(n1952), .I1(n2019), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34582_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n41435));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34582_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i36272_3_lut (.I0(n1852), .I1(n1919), .I2(n1877), .I3(GND_net), 
            .O(n1951));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36178_3_lut (.I0(n1951), .I1(n2018), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i723_3_lut_3_lut (.I0(n1067), .I1(n5893), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12862_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n36865), .I3(GND_net), .O(n17607));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13195_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n35431), .I3(GND_net), .O(n17940));   // verilog/coms.v(126[12] 289[6])
    defparam i13195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13189_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n35428), .I3(GND_net), .O(n17934));   // verilog/coms.v(126[12] 289[6])
    defparam i13189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976_adj_4628), 
            .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37381_1_lut (.I0(n2966_adj_4400), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n44233));
    defparam i37381_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13408_3_lut (.I0(setpoint[16]), .I1(n4394), .I2(n38059), 
            .I3(GND_net), .O(n18153));   // verilog/coms.v(126[12] 289[6])
    defparam i13408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1267_3_lut (.I0(n1858), .I1(n1925), .I2(n1877), .I3(GND_net), 
            .O(n1957));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1266_3_lut (.I0(n1857), .I1(n1924), .I2(n1877), .I3(GND_net), 
            .O(n1956));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i724_3_lut_3_lut (.I0(n1067), .I1(n5894), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1814 (.I0(bit_ctr[27]), .I1(n41271), .I2(n4472), 
            .I3(GND_net), .O(n34092));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1814.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i725_3_lut_3_lut (.I0(n1067), .I1(n5895), .I2(n515), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1265_3_lut (.I0(n1856), .I1(n1923), .I2(n1877), .I3(GND_net), 
            .O(n1955));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1263_rep_47_3_lut (.I0(n1854), .I1(n1921), .I2(n1877), 
            .I3(GND_net), .O(n1953));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1263_rep_47_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1815 (.I0(n41270), .I1(bit_ctr[21]), .I2(n4472), 
            .I3(GND_net), .O(n34090));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1815.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i722_3_lut_3_lut (.I0(n1067), .I1(n5892), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36181_3_lut (.I0(n1753), .I1(n1820), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13420_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4362), 
            .I3(n15917), .O(n18165));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13420_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i720_3_lut_3_lut (.I0(n1067), .I1(n5890), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4751));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34640_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n41493));
    defparam i34640_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4753));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4755));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34613_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n41466));
    defparam i34613_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i721_3_lut_3_lut (.I0(n1067), .I1(n5891), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i719_3_lut_3_lut (.I0(n1067), .I1(n5889), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13230_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n35435), .I3(GND_net), .O(n17975));   // verilog/coms.v(126[12] 289[6])
    defparam i13230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13196_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n35431), .I3(GND_net), .O(n17941));   // verilog/coms.v(126[12] 289[6])
    defparam i13196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13197_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n35431), .I3(GND_net), .O(n17942));   // verilog/coms.v(126[12] 289[6])
    defparam i13197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13198_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n35431), .I3(GND_net), .O(n17943));   // verilog/coms.v(126[12] 289[6])
    defparam i13198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13199_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n35431), .I3(GND_net), .O(n17944));   // verilog/coms.v(126[12] 289[6])
    defparam i13199_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    SB_LUT4 div_46_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4757));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13385_3_lut_4_lut (.I0(r_SM_Main_adj_5026[2]), .I1(r_SM_Main_adj_5026[0]), 
            .I2(n19634), .I3(r_SM_Main_adj_5026[1]), .O(n18130));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13385_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 div_46_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4774));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34570_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n41423));
    defparam i34570_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4776));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4778));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34540_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n41393));
    defparam i34540_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4780));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13416_3_lut (.I0(quadA_debounced_adj_4348), .I1(reg_B_adj_5035[1]), 
            .I2(n37455), .I3(GND_net), .O(n18161));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4586));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4796));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34576_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n41429));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34576_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i808_3_lut_3_lut (.I0(n1193), .I1(n5904), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i807_3_lut_3_lut (.I0(n1193), .I1(n5903), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4800));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34470_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n41323));
    defparam i34470_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4802));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4798));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i809_3_lut_3_lut (.I0(n1193), .I1(n5905), .I2(n516), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13155_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n35418), 
            .I3(GND_net), .O(n17900));   // verilog/coms.v(126[12] 289[6])
    defparam i13155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1256_3_lut (.I0(n1847), .I1(n1914), .I2(n1877), .I3(GND_net), 
            .O(n1946));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i805_3_lut_3_lut (.I0(n1193), .I1(n5901), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i804_3_lut_3_lut (.I0(n1193), .I1(n5900), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1255_3_lut (.I0(n1846), .I1(n1913), .I2(n1877), .I3(GND_net), 
            .O(n1945));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12718_4_lut (.I0(n541), .I1(r_Clock_Count_adj_5027[7]), .I2(n314), 
            .I3(r_SM_Main_adj_5026[2]), .O(n17463));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12718_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i806_3_lut_3_lut (.I0(n1193), .I1(n5902), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34510_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n41363));
    defparam i34510_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4821));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4825));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35080_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n41934));
    defparam i35080_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4827));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4823));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35130_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n41984));
    defparam i35130_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i23488_2_lut_4_lut (.I0(communication_counter[29]), .I1(n4_adj_4474), 
            .I2(communication_counter[31]), .I3(n4_adj_4396), .O(n6_adj_4343));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i23488_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 div_46_i803_3_lut_3_lut (.I0(n1193), .I1(n5899), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i802_3_lut_3_lut (.I0(n1193), .I1(n5898), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12721_4_lut (.I0(n541), .I1(r_Clock_Count_adj_5027[6]), .I2(n315), 
            .I3(r_SM_Main_adj_5026[2]), .O(n17466));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12721_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4590));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34564_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n41417));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34564_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i890_3_lut_3_lut (.I0(n1316), .I1(n5915), .I2(n1299), 
            .I3(GND_net), .O(n1419));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i889_3_lut_3_lut (.I0(n1316), .I1(n5914), .I2(n1298), 
            .I3(GND_net), .O(n1418));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i891_3_lut_3_lut (.I0(n1316), .I1(n5916), .I2(n517), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i887_3_lut_3_lut (.I0(n1316), .I1(n5912), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i886_3_lut_3_lut (.I0(n1316), .I1(n5911), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i888_3_lut_3_lut (.I0(n1316), .I1(n5913), .I2(n1297), 
            .I3(GND_net), .O(n1417));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i885_3_lut_3_lut (.I0(n1316), .I1(n5910), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i884_3_lut_3_lut (.I0(n1316), .I1(n5909), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i883_3_lut_3_lut (.I0(n1316), .I1(n5908), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1816 (.I0(bit_ctr[6]), .I1(n41285), .I2(n4472), 
            .I3(GND_net), .O(n34124));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1816.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4426), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34554_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n41407));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34554_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i22_3_lut_adj_1817 (.I0(bit_ctr[5]), .I1(n41284), .I2(n4472), 
            .I3(GND_net), .O(n34122));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1817.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1818 (.I0(bit_ctr[4]), .I1(n41283), .I2(n4472), 
            .I3(GND_net), .O(n34120));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1818.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_4951));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22_3_lut_adj_1819 (.I0(bit_ctr[3]), .I1(n41282), .I2(n4472), 
            .I3(GND_net), .O(n34118));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1819.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758_adj_4458), .I1(n1825), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1198_3_lut (.I0(n1757_adj_4457), .I1(n1824), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910), .I2(n2867), .I3(GND_net), 
            .O(n2942));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837), .I1(n2904), .I2(n2867), .I3(GND_net), 
            .O(n2936));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1935_3_lut (.I0(n2846), .I1(n2913), .I2(n2867), .I3(GND_net), 
            .O(n2945));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1937_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), .I3(GND_net), 
            .O(n2947));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1942_3_lut (.I0(n2853), .I1(n2920), .I2(n2867), .I3(GND_net), 
            .O(n2952_adj_4407));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1941_3_lut (.I0(n2852), .I1(n2919), .I2(n2867), .I3(GND_net), 
            .O(n2951_adj_4408));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4592));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i1938_3_lut (.I0(n2849), .I1(n2916), .I2(n2867), .I3(GND_net), 
            .O(n2948));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908), .I2(n2867), .I3(GND_net), 
            .O(n2940));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1936_3_lut (.I0(n2847), .I1(n2914), .I2(n2867), .I3(GND_net), 
            .O(n2946));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867), .I3(GND_net), 
            .O(n2950_adj_4409));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912), .I2(n2867), .I3(GND_net), 
            .O(n2944));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907), .I2(n2867), .I3(GND_net), 
            .O(n2939));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1943_3_lut (.I0(n2854), .I1(n2921), .I2(n2867), .I3(GND_net), 
            .O(n2953_adj_4406));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1939_3_lut (.I0(n2850), .I1(n2917), .I2(n2867), .I3(GND_net), 
            .O(n2949_adj_4410));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838), .I1(n2905), .I2(n2867), .I3(GND_net), 
            .O(n2937));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i970_3_lut_3_lut (.I0(n1436), .I1(n5927), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839), .I1(n2906), .I2(n2867), .I3(GND_net), 
            .O(n2938));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909), .I2(n2867), .I3(GND_net), 
            .O(n2941));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835), .I1(n2902), .I2(n2867), .I3(GND_net), 
            .O(n2934));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836), .I1(n2903), .I2(n2867), .I3(GND_net), 
            .O(n2935));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911), .I2(n2867), .I3(GND_net), 
            .O(n2943));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i967_3_lut_3_lut (.I0(n1436), .I1(n5924), .I2(n1417), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i968_3_lut_3_lut (.I0(n1436), .I1(n5925), .I2(n1418), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1820 (.I0(bit_ctr[2]), .I1(n41281), .I2(n4472), 
            .I3(GND_net), .O(n34116));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1820.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i964_3_lut_3_lut (.I0(n1436), .I1(n5921), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i963_3_lut_3_lut (.I0(n1436), .I1(n5920), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i966_3_lut_3_lut (.I0(n1436), .I1(n5923), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13182_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n35429), 
            .I3(GND_net), .O(n17927));   // verilog/coms.v(126[12] 289[6])
    defparam i13182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i971_3_lut_3_lut (.I0(n1436), .I1(n5928), .I2(n518), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13183_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n35429), 
            .I3(GND_net), .O(n17928));   // verilog/coms.v(126[12] 289[6])
    defparam i13183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i965_3_lut_3_lut (.I0(n1436), .I1(n5922), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867), .I3(GND_net), 
            .O(n2955_adj_4404));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855_adj_4434), .I1(n2922), .I2(n2867), 
            .I3(GND_net), .O(n2954_adj_4405));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2858), .I1(n2925), .I2(n2867), .I3(GND_net), 
            .O(n2957_adj_4402));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13184_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n35429), 
            .I3(GND_net), .O(n17929));   // verilog/coms.v(126[12] 289[6])
    defparam i13184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857), .I1(n2924), .I2(n2867), .I3(GND_net), 
            .O(n2956_adj_4403));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13185_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n35429), 
            .I3(GND_net), .O(n17930));   // verilog/coms.v(126[12] 289[6])
    defparam i13185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i962_3_lut_3_lut (.I0(n1436), .I1(n5919), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1821 (.I0(n2956_adj_4403), .I1(n2957_adj_4402), 
            .I2(n2958_adj_4401), .I3(GND_net), .O(n36517));
    defparam i1_3_lut_adj_1821.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1822 (.I0(n2933), .I1(n2954_adj_4405), .I2(n36517), 
            .I3(n2955_adj_4404), .O(n26_adj_4965));
    defparam i4_4_lut_adj_1822.LUT_INIT = 16'heaaa;
    SB_LUT4 i14_4_lut_adj_1823 (.I0(n2943), .I1(n2935), .I2(n2934), .I3(n2941), 
            .O(n36_adj_4963));
    defparam i14_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1824 (.I0(n2938), .I1(n2937), .I2(n2949_adj_4410), 
            .I3(n2953_adj_4406), .O(n34_adj_4964));
    defparam i12_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1825 (.I0(n2939), .I1(n36_adj_4963), .I2(n26_adj_4965), 
            .I3(n2944), .O(n40_adj_4959));
    defparam i18_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1826 (.I0(n2950_adj_4409), .I1(n2946), .I2(n2940), 
            .I3(n2948), .O(n38_adj_4961));
    defparam i16_4_lut_adj_1826.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2951_adj_4408), .I1(n34_adj_4964), .I2(n2952_adj_4407), 
            .I3(GND_net), .O(n39_adj_4960));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1827 (.I0(n2947), .I1(n2945), .I2(n2936), .I3(n2942), 
            .O(n37_adj_4962));
    defparam i15_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1828 (.I0(n37_adj_4962), .I1(n39_adj_4960), .I2(n38_adj_4961), 
            .I3(n40_adj_4959), .O(n2966_adj_4400));
    defparam i21_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i969_3_lut_3_lut (.I0(n1436), .I1(n5926), .I2(n1419), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34536_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n41389));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam i34536_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4601));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1047_3_lut_3_lut (.I0(n1553), .I1(n5939), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13186_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n35428), .I3(GND_net), .O(n17931));   // verilog/coms.v(126[12] 289[6])
    defparam i13186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1045_3_lut_3_lut (.I0(n1553), .I1(n5937), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13156_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n35418), 
            .I3(GND_net), .O(n17901));   // verilog/coms.v(126[12] 289[6])
    defparam i13156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13187_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n35428), .I3(GND_net), .O(n17932));   // verilog/coms.v(126[12] 289[6])
    defparam i13187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1042_3_lut_3_lut (.I0(n1553), .I1(n5934), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1048_3_lut_3_lut (.I0(n1553), .I1(n5940), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1041_3_lut_3_lut (.I0(n1553), .I1(n5933), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13188_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n35428), .I3(GND_net), .O(n17933));   // verilog/coms.v(126[12] 289[6])
    defparam i13188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1049_3_lut_3_lut (.I0(n1553), .I1(n5941), .I2(n519), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1044_3_lut_3_lut (.I0(n1553), .I1(n5936), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1043_3_lut_3_lut (.I0(n1553), .I1(n5935), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1040_3_lut_3_lut (.I0(n1553), .I1(n5932), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1039_3_lut_3_lut (.I0(n1553), .I1(n5931), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1046_3_lut_3_lut (.I0(n1553), .I1(n5938), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1124_3_lut_3_lut (.I0(n1667), .I1(n5954), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1118_3_lut_3_lut (.I0(n1667), .I1(n5948), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1122_3_lut_3_lut (.I0(n1667), .I1(n5952), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10_4_lut_adj_1829 (.I0(n2148), .I1(n2149), .I2(n2150), .I3(n2151), 
            .O(n24_adj_4916));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i10_4_lut_adj_1829.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1123_3_lut_3_lut (.I0(n1667), .I1(n5953), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1121_3_lut_3_lut (.I0(n1667), .I1(n5951), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1117_3_lut_3_lut (.I0(n1667), .I1(n5947), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1125_3_lut_3_lut (.I0(n1667), .I1(n5955), .I2(n520), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1120_3_lut_3_lut (.I0(n1667), .I1(n5950), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4542));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755_adj_4455), .I1(n1822), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_4950));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4541));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1195_3_lut (.I0(n1754_adj_4454), .I1(n1821), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4540));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4539));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36183_3_lut (.I0(n1653_adj_4460), .I1(n1720), .I2(n1679), 
            .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36184_3_lut (.I0(n1752), .I1(n1819), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i36184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_4949));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4538));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4537));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4536));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(173[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4535));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778_adj_4818), 
            .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1119_3_lut_3_lut (.I0(n1667), .I1(n5949), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1115_3_lut_3_lut (.I0(n1667), .I1(n5945), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1116_3_lut_3_lut (.I0(n1667), .I1(n5946), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1114_3_lut_3_lut (.I0(n1667), .I1(n5944), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1195_3_lut_3_lut (.I0(n1778), .I1(n5966), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1187_3_lut_3_lut (.I0(n1778), .I1(n5958), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1196_3_lut_3_lut (.I0(n1778), .I1(n5967), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1197_3_lut_3_lut (.I0(n1778), .I1(n5968), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1198_3_lut_3_lut (.I0(n1778), .I1(n5969), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n6_adj_4908), 
            .I3(r_Rx_Data), .O(n40_adj_4978));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hdccc;
    SB_LUT4 i8_4_lut_adj_1831 (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_4917));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i8_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n18067(n18067), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n18068(n18068), .n18069(n18069), .n18070(n18070), 
            .n18071(n18071), .n18072(n18072), .n18056(n18056), .n18057(n18057), 
            .n18058(n18058), .n18059(n18059), .n18060(n18060), .n18061(n18061), 
            .n18062(n18062), .n18063(n18063), .n18064(n18064), .n18065(n18065), 
            .n18066(n18066), .n18054(n18054), .n18055(n18055), .n18052(n18052), 
            .n18053(n18053), .n18050(n18050), .n18051(n18051), .data_o({quadA_debounced, 
            quadB_debounced}), .n2998({n2999, n3000, n3001, n3002, 
            n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
            n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
            n3019, n3020, n3021, n3022}), .GND_net(GND_net), .n17523(n17523), 
            .count_enable(count_enable), .n18101(n18101), .reg_B({reg_B}), 
            .n37457(n37457), .PIN_2_c_0(PIN_2_c_0), .n17526(n17526), .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(256[15] 261[4])
    SB_LUT4 div_46_i1192_3_lut_3_lut (.I0(n1778), .I1(n5963), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34499_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41313));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i34499_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_i1191_3_lut_3_lut (.I0(n1778), .I1(n5962), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i3_4_lut_adj_1832 (.I0(r_SM_Main[2]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(n44844), .O(n38007));
    defparam i3_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i34816_4_lut (.I0(n41313), .I1(r_SM_Main[0]), .I2(n35374), 
            .I3(r_Clock_Count[7]), .O(n41310));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i34816_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 div_46_i1194_3_lut_3_lut (.I0(n1778), .I1(n5965), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1199_3_lut_3_lut (.I0(n1778), .I1(n5970), .I2(n521), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1193_3_lut_3_lut (.I0(n1778), .I1(n5964), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i2_4_lut_adj_1833 (.I0(n41310), .I1(n40_adj_4978), .I2(n38007), 
            .I3(r_SM_Main[1]), .O(n35268));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_4_lut_adj_1833.LUT_INIT = 16'h0322;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n18075(n18075), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n18076(n18076), .n18077(n18077), .n18078(n18078), 
            .n18079(n18079), .n18080(n18080), .n18081(n18081), .n18095(n18095), 
            .n18096(n18096), .n18097(n18097), .n18093(n18093), .n18094(n18094), 
            .n18091(n18091), .n18092(n18092), .n18089(n18089), .n18090(n18090), 
            .n18087(n18087), .n18088(n18088), .n18085(n18085), .n18086(n18086), 
            .n18082(n18082), .n18083(n18083), .n18084(n18084), .n2948({n2949, 
            n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
            n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
            n2966, n2967, n2968, n2969, n2970, n2971, n2972}), 
            .GND_net(GND_net), .data_o({quadA_debounced_adj_4348, quadB_debounced_adj_4349}), 
            .n17525(n17525), .count_enable(count_enable_adj_4350), .n18161(n18161), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B_adj_5035}), .PIN_7_c_1(PIN_7_c_1), 
            .n37455(n37455), .n17539(n17539)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(264[15] 269[4])
    SB_LUT4 i12_4_lut_adj_1834 (.I0(n2145), .I1(n24_adj_4916), .I2(n18_adj_4918), 
            .I3(n2146), .O(n26_adj_4915));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i12_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1189_3_lut_3_lut (.I0(n1778), .I1(n5960), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1190_3_lut_3_lut (.I0(n1778), .I1(n5961), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1188_3_lut_3_lut (.I0(n1778), .I1(n5959), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1270_3_lut_3_lut (.I0(n1886), .I1(n5985), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_4948));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_4947));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_4946));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1261_3_lut_3_lut (.I0(n1886), .I1(n5976), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_4_lut_adj_1835 (.I0(n2153), .I1(n26_adj_4915), .I2(n22_adj_4917), 
            .I3(n2152), .O(n2174_adj_4589));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i13_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1259_3_lut_3_lut (.I0(n1886), .I1(n5974), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1258_3_lut_3_lut (.I0(n1886), .I1(n5973), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4534));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075_adj_4599), 
            .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13200_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n35431), .I3(GND_net), .O(n17945));   // verilog/coms.v(126[12] 289[6])
    defparam i13200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4533));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1269_3_lut_3_lut (.I0(n1886), .I1(n5984), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_4945));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i27_3_lut (.I0(n1138), .I1(n36199), .I2(state[0]), .I3(GND_net), 
            .O(n19_adj_4890));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1267_3_lut_3_lut (.I0(n1886), .I1(n5982), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4427), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1268_3_lut_3_lut (.I0(n1886), .I1(n5983), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_4944));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1265_3_lut_3_lut (.I0(n1886), .I1(n5980), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4532));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4943));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1266_3_lut_3_lut (.I0(n1886), .I1(n5981), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757_adj_4457));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13201_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n35431), .I3(GND_net), .O(n17946));   // verilog/coms.v(126[12] 289[6])
    defparam i13201_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13202_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n35432), .I3(GND_net), .O(n17947));   // verilog/coms.v(126[12] 289[6])
    defparam i13202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13203_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n35432), .I3(GND_net), .O(n17948));   // verilog/coms.v(126[12] 289[6])
    defparam i13203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4942));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13204_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n35432), .I3(GND_net), .O(n17949));   // verilog/coms.v(126[12] 289[6])
    defparam i13204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13205_3_lut (.I0(\data_in_frame[12] [3]), .I1(rx_data[3]), 
            .I2(n35432), .I3(GND_net), .O(n17950));   // verilog/coms.v(126[12] 289[6])
    defparam i13205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13206_3_lut (.I0(\data_in_frame[12] [4]), .I1(rx_data[4]), 
            .I2(n35432), .I3(GND_net), .O(n17951));   // verilog/coms.v(126[12] 289[6])
    defparam i13206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13207_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n35432), .I3(GND_net), .O(n17952));   // verilog/coms.v(126[12] 289[6])
    defparam i13207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13208_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n35432), .I3(GND_net), .O(n17953));   // verilog/coms.v(126[12] 289[6])
    defparam i13208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1264_3_lut_3_lut (.I0(n1886), .I1(n5979), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1271_3_lut_3_lut (.I0(n1886), .I1(n5986), .I2(n522), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1263_3_lut_3_lut (.I0(n1886), .I1(n5978), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1260_3_lut_3_lut (.I0(n1886), .I1(n5975), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1262_3_lut_3_lut (.I0(n1886), .I1(n5977), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1340_3_lut_3_lut (.I0(n1991), .I1(n6002), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1332_3_lut_3_lut (.I0(n1991), .I1(n5994), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1836 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n36545));
    defparam i1_3_lut_adj_1836.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_i1331_3_lut_3_lut (.I0(n1991), .I1(n5993), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1328_3_lut_3_lut (.I0(n1991), .I1(n5990), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1330_3_lut_3_lut (.I0(n1991), .I1(n5992), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4941));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755_adj_4455));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4531));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4530));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1329_3_lut_3_lut (.I0(n1991), .I1(n5991), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1327_3_lut_3_lut (.I0(n1991), .I1(n5989), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1335_3_lut_3_lut (.I0(n1991), .I1(n5997), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13209_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n35432), .I3(GND_net), .O(n17954));   // verilog/coms.v(126[12] 289[6])
    defparam i13209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12863_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n36865), .I3(GND_net), .O(n17608));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12864_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n36865), .I3(GND_net), .O(n17609));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12865_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n36865), .I3(GND_net), .O(n17610));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12866_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n36865), .I3(GND_net), .O(n17611));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12866_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12867_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n36865), .I3(GND_net), .O(n17612));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12867_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1336_3_lut_3_lut (.I0(n1991), .I1(n5998), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12868_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n36865), .I3(GND_net), .O(n17613));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12868_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12869_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n36865), .I3(GND_net), .O(n17614));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12869_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1334_3_lut_3_lut (.I0(n1991), .I1(n5996), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1339_3_lut_3_lut (.I0(n1991), .I1(n6001), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1338_3_lut_3_lut (.I0(n1991), .I1(n6000), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12870_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n36865), .I3(GND_net), .O(n17615));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12870_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12871_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n36865), .I3(GND_net), .O(n17616));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12871_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12872_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n36865), .I3(GND_net), .O(n17617));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12872_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12873_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n36865), .I3(GND_net), .O(n17618));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12873_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12874_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n36865), .I3(GND_net), .O(n17619));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12875_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n36865), .I3(GND_net), .O(n17620));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12875_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1337_3_lut_3_lut (.I0(n1991), .I1(n5999), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12876_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n36865), .I3(GND_net), .O(n17621));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24_3_lut_adj_1837 (.I0(n41269), .I1(bit_ctr[20]), .I2(n4472), 
            .I3(GND_net), .O(n34088));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1837.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4940));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12878_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n17068), .I3(GND_net), .O(n17623));   // verilog/coms.v(126[12] 289[6])
    defparam i12878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1341_3_lut_3_lut (.I0(n1991), .I1(n6003), .I2(n523), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1333_3_lut_3_lut (.I0(n1991), .I1(n5995), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1404_3_lut_3_lut (.I0(n2093), .I1(n6016), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1401_3_lut_3_lut (.I0(n2093), .I1(n6013), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37316_1_lut_2_lut (.I0(n3362), .I1(n10218), .I2(GND_net), 
            .I3(GND_net), .O(n44170));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i37316_1_lut_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_46_i1400_3_lut_3_lut (.I0(n2093), .I1(n6012), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1399_3_lut_3_lut (.I0(n2093), .I1(n6011), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1396_3_lut_3_lut (.I0(n2093), .I1(n6008), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1395_3_lut_3_lut (.I0(n2093), .I1(n6007), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1398_3_lut_3_lut (.I0(n2093), .I1(n6010), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1394_3_lut_3_lut (.I0(n2093), .I1(n6006), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1402_3_lut_3_lut (.I0(n2093), .I1(n6014), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1403_3_lut_3_lut (.I0(n2093), .I1(n6015), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1405_3_lut_3_lut (.I0(n2093), .I1(n6017), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1408_3_lut_3_lut (.I0(n2093), .I1(n6020), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1406_3_lut_3_lut (.I0(n2093), .I1(n6018), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1407_3_lut_3_lut (.I0(n2093), .I1(n6019), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1409_3_lut_3_lut (.I0(n2093), .I1(n6021), .I2(n524), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1397_3_lut_3_lut (.I0(n2093), .I1(n6009), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1470_3_lut_3_lut (.I0(n2192), .I1(n6035), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1459_3_lut_3_lut (.I0(n2192), .I1(n6024), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1471_3_lut_3_lut (.I0(n2192), .I1(n6036), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1467_3_lut_3_lut (.I0(n2192), .I1(n6032), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1465_3_lut_3_lut (.I0(n2192), .I1(n6030), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1475_3_lut_3_lut (.I0(n2192), .I1(n6040), .I2(n525), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1463_3_lut_3_lut (.I0(n2192), .I1(n6028), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1462_3_lut_3_lut (.I0(n2192), .I1(n6027), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1461_3_lut_3_lut (.I0(n2192), .I1(n6026), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1464_3_lut_3_lut (.I0(n2192), .I1(n6029), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1460_3_lut_3_lut (.I0(n2192), .I1(n6025), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1474_3_lut_3_lut (.I0(n2192), .I1(n6039), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1472_3_lut_3_lut (.I0(n2192), .I1(n6037), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1473_3_lut_3_lut (.I0(n2192), .I1(n6038), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1469_3_lut_3_lut (.I0(n2192), .I1(n6034), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1468_3_lut_3_lut (.I0(n2192), .I1(n6033), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1466_3_lut_3_lut (.I0(n2192), .I1(n6031), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1528_3_lut_3_lut (.I0(n2288), .I1(n6049), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1522_3_lut_3_lut (.I0(n2288), .I1(n6043), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1525_3_lut_3_lut (.I0(n2288), .I1(n6046), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1523_3_lut_3_lut (.I0(n2288), .I1(n6044), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1526_3_lut_3_lut (.I0(n2288), .I1(n6047), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1527_3_lut_3_lut (.I0(n2288), .I1(n6048), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1537_3_lut_3_lut (.I0(n2288), .I1(n6058), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1536_3_lut_3_lut (.I0(n2288), .I1(n6057), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1524_3_lut_3_lut (.I0(n2288), .I1(n6045), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1532_3_lut_3_lut (.I0(n2288), .I1(n6053), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1531_3_lut_3_lut (.I0(n2288), .I1(n6052), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1530_3_lut_3_lut (.I0(n2288), .I1(n6051), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1539_3_lut_3_lut (.I0(n2288), .I1(n6060), .I2(n526), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1529_3_lut_3_lut (.I0(n2288), .I1(n6050), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15930), 
            .O(n249));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_46_i1534_3_lut_3_lut (.I0(n2288), .I1(n6055), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754_adj_4454));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1127_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), .I3(GND_net), 
            .O(n1753));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam rem_4_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4529));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4528));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1838 (.I0(n97), .I1(n96), .I2(n95), .I3(n15940), 
            .O(n15977));
    defparam i1_2_lut_4_lut_adj_1838.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1839 (.I0(n96), .I1(n95), .I2(n15940), 
            .I3(GND_net), .O(n15933));
    defparam i1_2_lut_3_lut_adj_1839.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1535_3_lut_3_lut (.I0(n2288), .I1(n6056), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1840 (.I0(n94), .I1(n93), .I2(n92), .I3(n15946), 
            .O(n15940));
    defparam i1_2_lut_4_lut_adj_1840.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1841 (.I0(n93), .I1(n92), .I2(n15946), 
            .I3(GND_net), .O(n15943));
    defparam i1_2_lut_3_lut_adj_1841.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1533_3_lut_3_lut (.I0(n2288), .I1(n6054), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1842 (.I0(n91), .I1(n90), .I2(n89), .I3(n15986), 
            .O(n15946));
    defparam i1_2_lut_4_lut_adj_1842.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1538_3_lut_3_lut (.I0(n2288), .I1(n6059), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1595_3_lut_3_lut (.I0(n2381), .I1(n6075), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11_4_lut_adj_1843 (.I0(n2248), .I1(n2253), .I2(n2252), .I3(n2249), 
            .O(n26_adj_4910));   // verilog/TinyFPGA_B.v(78[6:33])
    defparam i11_4_lut_adj_1843.LUT_INIT = 16'hfffe;
    \pwm(32000000,20000,32000000,23,1)  PWM (.GND_net(GND_net), .VCC_net(VCC_net), 
            .PIN_19_c_0(PIN_19_c_0), .CLK_c(CLK_c), .\half_duty_new[0] (half_duty_new[0]), 
            .n18136(n18136), .\half_duty[0][6] (\half_duty[0] [6]), .n18137(n18137), 
            .\half_duty[0][7] (\half_duty[0] [7]), .n18134(n18134), .\half_duty[0][4] (\half_duty[0] [4]), 
            .n18135(n18135), .\half_duty[0][5] (\half_duty[0] [5]), .n18132(n18132), 
            .\half_duty[0][2] (\half_duty[0] [2]), .n18133(n18133), .\half_duty[0][3] (\half_duty[0] [3]), 
            .n18131(n18131), .\half_duty[0][1] (\half_duty[0] [1]), .n1144(n1144), 
            .\half_duty[0][0] (\half_duty[0] [0]), .\half_duty_new[1] (half_duty_new[1]), 
            .\half_duty_new[2] (half_duty_new[2]), .\half_duty_new[3] (half_duty_new[3]), 
            .\half_duty_new[4] (half_duty_new[4]), .\half_duty_new[5] (half_duty_new[5]), 
            .\half_duty_new[6] (half_duty_new[6]), .\half_duty_new[7] (half_duty_new[7]), 
            .pwm_setpoint({pwm_setpoint}), .n17531(n17531)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(155[43] 161[3])
    motorControl control (.GND_net(GND_net), .IntegralLimit({IntegralLimit}), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Ki[6] (Ki[6]), .\Kp[4] (Kp[4]), 
            .\Ki[7] (Ki[7]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .duty({duty}), .PWMLimit({PWMLimit}), .clk32MHz(clk32MHz), 
            .VCC_net(VCC_net), .n44224(n44224), .motor_state({motor_state}), 
            .n25(n25), .setpoint({setpoint})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(236[16] 249[4])
    SB_LUT4 div_46_i1584_3_lut_3_lut (.I0(n2381), .I1(n6064), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1583_3_lut_3_lut (.I0(n2381), .I1(n6063), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1587_3_lut_3_lut (.I0(n2381), .I1(n6067), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1588_3_lut_3_lut (.I0(n2381), .I1(n6068), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1585_3_lut_3_lut (.I0(n2381), .I1(n6065), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1586_3_lut_3_lut (.I0(n2381), .I1(n6066), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1601_3_lut_3_lut (.I0(n2381), .I1(n6081), .I2(n527), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1844 (.I0(n90), .I1(n89), .I2(n15986), 
            .I3(GND_net), .O(n15950));
    defparam i1_2_lut_3_lut_adj_1844.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1596_3_lut_3_lut (.I0(n2381), .I1(n6076), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1845 (.I0(n88), .I1(n87), .I2(n86), .I3(n15959), 
            .O(n15986));
    defparam i1_2_lut_4_lut_adj_1845.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1592_3_lut_3_lut (.I0(n2381), .I1(n6072), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1600_3_lut_3_lut (.I0(n2381), .I1(n6080), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1599_3_lut_3_lut (.I0(n2381), .I1(n6079), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1598_3_lut_3_lut (.I0(n2381), .I1(n6078), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1846 (.I0(n87), .I1(n86), .I2(n15959), 
            .I3(GND_net), .O(n15989));
    defparam i1_2_lut_3_lut_adj_1846.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1591_3_lut_3_lut (.I0(n2381), .I1(n6071), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1590_3_lut_3_lut (.I0(n2381), .I1(n6070), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1597_3_lut_3_lut (.I0(n2381), .I1(n6077), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1589_3_lut_3_lut (.I0(n2381), .I1(n6069), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1594_3_lut_3_lut (.I0(n2381), .I1(n6074), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1593_3_lut_3_lut (.I0(n2381), .I1(n6073), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1655_3_lut_3_lut (.I0(n2471), .I1(n6097), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1642_3_lut_3_lut (.I0(n2471), .I1(n6084), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1643_3_lut_3_lut (.I0(n2471), .I1(n6085), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1847 (.I0(n86), .I1(n15959), .I2(GND_net), .I3(GND_net), 
            .O(n15953));
    defparam i1_2_lut_adj_1847.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_i1644_3_lut_3_lut (.I0(n2471), .I1(n6086), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(252[21:53])
    defparam div_46_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, bit_ctr, VCC_net, 
            GND_net, timer, n41296, n19, n34116, n34118, n34120, 
            n34122, n34124, n34090, n34092, n34148, n34084, n34144, 
            n34146, n34140, n34142, n34136, n34138, n34132, n34134, 
            n34126, n34128, n34130, n34114, n34112, n34106, n34108, 
            n34110, n34080, n34082, n34104, n34098, n34094, n34096, 
            n41295, n41284, \neo_pixel_transmitter.t0 , n41294, n41283, 
            n41293, n41292, n4, start, \state[0] , n106, \state[1] , 
            n35266, n41291, n41282, n41290, n41281, n41289, n41288, 
            n34088, n17621, n17620, n17619, n17618, n17617, n17616, 
            n17615, n17614, n17613, n17612, n17611, n17610, n17609, 
            n17608, n41280, PIN_8_c, n36850, n41274, n41273, n17607, 
            n41287, n17606, n17605, n17604, n17603, n41266, n11, 
            n41286, n41267, n17058, n17312, n41271, n41272, n41285, 
            n34150, n17389, n17602, n17601, n17600, n17599, n17598, 
            n17597, n17596, n17595, n17594, n17593, n17592, n17591, 
            n17578, n41279, n41278, n41277, n41276, \one_wire_N_513[11] , 
            n41275, \one_wire_N_513[8] , n41270, \one_wire_N_513[7] , 
            \one_wire_N_513[6] , \one_wire_N_513[5] , n41269, n41268, 
            n41297, n25771, n1138, n12, n8, \color[20] , \color[4] , 
            \color[10] , \color[11] , \color[9] , \color[17] , \color[18] , 
            \color[19] , \color[1] , \color[2] , \color[3] , \color[12] , 
            \state_3__N_362[1] , n4472, n25711, n36199, n36306, n36865) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output [31:0]bit_ctr;
    input VCC_net;
    input GND_net;
    output [31:0]timer;
    output n41296;
    input n19;
    input n34116;
    input n34118;
    input n34120;
    input n34122;
    input n34124;
    input n34090;
    input n34092;
    input n34148;
    input n34084;
    input n34144;
    input n34146;
    input n34140;
    input n34142;
    input n34136;
    input n34138;
    input n34132;
    input n34134;
    input n34126;
    input n34128;
    input n34130;
    input n34114;
    input n34112;
    input n34106;
    input n34108;
    input n34110;
    input n34080;
    input n34082;
    input n34104;
    input n34098;
    input n34094;
    input n34096;
    output n41295;
    output n41284;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output n41294;
    output n41283;
    output n41293;
    output n41292;
    output n4;
    output start;
    output \state[0] ;
    output n106;
    output \state[1] ;
    input n35266;
    output n41291;
    output n41282;
    output n41290;
    output n41281;
    output n41289;
    output n41288;
    input n34088;
    input n17621;
    input n17620;
    input n17619;
    input n17618;
    input n17617;
    input n17616;
    input n17615;
    input n17614;
    input n17613;
    input n17612;
    input n17611;
    input n17610;
    input n17609;
    input n17608;
    output n41280;
    output PIN_8_c;
    input n36850;
    output n41274;
    output n41273;
    input n17607;
    output n41287;
    input n17606;
    input n17605;
    input n17604;
    input n17603;
    output n41266;
    input n11;
    output n41286;
    output n41267;
    output n17058;
    output n17312;
    output n41271;
    output n41272;
    output n41285;
    input n34150;
    input n17389;
    input n17602;
    input n17601;
    input n17600;
    input n17599;
    input n17598;
    input n17597;
    input n17596;
    input n17595;
    input n17594;
    input n17593;
    input n17592;
    input n17591;
    input n17578;
    output n41279;
    output n41278;
    output n41277;
    output n41276;
    output \one_wire_N_513[11] ;
    output n41275;
    output \one_wire_N_513[8] ;
    output n41270;
    output \one_wire_N_513[7] ;
    output \one_wire_N_513[6] ;
    output \one_wire_N_513[5] ;
    output n41269;
    output n41268;
    output n41297;
    output n25771;
    output n1138;
    output n12;
    output n8;
    input \color[20] ;
    input \color[4] ;
    input \color[10] ;
    input \color[11] ;
    input \color[9] ;
    input \color[17] ;
    input \color[18] ;
    input \color[19] ;
    input \color[1] ;
    input \color[2] ;
    input \color[3] ;
    input \color[12] ;
    output \state_3__N_362[1] ;
    output n4472;
    output n25711;
    output n36199;
    input n36306;
    output n36865;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n29989, n3099, n3116, n29990, n29750, n2007, n2027, n29751, 
        n2107, n2008, n29749, n3199, n3100, n29988, n3200, n3101, 
        n29987, n2108, n2009, n44218, n29748, \neo_pixel_transmitter.done_N_570 , 
        n38137, n3201, n3102, n29986, n2109;
    wire [31:0]n133;
    
    wire n29242, n3202, n3103, n29985, n1994, n1895, n1928, n29747, 
        n29241, n29233, n29234, n28634;
    wire [31:0]n1;
    
    wire n28635, n1995, n1896, n29746, n29232, n3203, n3104, n29984, 
        n1996, n1897, n29745, n3204, n3105, n29983, n1997, n1898, 
        n29744, n29240, n3205, n3106, n29982, n29239, n29231, 
        n28443, n29230, n1998, n1899, n29743, n3206, n3107, n29981, 
        n1999, n1900, n29742, n29229, n29238, n29228;
    wire [31:0]one_wire_N_513;
    
    wire n28633, n29227, n28632, n2907, n2909, n33, n3207, n3108, 
        n29980, n2000, n1901, n29741, n29237, n3208, n3109, n44217, 
        n29979, n2001, n1902, n29740, n3209, n2002, n1903, n29739, 
        n2003, n1904, n29738, n3083, n2984, n3017, n29978, n3084, 
        n2985, n29977, n2004, n1905, n29737, n29236, n2005, n1906, 
        n29736, n2900, n2891, n2897, n2888, n41, n2906, n2887, 
        n2892, n38, n2896, n2885, n2905, n2902, n43, n2899, 
        n2890, n2898, n2908, n40, n29226, n2889, n2901, n46, 
        n2886, n2894, n2895, n2903, n39, n2904, n2893, n47, 
        n2918, n3085, n2986, n29976, n30771, n28631, n4_c, n44220, 
        n29225, n29224, n29223, n1699, n1709, n17, n1698, n1707, 
        n1703, n1705, n21, n1704, n1701, n1708, n20, n1702, 
        n1697, n24, n1700, n1706, n1730, n29222, n1829, n44221, 
        n29221, n29220, n28444, n1509, n25571, n1506, n1502, n1501, 
        n18, n1503, n1507, n16, n29219, n1504, n1508, n1505, 
        n20_adj_4175, n29218, n29217, n1500, n1499, n1532, n29216, 
        n3086, n2987, n29975, n2006, n1907, n29735, n29215, n29214, 
        n29213, n29212, n28442, n28431, n1908, n29734, n29235, 
        n3087, n2988, n29974, n1909, n44219, n29733, n3088, n2989, 
        n29973, n3089, n2990, n29972, n1796, n29732, n3090, n2991, 
        n29971, n1797, n29731, n3091, n2992, n29970, n1798, n29730, 
        n1799, n29729, n3092, n2993, n29969, n1800, n29728, n3093, 
        n2994, n29968, n3094, n2995, n29967, n1801, n29727, n1802, 
        n29726, n1806, n1804, n24_adj_4177, n1807, n1808, n22, 
        n1803, n1805, n23, n3095, n2996, n29966, n28432, n1809, 
        n21_adj_4178, n29725, n3096, n2997, n29965, n29724, n3097, 
        n2998, n29964, n29723, n29722, n3098, n2999, n29963, n3000, 
        n29962, n29721, n3001, n29961, n2791, n2795, n2802, n2799, 
        n40_adj_4179, n29720, n2786, n2801, n2807, n2803, n38_adj_4180, 
        n3002, n29960, n29719, n3003, n29959, n2793, n2806, n2794, 
        n2787, n39_adj_4181, n29718, n29717, n3004, n29958, n29716, 
        n3005, n29957, n3006, n29956, n26, n19_adj_4182, n16_adj_4183, 
        n29715, n2796, n2798, n2788, n2800, n37, n24_adj_4184, 
        n28, n3007, n29955, n29714, n2808, n2809, n36, n2805, 
        n2804, n35, n46_adj_4185, n3008, n29954, n29713, n28441, 
        n3009, n29953, n2797, n2789, n2790, n2792, n41_adj_4186, 
        n29712, n29711, n2596, n2609, n28_adj_4187, n2595, n2590, 
        n2592, n2599, n35_adj_4188, n2593, n2605, n2589, n2608, 
        n34, n2606, n2603, n40_adj_4189, n2591, n2588, n2594, 
        n2598, n38_adj_4190, n29710, n2602, n2607, n39_adj_4191, 
        n2597, n2600, n2601, n2604, n37_adj_4192, n2621, n2819, 
        n29952, n2720, n44230, n29951, n29709, n29950, n28430, 
        n29708, n29949, n29948, n29707, n29947, n44222, n29706, 
        n28440, n29946, n1598, n1631, n29705, n1599, n29704, n29945, 
        n29944, n1600, n29703, n44223, n29943, n1601, n29702, 
        n29942, n1602, n29701, n29941, n1603, n29700, n1604, n29699, 
        n29940, n28439, n1605, n29698, n29939, n1606, n29697, 
        n29938, n1607, n29696, n1608, n29695, n29937, n1609, n44225, 
        n29694, n29936, n29935, n29934, n29933, n29932, n29931, 
        n29930, n29929, n29928, n29927, n29926, n29925, n25417, 
        n35446, n21_adj_4194, n23_adj_4195, n22_adj_4196, n24_adj_4197, 
        n36_adj_4198, n25, n27, n26_adj_4199, n28_adj_4200, n37_adj_4201, 
        n29_adj_4202, n30_adj_4203, n15928, n112, n29924, n29923, 
        n1409, n25569, n1405, n1403, n1406, n16_adj_4204, n1402, 
        n1404, n1400, n1407, n17_adj_4205, n1408, n1401, n1433, 
        n29922, n29921, n29920, n2693, n2704, n28_adj_4206, n2699, 
        n2706, n2694, n2691, n38_adj_4207, n2709, n25667, n2701, 
        n2696, n2697, n36_adj_4208, n28438, n2700, n2705, n42, 
        n29919, n2702, n2690, n2689, n2708, n40_adj_4209, n2687, 
        n2703, n2695, n41_adj_4210, n2688, n2698, n2692, n2707, 
        n39_adj_4211, n28511, n29918, n28510, n28429, n29917, n28437, 
        n29916, n29915, n29914, n25553, n708, n29913, n29912, 
        n29911, n29910, n29909, n28509, n29908, n44227, n28508, 
        n29907, n29906, n28507, n28428, n29905, n29904, n29903, 
        n28506, n28606, n20_adj_4212, n13, n18_adj_4213, n29902, 
        n22_adj_4214, n29901, n29900, n28436, n29899, n29898, n28605, 
        n29897, n29896, n28505, n29895, n28604, n29894, n29893, 
        n29892, n29891, n29890, n28603, n29889, n28504, n29888, 
        n29887, n29886, n28602, n29885, n29884, n29883, n28601, 
        n28503, n29882, n28502, n28435, n29881, n29880, n29879, 
        n29878, n29877, n29876, n29875, n44229, n28501, n29874, 
        n28427, n29873, n29872, \neo_pixel_transmitter.done_N_576 , 
        n17075, n29871, n29870, n29869, n29868, n29867, n28600, 
        n29866, n29865, n29864, n29863, n28599, n29862, n28598, 
        n29861, n28661, n28457, n28660, n29860, n28659, n44231, 
        n28597, n44232, n29859, n28456, n28658, n2489, n2522, 
        n29858, n2490, n29857, n2491, n29856, n28657, n28656, 
        n2492, n29855, n28655, n28654, n2493, n29854, n28653, 
        n2494, n29853, n2495, n29852, n28652, n2496, n29851, n2497, 
        n29850, n28651, n2498, n29849, n2499, n29848, n2500, n29847, 
        n2501, n29846, n2502, n29845, n2503, n29844, n2504, n29843, 
        n2505, n29842, n2506, n29841, n28650, n2507, n29840, n2508, 
        n29839, n25651, n28_adj_4217, n26_adj_4218, n27_adj_4219, 
        n25_adj_4220, n36_adj_4221, n46_adj_4222, n42_adj_4223, n33_adj_4224, 
        n43_adj_4225, n50, n48, n49, n47_adj_4226, n2509, n44234, 
        n29838, n28434, n28649, n2390, n2423, n29837, n2391, n29836, 
        n2392, n29835, n2393, n29834;
    wire [31:0]n971;
    
    wire n905, n28867, n906, n28866, n2394, n29833, n2395, n29832, 
        n2396, n29831, n2397, n29830, n36288, n28865, n2398, n29829, 
        n17229, n28864, n28648, n2399, n29828, n2400, n29827, 
        n28455, n2401, n29826, n2402, n29825, n28433, n14415, 
        n28863, n2403, n29824, n28454, n2404, n29823;
    wire [3:0]state_3__N_362;
    
    wire n2405, n29822, n2406, n29821, n2407, n29820, n1103, n4_adj_4228, 
        n1037, n28862, n1104, n1005, n28861, n2408, n29819, n1105, 
        n1006, n28860, n2409, n44235, n29818, n28647, n28453, 
        n1106, n1007, n28859, n1107, n1008, n28858, n1108, n1009, 
        n44236, n28857, n1109, n2291, n2324, n29817, n2292, n29816, 
        n2293, n29815, n2294, n29814, n2295, n29813, n2296, n29812, 
        n2297, n29811, n28452, n2298, n29810, n2299, n29809, n2300, 
        n29808, n2301, n29807, n2302, n29806, n2303, n29805, n28646, 
        n28645, n2304, n29804, n2305, n29803, n2306, n29802, n28451, 
        n2307, n29801, n2308, n29800, n2309, n44237, n29799, n2192, 
        n2225, n29798, n2193, n29797, n2194, n29796, n2195, n29795, 
        n1202, n1136, n28807, n1203, n28806, n28644, n2196, n29794, 
        n1204, n28805, n1205, n28804, n1206, n28803, n2197, n29793, 
        n1207, n28802, n1208, n44239, n28801, n1209, n2198, n29792, 
        n2199, n29791, n28643, n2200, n29790, n2201, n29789, n2202, 
        n29788, n2203, n29787, n1301, n1235, n28792, n1302, n28791, 
        n1303, n28790, n1304, n28789, n1305, n28788, n1306, n28787, 
        n2204, n29786, n28642, n2205, n29785, n1307, n28786, n1308, 
        n44240, n28785, n1309, n2206, n29784, n1334, n28784, n28783, 
        n28782, n2207, n29783, n28781, n28780, n28779, n28778, 
        n28450, n28777, n44241, n28776, n28449, n2208, n29782, 
        n2209, n44238, n29781, n28641, n2093, n2126, n29780, n2094, 
        n29779, n2095, n29778, n2096, n29777, n2097, n29776, n2098, 
        n29775, n2099, n29774, n2100, n29773, n2101, n29772, n28640, 
        n28448, n28639, n28638, n2102, n29771, n2103, n29770, 
        n28447, n2104, n29769, n3182, n30005, n2105, n29768, n28637, 
        n3183, n30004, n2106, n29767, n28636, n3184, n30003, n29766, 
        n29765, n28446, n3185, n30002, n44242, n29764, n3186, 
        n30001, n3187, n30000, n29763, n29762, n29761, n28445, 
        n3188, n29999, n29760, n29759, n3189, n29998, n29758, 
        n3190, n29997, n29757, n3191, n29996, n3192, n29995, n29756, 
        n29755, n3193, n29994, n29754, n3194, n29993, n29753, 
        n3195, n29992, n3196, n29991, n29752, n3197, n3198, n37679, 
        n30650, n15775, n4_adj_4242, n15887, n25777, n36211, n838, 
        n13454, n36197, n608, n36189, n36154, n60, n14417, n807, 
        n18_adj_4244, n25655, n30_adj_4245, n28_adj_4246, n29_adj_4247, 
        n27_adj_4248, n10_adj_4249, n12_adj_4250, n16_adj_4251, n14_adj_4252, 
        n9_adj_4253, n25561, n12_adj_4254, n28_adj_4255, n32_adj_4256, 
        n30_adj_4257, n31_adj_4258, n29_adj_4259, n22_adj_4260, n30_adj_4261, 
        n34_adj_4262, n32_adj_4263, n33_adj_4264, n31_adj_4265, n31958, 
        n39093, n39101, n6_adj_4266, n41043, n25645, n48_adj_4267, 
        n46_adj_4268, n47_adj_4269, n45, n44, n43_adj_4270, n54, 
        n49_adj_4271, n25737, n1141, n41235, n41231, n9_adj_4273, 
        n45277, n42667, n18_adj_4274, n45271, n17_adj_4275, n3_adj_4276, 
        n2_adj_4277, n42462, n39195;
    wire [4:0]color_bit_N_556;
    
    wire n41303, n43057, n22_adj_4278, n32_adj_4279, n25671, n36_adj_4280, 
        n34_adj_4281, n35_adj_4282, n33_adj_4283, n26_adj_4284, n33_adj_4285, 
        n22_adj_4286, n38_adj_4287, n36_adj_4288, n37_adj_4289, n35_adj_4290, 
        n30_adj_4291, n48_adj_4292, n46_adj_4293, n47_adj_4294, n45_adj_4295, 
        n44_adj_4296, n43_adj_4297, n54_adj_4298, n49_adj_4299, n4443, 
        n31_adj_4300, n41_adj_4301, n40_adj_4302, n45_adj_4303, n44_adj_4304, 
        n43_adj_4305, n47_adj_4306, n49_adj_4307, n6_adj_4308, n6_adj_4309, 
        n36207, n37638;
    
    SB_CARRY mod_5_add_2143_13 (.CI(n29989), .I0(n3099), .I1(n3116), .CO(n29990));
    SB_CARRY mod_5_add_1406_5 (.CI(n29750), .I0(n2007), .I1(n2027), .CO(n29751));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n29749), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n29749), .I0(n2008), .I1(n2027), .CO(n29750));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n29988), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n29988), .I0(n3100), .I1(n3116), .CO(n29989));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n29987), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n29987), .I0(n3101), .I1(n3116), .CO(n29988));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n44218), 
            .I3(n29748), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n38137), .D(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_3 (.CI(n29748), .I0(n2009), .I1(n44218), .CO(n29749));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n29986), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n44218), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1200_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n29242), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_10 (.CI(n29986), .I0(n3102), .I1(n3116), .CO(n29987));
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n44218), 
            .CO(n29748));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n29985), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n29747), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1200_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n29241), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_24 (.CI(n29233), .I0(GND_net), .I1(timer[22]), 
            .CO(n29234));
    SB_CARRY sub_14_add_2_6 (.CI(n28634), .I0(timer[4]), .I1(n1[4]), .CO(n28635));
    SB_CARRY mod_5_add_2143_9 (.CI(n29985), .I0(n3103), .I1(n3116), .CO(n29986));
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n29746), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1200_add_4_32 (.CI(n29241), .I0(GND_net), .I1(timer[30]), 
            .CO(n29242));
    SB_LUT4 timer_1200_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n29232), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n29984), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n29746), .I0(n1896), .I1(n1928), .CO(n29747));
    SB_CARRY timer_1200_add_4_23 (.CI(n29232), .I0(GND_net), .I1(timer[21]), 
            .CO(n29233));
    SB_CARRY mod_5_add_2143_8 (.CI(n29984), .I0(n3104), .I1(n3116), .CO(n29985));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n29745), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n29983), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n29745), .I0(n1897), .I1(n1928), .CO(n29746));
    SB_CARRY mod_5_add_2143_7 (.CI(n29983), .I0(n3105), .I1(n3116), .CO(n29984));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n29744), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1200_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n29240), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_31 (.CI(n29240), .I0(GND_net), .I1(timer[29]), 
            .CO(n29241));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n29982), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n29744), .I0(n1898), .I1(n1928), .CO(n29745));
    SB_LUT4 timer_1200_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n29239), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1200_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n29231), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_19_lut (.I0(n19), .I1(bit_ctr[17]), .I2(GND_net), .I3(n28443), 
            .O(n41296)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1200_add_4_22 (.CI(n29231), .I0(GND_net), .I1(timer[20]), 
            .CO(n29232));
    SB_LUT4 timer_1200_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n29230), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_21 (.CI(n29230), .I0(GND_net), .I1(timer[19]), 
            .CO(n29231));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n29743), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n29982), .I0(n3106), .I1(n3116), .CO(n29983));
    SB_CARRY mod_5_add_1339_13 (.CI(n29743), .I0(n1899), .I1(n1928), .CO(n29744));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n29981), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n29742), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1200_add_4_30 (.CI(n29239), .I0(GND_net), .I1(timer[28]), 
            .CO(n29240));
    SB_LUT4 timer_1200_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n29229), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_20 (.CI(n29229), .I0(GND_net), .I1(timer[18]), 
            .CO(n29230));
    SB_LUT4 timer_1200_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n29238), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1200_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n29228), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n28633), .O(one_wire_N_513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_19 (.CI(n29228), .I0(GND_net), .I1(timer[17]), 
            .CO(n29229));
    SB_CARRY timer_1200_add_4_29 (.CI(n29238), .I0(GND_net), .I1(timer[27]), 
            .CO(n29239));
    SB_LUT4 timer_1200_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n29227), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n28633), .I0(timer[3]), .I1(n1[3]), .CO(n28634));
    SB_CARRY timer_1200_add_4_18 (.CI(n29227), .I0(GND_net), .I1(timer[16]), 
            .CO(n29228));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n28632), .O(one_wire_N_513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_2143_5 (.CI(n29981), .I0(n3107), .I1(n3116), .CO(n29982));
    SB_CARRY mod_5_add_1339_12 (.CI(n29742), .I0(n1900), .I1(n1928), .CO(n29743));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n29980), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n29980), .I0(n3108), .I1(n3116), .CO(n29981));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n29741), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1200_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n29237), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_11 (.CI(n29741), .I0(n1901), .I1(n1928), .CO(n29742));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n44217), 
            .I3(n29979), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n29740), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n29740), .I0(n1902), .I1(n1928), .CO(n29741));
    SB_CARRY mod_5_add_2143_3 (.CI(n29979), .I0(n3109), .I1(n44217), .CO(n29980));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n44217), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n29739), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1200_add_4_28 (.CI(n29237), .I0(GND_net), .I1(timer[26]), 
            .CO(n29238));
    SB_CARRY mod_5_add_1339_9 (.CI(n29739), .I0(n1903), .I1(n1928), .CO(n29740));
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n44217), 
            .CO(n29979));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n29738), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n29978), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n29738), .I0(n1904), .I1(n1928), .CO(n29739));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n29977), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n29737), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1200_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n29236), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_27 (.CI(n29977), .I0(n2985), .I1(n3017), .CO(n29978));
    SB_CARRY mod_5_add_1339_7 (.CI(n29737), .I0(n1905), .I1(n1928), .CO(n29738));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n29736), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1200_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n29226), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut (.I0(n41), .I1(n33), .I2(n2889), .I3(n2901), .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n34116));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i14_4_lut (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n34118));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n34120));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n34122));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n34124));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i22_4_lut (.I0(n43), .I1(n2904), .I2(n38), .I3(n2893), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_4 (.CI(n28632), .I0(timer[2]), .I1(n1[2]), .CO(n28633));
    SB_CARRY timer_1200_add_4_17 (.CI(n29226), .I0(GND_net), .I1(timer[15]), 
            .CO(n29227));
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n34090));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n34092));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n34148));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n34084));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n34144));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n34146));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n34140));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n34142));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n34136));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n34138));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n34132));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n34134));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n34126));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n34128));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n34130));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n34114));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n34112));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n34106));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n34108));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n34110));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(VCC_net), 
            .D(n34080));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(VCC_net), 
            .D(n34082));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n34104));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n29976), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n34098));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n34094));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n34096));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_c), .I1(timer[1]), .I2(n1[1]), 
            .I3(n28631), .O(n30771)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i37368_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44220));
    defparam i37368_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1200_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n29225), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_16 (.CI(n29225), .I0(GND_net), .I1(timer[14]), 
            .CO(n29226));
    SB_LUT4 timer_1200_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n29224), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_15 (.CI(n29224), .I0(GND_net), .I1(timer[13]), 
            .CO(n29225));
    SB_LUT4 timer_1200_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n29223), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_14 (.CI(n29223), .I0(GND_net), .I1(timer[12]), 
            .CO(n29224));
    SB_LUT4 i4_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n17));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n21), .I1(n17), .I2(n1702), .I3(n1697), .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n1700), .I1(n24), .I2(n20), .I3(n1706), .O(n1730));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1200_add_4_27 (.CI(n29236), .I0(GND_net), .I1(timer[25]), 
            .CO(n29237));
    SB_LUT4 timer_1200_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n29222), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37369_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44221));
    defparam i37369_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1200_add_4_13 (.CI(n29222), .I0(GND_net), .I1(timer[11]), 
            .CO(n29223));
    SB_LUT4 timer_1200_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n29221), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_26 (.CI(n29976), .I0(n2986), .I1(n3017), .CO(n29977));
    SB_CARRY timer_1200_add_4_12 (.CI(n29221), .I0(GND_net), .I1(timer[10]), 
            .CO(n29222));
    SB_LUT4 timer_1200_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n29220), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_11 (.CI(n29220), .I0(GND_net), .I1(timer[9]), 
            .CO(n29221));
    SB_CARRY add_21_19 (.CI(n28443), .I0(bit_ctr[17]), .I1(GND_net), .CO(n28444));
    SB_LUT4 i20842_2_lut (.I0(bit_ctr[20]), .I1(n1509), .I2(GND_net), 
            .I3(GND_net), .O(n25571));
    defparam i20842_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut (.I0(n1506), .I1(n1502), .I2(n25571), .I3(n1501), 
            .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1339_6 (.CI(n29736), .I0(n1906), .I1(n1928), .CO(n29737));
    SB_LUT4 i5_2_lut (.I0(n1503), .I1(n1507), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 timer_1200_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n29219), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_10 (.CI(n29219), .I0(GND_net), .I1(timer[8]), 
            .CO(n29220));
    SB_LUT4 i9_4_lut (.I0(n1504), .I1(n18), .I2(n1508), .I3(n1505), 
            .O(n20_adj_4175));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1200_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n29218), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_9 (.CI(n29218), .I0(GND_net), .I1(timer[7]), 
            .CO(n29219));
    SB_LUT4 timer_1200_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n29217), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_8 (.CI(n29217), .I0(GND_net), .I1(timer[6]), 
            .CO(n29218));
    SB_LUT4 i10_4_lut (.I0(n1500), .I1(n20_adj_4175), .I2(n16), .I3(n1499), 
            .O(n1532));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1200_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n29216), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n29975), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n29735), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n29735), .I0(n1907), .I1(n1928), .CO(n29736));
    SB_CARRY timer_1200_add_4_7 (.CI(n29216), .I0(GND_net), .I1(timer[5]), 
            .CO(n29217));
    SB_LUT4 timer_1200_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n29215), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_6 (.CI(n29215), .I0(GND_net), .I1(timer[4]), 
            .CO(n29216));
    SB_LUT4 timer_1200_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n29214), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_5 (.CI(n29214), .I0(GND_net), .I1(timer[3]), 
            .CO(n29215));
    SB_LUT4 timer_1200_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n29213), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_4 (.CI(n29213), .I0(GND_net), .I1(timer[2]), 
            .CO(n29214));
    SB_LUT4 timer_1200_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n29212), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1200_add_4_3 (.CI(n29212), .I0(GND_net), .I1(timer[1]), 
            .CO(n29213));
    SB_LUT4 timer_1200_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_18_lut (.I0(n19), .I1(bit_ctr[16]), .I2(GND_net), .I3(n28442), 
            .O(n41295)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n28431), 
            .O(n41284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1200_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n29212));
    SB_CARRY mod_5_add_2076_25 (.CI(n29975), .I0(n2987), .I1(n3017), .CO(n29976));
    SB_CARRY sub_14_add_2_3 (.CI(n28631), .I0(timer[1]), .I1(n1[1]), .CO(n28632));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n29734), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1200_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n29235), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n29974), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n29734), .I0(n1908), .I1(n1928), .CO(n29735));
    SB_CARRY mod_5_add_2076_24 (.CI(n29974), .I0(n2988), .I1(n3017), .CO(n29975));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n44219), 
            .I3(n29733), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n29973), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_3 (.CI(n29733), .I0(n1909), .I1(n44219), .CO(n29734));
    SB_CARRY mod_5_add_2076_23 (.CI(n29973), .I0(n2989), .I1(n3017), .CO(n29974));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n44219), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1200_add_4_26 (.CI(n29235), .I0(GND_net), .I1(timer[24]), 
            .CO(n29236));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_513[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_c)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n29972), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n44219), 
            .CO(n29733));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n28631));
    SB_LUT4 timer_1200_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n29234), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_22 (.CI(n29972), .I0(n2990), .I1(n3017), .CO(n29973));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n29732), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n29971), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n29731), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n29971), .I0(n2991), .I1(n3017), .CO(n29972));
    SB_CARRY mod_5_add_1272_15 (.CI(n29731), .I0(n1797), .I1(n1829), .CO(n29732));
    SB_CARRY timer_1200_add_4_25 (.CI(n29234), .I0(GND_net), .I1(timer[23]), 
            .CO(n29235));
    SB_LUT4 timer_1200_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n29233), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1200_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n29970), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n29730), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n29970), .I0(n2992), .I1(n3017), .CO(n29971));
    SB_CARRY mod_5_add_1272_14 (.CI(n29730), .I0(n1798), .I1(n1829), .CO(n29731));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n29729), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n29729), .I0(n1799), .I1(n1829), .CO(n29730));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n29969), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n29728), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n29969), .I0(n2993), .I1(n3017), .CO(n29970));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n29968), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n29968), .I0(n2994), .I1(n3017), .CO(n29969));
    SB_CARRY mod_5_add_1272_12 (.CI(n29728), .I0(n1800), .I1(n1829), .CO(n29729));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n29967), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n29967), .I0(n2995), .I1(n3017), .CO(n29968));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n29727), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n29727), .I0(n1801), .I1(n1829), .CO(n29728));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n29726), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1472 (.I0(n1806), .I1(n1804), .I2(n1796), .I3(n1799), 
            .O(n24_adj_4177));
    defparam i10_4_lut_adj_1472.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1473 (.I0(n1807), .I1(n1797), .I2(n1802), .I3(n1808), 
            .O(n22));
    defparam i8_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1474 (.I0(n1803), .I1(n1801), .I2(n1800), .I3(n1805), 
            .O(n23));
    defparam i9_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n29966), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n29726), .I0(n1802), .I1(n1829), .CO(n29727));
    SB_CARRY add_21_7 (.CI(n28431), .I0(bit_ctr[5]), .I1(GND_net), .CO(n28432));
    SB_LUT4 i7_3_lut_adj_1475 (.I0(n1798), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4178));
    defparam i7_3_lut_adj_1475.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_2076_16 (.CI(n29966), .I0(n2996), .I1(n3017), .CO(n29967));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n29725), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n29965), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n29725), .I0(n1803), .I1(n1829), .CO(n29726));
    SB_CARRY mod_5_add_2076_15 (.CI(n29965), .I0(n2997), .I1(n3017), .CO(n29966));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n29724), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut (.I0(n21_adj_4178), .I1(n23), .I2(n22), .I3(n24_adj_4177), 
            .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n29964), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n29724), .I0(n1804), .I1(n1829), .CO(n29725));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n29723), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n29723), .I0(n1805), .I1(n1829), .CO(n29724));
    SB_CARRY mod_5_add_2076_14 (.CI(n29964), .I0(n2998), .I1(n3017), .CO(n29965));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n29722), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n29963), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n28442), .I0(bit_ctr[16]), .I1(GND_net), .CO(n28443));
    SB_CARRY mod_5_add_2076_13 (.CI(n29963), .I0(n2999), .I1(n3017), .CO(n29964));
    SB_CARRY mod_5_add_1272_6 (.CI(n29722), .I0(n1806), .I1(n1829), .CO(n29723));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n29962), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n29962), .I0(n3000), .I1(n3017), .CO(n29963));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n29721), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n29721), .I0(n1807), .I1(n1829), .CO(n29722));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n29961), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1476 (.I0(n2791), .I1(n2795), .I2(n2802), .I3(n2799), 
            .O(n40_adj_4179));
    defparam i16_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_11 (.CI(n29961), .I0(n3001), .I1(n3017), .CO(n29962));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n29720), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1477 (.I0(n2786), .I1(n2801), .I2(n2807), .I3(n2803), 
            .O(n38_adj_4180));
    defparam i14_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n29960), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n29960), .I0(n3002), .I1(n3017), .CO(n29961));
    SB_CARRY mod_5_add_1272_4 (.CI(n29720), .I0(n1808), .I1(n1829), .CO(n29721));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n44221), 
            .I3(n29719), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n29959), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1478 (.I0(n2793), .I1(n2806), .I2(n2794), .I3(n2787), 
            .O(n39_adj_4181));
    defparam i15_4_lut_adj_1478.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1272_3 (.CI(n29719), .I0(n1809), .I1(n44221), .CO(n29720));
    SB_CARRY mod_5_add_2076_9 (.CI(n29959), .I0(n3003), .I1(n3017), .CO(n29960));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n44221), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n44221), 
            .CO(n29719));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n29718), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n29717), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n29717), .I0(n1698), .I1(n1730), .CO(n29718));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n29958), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n29958), .I0(n3004), .I1(n3017), .CO(n29959));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n29716), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n29716), .I0(n1699), .I1(n1730), .CO(n29717));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n29957), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n29957), .I0(n3005), .I1(n3017), .CO(n29958));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n29956), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_6 (.CI(n29956), .I0(n3006), .I1(n3017), .CO(n29957));
    SB_LUT4 i11_4_lut_adj_1479 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26));
    defparam i11_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1480 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4182));
    defparam i4_3_lut_adj_1480.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4183));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n29715), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1481 (.I0(n2796), .I1(n2798), .I2(n2788), .I3(n2800), 
            .O(n37));
    defparam i13_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1482 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4184));
    defparam i9_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1483 (.I0(n19_adj_4182), .I1(n26), .I2(n1905), 
            .I3(n1903), .O(n28));
    defparam i13_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1484 (.I0(n1896), .I1(n28), .I2(n24_adj_4184), 
            .I3(n16_adj_4183), .O(n1928));
    defparam i14_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n29955), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n29955), .I0(n3007), .I1(n3017), .CO(n29956));
    SB_CARRY mod_5_add_1205_12 (.CI(n29715), .I0(n1700), .I1(n1730), .CO(n29716));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n29714), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_3_lut (.I0(bit_ctr[7]), .I1(n2808), .I2(n2809), .I3(GND_net), 
            .O(n36));
    defparam i12_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i11_2_lut (.I0(n2805), .I1(n2804), .I2(GND_net), .I3(GND_net), 
            .O(n35));
    defparam i11_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i22_4_lut_adj_1485 (.I0(n37), .I1(n39_adj_4181), .I2(n38_adj_4180), 
            .I3(n40_adj_4179), .O(n46_adj_4185));
    defparam i22_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n29954), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n29714), .I0(n1701), .I1(n1730), .CO(n29715));
    SB_CARRY mod_5_add_2076_4 (.CI(n29954), .I0(n3008), .I1(n3017), .CO(n29955));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n29713), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(n19), .I1(bit_ctr[15]), .I2(GND_net), .I3(n28441), 
            .O(n41294)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n44220), 
            .I3(n29953), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i17_4_lut (.I0(n2797), .I1(n2789), .I2(n2790), .I3(n2792), 
            .O(n41_adj_4186));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1205_10 (.CI(n29713), .I0(n1702), .I1(n1730), .CO(n29714));
    SB_CARRY mod_5_add_2076_3 (.CI(n29953), .I0(n3009), .I1(n44220), .CO(n29954));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n44220), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n29712), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n29712), .I0(n1703), .I1(n1730), .CO(n29713));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n44220), 
            .CO(n29953));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n29711), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_3_lut (.I0(n2596), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n28_adj_4187));
    defparam i6_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1486 (.I0(n2595), .I1(n2590), .I2(n2592), .I3(n2599), 
            .O(n35_adj_4188));
    defparam i13_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1487 (.I0(n2593), .I1(n2605), .I2(n2589), .I3(n2608), 
            .O(n34));
    defparam i12_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1205_8 (.CI(n29711), .I0(n1704), .I1(n1730), .CO(n29712));
    SB_LUT4 i18_4_lut_adj_1488 (.I0(n35_adj_4188), .I1(n2606), .I2(n28_adj_4187), 
            .I3(n2603), .O(n40_adj_4189));
    defparam i18_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1489 (.I0(n2591), .I1(n2588), .I2(n2594), .I3(n2598), 
            .O(n38_adj_4190));
    defparam i16_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n29710), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_3_lut (.I0(n2602), .I1(n34), .I2(n2607), .I3(GND_net), 
            .O(n39_adj_4191));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1490 (.I0(n2597), .I1(n2600), .I2(n2601), .I3(n2604), 
            .O(n37_adj_4192));
    defparam i15_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1491 (.I0(n37_adj_4192), .I1(n39_adj_4191), .I2(n38_adj_4190), 
            .I3(n40_adj_4189), .O(n2621));
    defparam i21_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_4186), .I1(n46_adj_4185), .I2(n35), 
            .I3(n36), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n29952), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i37378_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44230));
    defparam i37378_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n29951), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n29710), .I0(n1705), .I1(n1730), .CO(n29711));
    SB_CARRY add_21_17 (.CI(n28441), .I0(bit_ctr[15]), .I1(GND_net), .CO(n28442));
    SB_CARRY mod_5_add_2009_26 (.CI(n29951), .I0(n2886), .I1(n2918), .CO(n29952));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n29709), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n29950), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n28430), 
            .O(n41283)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1205_6 (.CI(n29709), .I0(n1706), .I1(n1730), .CO(n29710));
    SB_CARRY mod_5_add_2009_25 (.CI(n29950), .I0(n2887), .I1(n2918), .CO(n29951));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n29708), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n29949), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n29949), .I0(n2888), .I1(n2918), .CO(n29950));
    SB_CARRY mod_5_add_1205_5 (.CI(n29708), .I0(n1707), .I1(n1730), .CO(n29709));
    SB_LUT4 i37367_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44219));
    defparam i37367_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n29948), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n28430), .I0(bit_ctr[4]), .I1(GND_net), .CO(n28431));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n29707), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n29948), .I0(n2889), .I1(n2918), .CO(n29949));
    SB_CARRY mod_5_add_1205_4 (.CI(n29707), .I0(n1708), .I1(n1730), .CO(n29708));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n29947), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n44222), 
            .I3(n29706), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_22 (.CI(n29947), .I0(n2890), .I1(n2918), .CO(n29948));
    SB_CARRY mod_5_add_1205_3 (.CI(n29706), .I0(n1709), .I1(n44222), .CO(n29707));
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n28440), 
            .O(n41293)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_16 (.CI(n28440), .I0(bit_ctr[14]), .I1(GND_net), .CO(n28441));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n29946), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n44222), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_21 (.CI(n29946), .I0(n2891), .I1(n2918), .CO(n29947));
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n44222), 
            .CO(n29706));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n29705), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n29704), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n29945), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n29945), .I0(n2892), .I1(n2918), .CO(n29946));
    SB_CARRY mod_5_add_1138_13 (.CI(n29704), .I0(n1599), .I1(n1631), .CO(n29705));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n29944), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n29703), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n29944), .I0(n2893), .I1(n2918), .CO(n29945));
    SB_CARRY mod_5_add_1138_12 (.CI(n29703), .I0(n1600), .I1(n1631), .CO(n29704));
    SB_LUT4 i37371_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44223));
    defparam i37371_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n29943), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n29702), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n29943), .I0(n2894), .I1(n2918), .CO(n29944));
    SB_CARRY mod_5_add_1138_11 (.CI(n29702), .I0(n1601), .I1(n1631), .CO(n29703));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n29942), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n29701), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n29942), .I0(n2895), .I1(n2918), .CO(n29943));
    SB_CARRY mod_5_add_1138_10 (.CI(n29701), .I0(n1602), .I1(n1631), .CO(n29702));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n29941), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n29700), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n29700), .I0(n1603), .I1(n1631), .CO(n29701));
    SB_CARRY mod_5_add_2009_16 (.CI(n29941), .I0(n2896), .I1(n2918), .CO(n29942));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n29699), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n29940), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n29699), .I0(n1604), .I1(n1631), .CO(n29700));
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n28439), 
            .O(n41292)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n29698), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n29940), .I0(n2897), .I1(n2918), .CO(n29941));
    SB_CARRY mod_5_add_1138_7 (.CI(n29698), .I0(n1605), .I1(n1631), .CO(n29699));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n29939), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n29939), .I0(n2898), .I1(n2918), .CO(n29940));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n29697), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n29938), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n29697), .I0(n1606), .I1(n1631), .CO(n29698));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n29696), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n29696), .I0(n1607), .I1(n1631), .CO(n29697));
    SB_CARRY mod_5_add_2009_13 (.CI(n29938), .I0(n2899), .I1(n2918), .CO(n29939));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n29695), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n29695), .I0(n1608), .I1(n1631), .CO(n29696));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n29937), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n29937), .I0(n2900), .I1(n2918), .CO(n29938));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n44225), 
            .I3(n29694), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n29694), .I0(n1609), .I1(n44225), .CO(n29695));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n29936), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n29936), .I0(n2901), .I1(n2918), .CO(n29937));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n29935), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n44225), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_10 (.CI(n29935), .I0(n2902), .I1(n2918), .CO(n29936));
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n44225), 
            .CO(n29694));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n29934), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n29934), .I0(n2903), .I1(n2918), .CO(n29935));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n29933), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n29933), .I0(n2904), .I1(n2918), .CO(n29934));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n29932), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n29932), .I0(n2905), .I1(n2918), .CO(n29933));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n29931), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n29931), .I0(n2906), .I1(n2918), .CO(n29932));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n29930), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n29930), .I0(n2907), .I1(n2918), .CO(n29931));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n29929), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n29929), .I0(n2908), .I1(n2918), .CO(n29930));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n44223), 
            .I3(n29928), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n29928), .I0(n2909), .I1(n44223), .CO(n29929));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n44223), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n44223), 
            .CO(n29928));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n29927), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n29926), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n29926), .I0(n2787), .I1(n2819), .CO(n29927));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n29925), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(one_wire_N_513[9]), .I1(one_wire_N_513[10]), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'heeee;
    SB_LUT4 i20694_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n25417));
    defparam i20694_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i36628_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n35446));
    defparam i36628_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16_4_lut_adj_1493 (.I0(n21_adj_4194), .I1(n23_adj_4195), .I2(n22_adj_4196), 
            .I3(n24_adj_4197), .O(n36_adj_4198));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1494 (.I0(n25), .I1(n27), .I2(n26_adj_4199), 
            .I3(n28_adj_4200), .O(n37_adj_4201));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37_adj_4201), .I1(n29_adj_4202), .I2(n36_adj_4198), 
            .I3(n30_adj_4203), .O(n15928));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_513[4]), .I1(one_wire_N_513[3]), .I2(n35446), 
            .I3(n30771), .O(n112));
    defparam i1_4_lut.LUT_INIT = 16'h5155;
    SB_LUT4 i1_4_lut_adj_1495 (.I0(n112), .I1(n35446), .I2(one_wire_N_513[2]), 
            .I3(one_wire_N_513[3]), .O(n106));
    defparam i1_4_lut_adj_1495.LUT_INIT = 16'haeee;
    SB_LUT4 i37351_3_lut (.I0(\state[1] ), .I1(n35266), .I2(n15928), .I3(GND_net), 
            .O(n38137));
    defparam i37351_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i37366_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44218));
    defparam i37366_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_24 (.CI(n29925), .I0(n2788), .I1(n2819), .CO(n29926));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n29924), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n29924), .I0(n2789), .I1(n2819), .CO(n29925));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n29923), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20840_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n25569));
    defparam i20840_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1942_22 (.CI(n29923), .I0(n2790), .I1(n2819), .CO(n29924));
    SB_LUT4 i6_4_lut (.I0(n1405), .I1(n25569), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4204));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1496 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4205));
    defparam i7_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1497 (.I0(n17_adj_4205), .I1(n1408), .I2(n16_adj_4204), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n29922), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n29922), .I0(n2791), .I1(n2819), .CO(n29923));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n29921), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n29921), .I0(n2792), .I1(n2819), .CO(n29922));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n29920), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_2_lut_adj_1498 (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4206));
    defparam i5_2_lut_adj_1498.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1499 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4207));
    defparam i15_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_15 (.CI(n28439), .I0(bit_ctr[13]), .I1(GND_net), .CO(n28440));
    SB_LUT4 i20937_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n25667));
    defparam i20937_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1500 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n25667), 
            .O(n36_adj_4208));
    defparam i13_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n28438), 
            .O(n41291)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_19 (.CI(n29920), .I0(n2793), .I1(n2819), .CO(n29921));
    SB_LUT4 i19_4_lut_adj_1501 (.I0(n2700), .I1(n38_adj_4207), .I2(n28_adj_4206), 
            .I3(n2705), .O(n42));
    defparam i19_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n29919), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n29919), .I0(n2794), .I1(n2819), .CO(n29920));
    SB_LUT4 i17_4_lut_adj_1502 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4209));
    defparam i17_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1503 (.I0(n2687), .I1(n36_adj_4208), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4210));
    defparam i18_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1504 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4211));
    defparam i16_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1505 (.I0(n39_adj_4211), .I1(n41_adj_4210), .I2(n40_adj_4209), 
            .I3(n42), .O(n2720));
    defparam i22_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n28511), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n29918), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n28510), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n28429), 
            .O(n41282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_14 (.CI(n28438), .I0(bit_ctr[12]), .I1(GND_net), .CO(n28439));
    SB_CARRY mod_5_add_1942_17 (.CI(n29918), .I0(n2795), .I1(n2819), .CO(n29919));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n29917), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(n19), .I1(bit_ctr[11]), .I2(GND_net), .I3(n28437), 
            .O(n41290)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_5 (.CI(n28429), .I0(bit_ctr[3]), .I1(GND_net), .CO(n28430));
    SB_CARRY mod_5_add_1942_16 (.CI(n29917), .I0(n2796), .I1(n2819), .CO(n29918));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n29916), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n29916), .I0(n2797), .I1(n2819), .CO(n29917));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n29915), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n29915), .I0(n2798), .I1(n2819), .CO(n29916));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n29914), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n29914), .I0(n2799), .I1(n2819), .CO(n29915));
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n25553), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hd622;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n29913), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n29913), .I0(n2800), .I1(n2819), .CO(n29914));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n29912), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n29912), .I0(n2801), .I1(n2819), .CO(n29913));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n29911), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n29911), .I0(n2802), .I1(n2819), .CO(n29912));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n29910), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n28510), .I0(n1500), .I1(n1532), .CO(n28511));
    SB_CARRY mod_5_add_1942_9 (.CI(n29910), .I0(n2803), .I1(n2819), .CO(n29911));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n29909), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n29909), .I0(n2804), .I1(n2819), .CO(n29910));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n28509), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n29908), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n28509), .I0(n1501), .I1(n1532), .CO(n28510));
    SB_LUT4 i37375_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44227));
    defparam i37375_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n28508), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1200__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY add_21_13 (.CI(n28437), .I0(bit_ctr[11]), .I1(GND_net), .CO(n28438));
    SB_CARRY mod_5_add_1071_10 (.CI(n28508), .I0(n1502), .I1(n1532), .CO(n28509));
    SB_CARRY mod_5_add_1942_7 (.CI(n29908), .I0(n2805), .I1(n2819), .CO(n29909));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n29907), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i37373_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44225));
    defparam i37373_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_6 (.CI(n29907), .I0(n2806), .I1(n2819), .CO(n29908));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n29906), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n29906), .I0(n2807), .I1(n2819), .CO(n29907));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n28507), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n28428), 
            .O(n41281)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n29905), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n29905), .I0(n2808), .I1(n2819), .CO(n29906));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n44227), 
            .I3(n29904), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n29904), .I0(n2809), .I1(n44227), .CO(n29905));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n44227), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1071_9 (.CI(n28507), .I0(n1503), .I1(n1532), .CO(n28508));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n44227), 
            .CO(n29904));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n29903), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n28506), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28606), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut_adj_1506 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4212));
    defparam i8_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), .I3(GND_net), 
            .O(n13));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4213));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n29902), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1507 (.I0(n13), .I1(n20_adj_4212), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4214));
    defparam i10_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_24 (.CI(n29902), .I0(n2688), .I1(n2720), .CO(n29903));
    SB_LUT4 i11_4_lut_adj_1508 (.I0(n1601), .I1(n22_adj_4214), .I2(n18_adj_4213), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n29901), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n29901), .I0(n2689), .I1(n2720), .CO(n29902));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n29900), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n29900), .I0(n2690), .I1(n2720), .CO(n29901));
    SB_CARRY mod_5_add_1071_8 (.CI(n28506), .I0(n1504), .I1(n1532), .CO(n28507));
    SB_LUT4 i37370_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44222));
    defparam i37370_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_12_lut (.I0(n19), .I1(bit_ctr[10]), .I2(GND_net), .I3(n28436), 
            .O(n41289)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n29899), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n29899), .I0(n2691), .I1(n2720), .CO(n29900));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n29898), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n29898), .I0(n2692), .I1(n2720), .CO(n29899));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28605), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n29897), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n29897), .I0(n2693), .I1(n2720), .CO(n29898));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n29896), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28605), .I0(n1401), .I1(n1433), .CO(n28606));
    SB_CARRY add_21_4 (.CI(n28428), .I0(bit_ctr[2]), .I1(GND_net), .CO(n28429));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n28505), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n29896), .I0(n2694), .I1(n2720), .CO(n29897));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n29895), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28604), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n28604), .I0(n1402), .I1(n1433), .CO(n28605));
    SB_CARRY mod_5_add_1071_7 (.CI(n28505), .I0(n1505), .I1(n1532), .CO(n28506));
    SB_CARRY mod_5_add_1875_17 (.CI(n29895), .I0(n2695), .I1(n2720), .CO(n29896));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n29894), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n29894), .I0(n2696), .I1(n2720), .CO(n29895));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n29893), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n29893), .I0(n2697), .I1(n2720), .CO(n29894));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n29892), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n29892), .I0(n2698), .I1(n2720), .CO(n29893));
    SB_CARRY add_21_12 (.CI(n28436), .I0(bit_ctr[10]), .I1(GND_net), .CO(n28437));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n29891), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n29891), .I0(n2699), .I1(n2720), .CO(n29892));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n29890), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n29890), .I0(n2700), .I1(n2720), .CO(n29891));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28603), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n29889), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n28504), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n29889), .I0(n2701), .I1(n2720), .CO(n29890));
    SB_CARRY mod_5_add_1004_9 (.CI(n28603), .I0(n1403), .I1(n1433), .CO(n28604));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n29888), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n29888), .I0(n2702), .I1(n2720), .CO(n29889));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n29887), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n29887), .I0(n2703), .I1(n2720), .CO(n29888));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n29886), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28602), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n28602), .I0(n1404), .I1(n1433), .CO(n28603));
    SB_CARRY mod_5_add_1875_8 (.CI(n29886), .I0(n2704), .I1(n2720), .CO(n29887));
    SB_CARRY mod_5_add_1071_6 (.CI(n28504), .I0(n1506), .I1(n1532), .CO(n28505));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n29885), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n29885), .I0(n2705), .I1(n2720), .CO(n29886));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n29884), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n29884), .I0(n2706), .I1(n2720), .CO(n29885));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n29883), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28601), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n28503), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n28503), .I0(n1507), .I1(n1532), .CO(n28504));
    SB_CARRY mod_5_add_1875_5 (.CI(n29883), .I0(n2707), .I1(n2720), .CO(n29884));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n29882), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n28502), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n28502), .I0(n1508), .I1(n1532), .CO(n28503));
    SB_LUT4 add_21_11_lut (.I0(n19), .I1(bit_ctr[9]), .I2(GND_net), .I3(n28435), 
            .O(n41288)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_4 (.CI(n29882), .I0(n2708), .I1(n2720), .CO(n29883));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n44230), 
            .I3(n29881), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n29881), .I0(n2709), .I1(n44230), .CO(n29882));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n44230), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n44230), 
            .CO(n29881));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n29880), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n29879), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n29879), .I0(n2589), .I1(n2621), .CO(n29880));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n29878), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n29878), .I0(n2590), .I1(n2621), .CO(n29879));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n29877), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n29877), .I0(n2591), .I1(n2621), .CO(n29878));
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n34088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17620));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17619));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17618));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17617));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17616));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17615));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17614));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17613));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17612));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17611));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17610));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17609));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17608));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n29876), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n28601), .I0(n1405), .I1(n1433), .CO(n28602));
    SB_CARRY mod_5_add_1808_20 (.CI(n29876), .I0(n2592), .I1(n2621), .CO(n29877));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n29875), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n29875), .I0(n2593), .I1(n2621), .CO(n29876));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n44229), 
            .I3(n28501), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n29874), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n29874), .I0(n2594), .I1(n2621), .CO(n29875));
    SB_LUT4 add_21_3_lut (.I0(n19), .I1(bit_ctr[1]), .I2(GND_net), .I3(n28427), 
            .O(n41280)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_11 (.CI(n28435), .I0(bit_ctr[9]), .I1(GND_net), .CO(n28436));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n29873), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n29873), .I0(n2595), .I1(n2621), .CO(n29874));
    SB_CARRY mod_5_add_1071_3 (.CI(n28501), .I0(n1509), .I1(n44229), .CO(n28502));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n29872), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n29872), .I0(n2596), .I1(n2621), .CO(n29873));
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n17075), .D(\neo_pixel_transmitter.done_N_576 ), 
            .R(n36850));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n29871), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n44229), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_15 (.CI(n29871), .I0(n2597), .I1(n2621), .CO(n29872));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n29870), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n29870), .I0(n2598), .I1(n2621), .CO(n29871));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n29869), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n29869), .I0(n2599), .I1(n2621), .CO(n29870));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n29868), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n29868), .I0(n2600), .I1(n2621), .CO(n29869));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n29867), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28600), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n29867), .I0(n2601), .I1(n2621), .CO(n29868));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n29866), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n29866), .I0(n2602), .I1(n2621), .CO(n29867));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n29865), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n29865), .I0(n2603), .I1(n2621), .CO(n29866));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n29864), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n29864), .I0(n2604), .I1(n2621), .CO(n29865));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n29863), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28600), .I0(n1406), .I1(n1433), .CO(n28601));
    SB_CARRY mod_5_add_1808_7 (.CI(n29863), .I0(n2605), .I1(n2621), .CO(n29864));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28599), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n29862), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n28599), .I0(n1407), .I1(n1433), .CO(n28600));
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n44229), 
            .CO(n28501));
    SB_CARRY mod_5_add_1808_6 (.CI(n29862), .I0(n2606), .I1(n2621), .CO(n29863));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28598), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n29861), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n29861), .I0(n2607), .I1(n2621), .CO(n29862));
    SB_CARRY mod_5_add_1004_4 (.CI(n28598), .I0(n1408), .I1(n1433), .CO(n28599));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_513[22]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n28661), .O(n22_adj_4196)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n28457), 
            .O(n41274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_513[17]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n28660), .O(n24_adj_4197)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n29860), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_32 (.CI(n28660), .I0(timer[30]), .I1(n1[30]), 
            .CO(n28661));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_513[12]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n28659), .O(n26_adj_4199)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_4 (.CI(n29860), .I0(n2608), .I1(n2621), .CO(n29861));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n44231), 
            .I3(n28597), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n28597), .I0(n1409), .I1(n44231), .CO(n28598));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n44232), 
            .I3(n29859), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n44231), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n28456), 
            .O(n41273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_31 (.CI(n28659), .I0(timer[29]), .I1(n1[29]), 
            .CO(n28660));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n44231), 
            .CO(n28597));
    SB_CARRY mod_5_add_1808_3 (.CI(n29859), .I0(n2609), .I1(n44232), .CO(n29860));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n44232), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n44232), 
            .CO(n29859));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_513[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n28658), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n28658), .I0(timer[28]), .I1(n1[28]), 
            .CO(n28659));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n29858), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n29857), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n29857), .I0(n2490), .I1(n2522), .CO(n29858));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n29856), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_513[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n28657), .O(n21_adj_4194)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n28657), .I0(timer[27]), .I1(n1[27]), 
            .CO(n28658));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n28656), .O(one_wire_N_513[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n29856), .I0(n2491), .I1(n2522), .CO(n29857));
    SB_CARRY sub_14_add_2_28 (.CI(n28656), .I0(timer[26]), .I1(n1[26]), 
            .CO(n28657));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n29855), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_27_lut (.I0(one_wire_N_513[13]), .I1(timer[25]), 
            .I2(n1[25]), .I3(n28655), .O(n23_adj_4195)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n28655), .I0(timer[25]), .I1(n1[25]), 
            .CO(n28656));
    SB_LUT4 sub_14_add_2_26_lut (.I0(one_wire_N_513[19]), .I1(timer[24]), 
            .I2(n1[24]), .I3(n28654), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_20 (.CI(n29855), .I0(n2492), .I1(n2522), .CO(n29856));
    SB_CARRY sub_14_add_2_26 (.CI(n28654), .I0(timer[24]), .I1(n1[24]), 
            .CO(n28655));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n29854), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_513[20]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n28653), .O(n30_adj_4203)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n28653), .I0(timer[23]), .I1(n1[23]), 
            .CO(n28654));
    SB_CARRY mod_5_add_1741_19 (.CI(n29854), .I0(n2493), .I1(n2522), .CO(n29855));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n29853), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n29853), .I0(n2494), .I1(n2522), .CO(n29854));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n29852), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n28652), .O(one_wire_N_513[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_17 (.CI(n29852), .I0(n2495), .I1(n2522), .CO(n29853));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n29851), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n29851), .I0(n2496), .I1(n2522), .CO(n29852));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n29850), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_24 (.CI(n28652), .I0(timer[22]), .I1(n1[22]), 
            .CO(n28653));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_513[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n28651), .O(n28_adj_4200)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_15 (.CI(n29850), .I0(n2497), .I1(n2522), .CO(n29851));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n29849), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_23 (.CI(n28651), .I0(timer[21]), .I1(n1[21]), 
            .CO(n28652));
    SB_CARRY mod_5_add_1741_14 (.CI(n29849), .I0(n2498), .I1(n2522), .CO(n29850));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n29848), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n29848), .I0(n2499), .I1(n2522), .CO(n29849));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n29847), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n29847), .I0(n2500), .I1(n2522), .CO(n29848));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n29846), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n29846), .I0(n2501), .I1(n2522), .CO(n29847));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n29845), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n29845), .I0(n2502), .I1(n2522), .CO(n29846));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n29844), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n29844), .I0(n2503), .I1(n2522), .CO(n29845));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n29843), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n29843), .I0(n2504), .I1(n2522), .CO(n29844));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n29842), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n29842), .I0(n2505), .I1(n2522), .CO(n29843));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n29841), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_22_lut (.I0(GND_net), .I1(timer[20]), .I2(n1[20]), 
            .I3(n28650), .O(one_wire_N_513[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n29841), .I0(n2506), .I1(n2522), .CO(n29842));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n29840), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n29840), .I0(n2507), .I1(n2522), .CO(n29841));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n29839), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n28650), .I0(timer[20]), .I1(n1[20]), 
            .CO(n28651));
    SB_LUT4 i20921_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n25651));
    defparam i20921_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1509 (.I0(n2004), .I1(n1998), .I2(n2006), .I3(n2002), 
            .O(n28_adj_4217));
    defparam i12_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1510 (.I0(n1995), .I1(n2003), .I2(n2007), .I3(n25651), 
            .O(n26_adj_4218));
    defparam i10_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1511 (.I0(n1994), .I1(n2005), .I2(n1996), .I3(n1997), 
            .O(n27_adj_4219));
    defparam i11_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1512 (.I0(n2008), .I1(n2000), .I2(n1999), .I3(n2001), 
            .O(n25_adj_4220));
    defparam i9_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1513 (.I0(n25_adj_4220), .I1(n27_adj_4219), .I2(n26_adj_4218), 
            .I3(n28_adj_4217), .O(n2027));
    defparam i15_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_2_lut (.I0(n3088), .I1(n3108), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_4221));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1514 (.I0(n3086), .I1(n3094), .I2(n3093), .I3(n3085), 
            .O(n46_adj_4222));
    defparam i19_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1515 (.I0(n3102), .I1(n3084), .I2(n3091), .I3(n3106), 
            .O(n42_adj_4223));
    defparam i15_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut_adj_1516 (.I0(n3099), .I1(bit_ctr[4]), .I2(n3109), 
            .I3(GND_net), .O(n33_adj_4224));
    defparam i6_3_lut_adj_1516.LUT_INIT = 16'heaea;
    SB_LUT4 i16_4_lut_adj_1517 (.I0(n3104), .I1(n3083), .I2(n3092), .I3(n3101), 
            .O(n43_adj_4225));
    defparam i16_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1518 (.I0(n3103), .I1(n46_adj_4222), .I2(n36_adj_4221), 
            .I3(n3087), .O(n50));
    defparam i23_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1519 (.I0(n3097), .I1(n42_adj_4223), .I2(n3100), 
            .I3(n3089), .O(n48));
    defparam i21_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1520 (.I0(n43_adj_4225), .I1(n33_adj_4224), .I2(n3098), 
            .I3(n3095), .O(n49));
    defparam i22_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n3107), .I1(n3090), .I2(n3105), .I3(n3096), 
            .O(n47_adj_4226));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17607));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_4 (.CI(n29839), .I0(n2508), .I1(n2522), .CO(n29840));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n44234), 
            .I3(n29838), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_10_lut (.I0(n19), .I1(bit_ctr[8]), .I2(GND_net), .I3(n28434), 
            .O(n41287)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n28649), .O(one_wire_N_513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n29838), .I0(n2509), .I1(n44234), .CO(n29839));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n44234), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_32 (.CI(n28456), .I0(bit_ctr[30]), .I1(GND_net), .CO(n28457));
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n44234), 
            .CO(n29838));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n29837), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17606));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17605));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n29836), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n28427), .I0(bit_ctr[1]), .I1(GND_net), .CO(n28428));
    SB_CARRY mod_5_add_1674_21 (.CI(n29836), .I0(n2391), .I1(n2423), .CO(n29837));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n29835), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n29835), .I0(n2392), .I1(n2423), .CO(n29836));
    SB_CARRY sub_14_add_2_21 (.CI(n28649), .I0(timer[19]), .I1(n1[19]), 
            .CO(n28650));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n29834), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n29834), .I0(n2393), .I1(n2423), .CO(n29835));
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17604));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n28867), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28866), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n29833), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n29833), .I0(n2394), .I1(n2423), .CO(n29834));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n29832), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_6 (.CI(n28866), .I0(n906), .I1(VCC_net), .CO(n28867));
    SB_CARRY mod_5_add_1674_17 (.CI(n29832), .I0(n2395), .I1(n2423), .CO(n29833));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n29831), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_10 (.CI(n28434), .I0(bit_ctr[8]), .I1(GND_net), .CO(n28435));
    SB_CARRY mod_5_add_1674_16 (.CI(n29831), .I0(n2396), .I1(n2423), .CO(n29832));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n29830), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n36288), .I2(VCC_net), 
            .I3(n28865), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_15 (.CI(n29830), .I0(n2397), .I1(n2423), .CO(n29831));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n29829), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n29829), .I0(n2398), .I1(n2423), .CO(n29830));
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17603));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_669_5 (.CI(n28865), .I0(n36288), .I1(VCC_net), 
            .CO(n28866));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17229), .I2(VCC_net), 
            .I3(n28864), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n28648), .O(one_wire_N_513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n29828), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n29828), .I0(n2399), .I1(n2423), .CO(n29829));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n29827), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_31_lut (.I0(n11), .I1(bit_ctr[29]), .I2(GND_net), .I3(n28455), 
            .O(n41266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_12 (.CI(n29827), .I0(n2400), .I1(n2423), .CO(n29828));
    SB_CARRY mod_5_add_669_4 (.CI(n28864), .I0(n17229), .I1(VCC_net), 
            .CO(n28865));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n29826), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n29826), .I0(n2401), .I1(n2423), .CO(n29827));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n29825), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n28433), 
            .O(n41286)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_10 (.CI(n29825), .I0(n2402), .I1(n2423), .CO(n29826));
    SB_CARRY add_21_31 (.CI(n28455), .I0(bit_ctr[29]), .I1(GND_net), .CO(n28456));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14415), .I2(GND_net), 
            .I3(n28863), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n29824), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(n11), .I1(bit_ctr[28]), .I2(GND_net), .I3(n28454), 
            .O(n41267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_9 (.CI(n28433), .I0(bit_ctr[7]), .I1(GND_net), .CO(n28434));
    SB_CARRY mod_5_add_669_3 (.CI(n28863), .I0(n14415), .I1(GND_net), 
            .CO(n28864));
    SB_CARRY mod_5_add_1674_9 (.CI(n29824), .I0(n2403), .I1(n2423), .CO(n29825));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n29823), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n29823), .I0(n2404), .I1(n2423), .CO(n29824));
    SB_DFF timer_1200__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17058), .D(state_3__N_362[0]), 
            .S(n17312));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n29822), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_20 (.CI(n28648), .I0(timer[18]), .I1(n1[18]), 
            .CO(n28649));
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28863));
    SB_CARRY mod_5_add_1674_7 (.CI(n29822), .I0(n2405), .I1(n2423), .CO(n29823));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n29821), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n29821), .I0(n2406), .I1(n2423), .CO(n29822));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n29820), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1200__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4228), .I1(n4_adj_4228), .I2(n1037), 
            .I3(n28862), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n29820), .I0(n2407), .I1(n2423), .CO(n29821));
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28861), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n29819), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28861), .I0(n1005), .I1(n1037), .CO(n28862));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28860), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n29819), .I0(n2408), .I1(n2423), .CO(n29820));
    SB_CARRY mod_5_add_736_6 (.CI(n28860), .I0(n1006), .I1(n1037), .CO(n28861));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n44235), 
            .I3(n29818), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n29818), .I0(n2409), .I1(n44235), .CO(n29819));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n44235), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n1[17]), 
            .I3(n28647), .O(one_wire_N_513[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n28454), .I0(bit_ctr[28]), .I1(GND_net), .CO(n28455));
    SB_LUT4 add_21_29_lut (.I0(n19), .I1(bit_ctr[27]), .I2(GND_net), .I3(n28453), 
            .O(n41271)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n44235), 
            .CO(n29818));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28859), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28859), .I0(n1007), .I1(n1037), .CO(n28860));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28858), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n28858), .I0(n1008), .I1(n1037), .CO(n28859));
    SB_CARRY add_21_29 (.CI(n28453), .I0(bit_ctr[27]), .I1(GND_net), .CO(n28454));
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n41272)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n28432), 
            .O(n41285)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_DFF timer_1200__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1200__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n34150));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17389));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17602));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17601));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17600));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17599));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17598));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17597));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17596));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17595));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17594));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17592));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17591));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17578));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n44236), 
            .I3(n28857), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n28857), .I0(n1009), .I1(n44236), .CO(n28858));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n44236), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n44236), 
            .CO(n28857));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n29817), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n29816), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n29816), .I0(n2292), .I1(n2324), .CO(n29817));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n29815), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n29815), .I0(n2293), .I1(n2324), .CO(n29816));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n29814), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n29814), .I0(n2294), .I1(n2324), .CO(n29815));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n29813), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n29813), .I0(n2295), .I1(n2324), .CO(n29814));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n29812), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n29812), .I0(n2296), .I1(n2324), .CO(n29813));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n29811), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n29811), .I0(n2297), .I1(n2324), .CO(n29812));
    SB_LUT4 add_21_28_lut (.I0(n19), .I1(bit_ctr[26]), .I2(GND_net), .I3(n28452), 
            .O(n41279)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n29810), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n29810), .I0(n2298), .I1(n2324), .CO(n29811));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n29809), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n29809), .I0(n2299), .I1(n2324), .CO(n29810));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n29808), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n29808), .I0(n2300), .I1(n2324), .CO(n29809));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n29807), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n29807), .I0(n2301), .I1(n2324), .CO(n29808));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n29806), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n29806), .I0(n2302), .I1(n2324), .CO(n29807));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n29805), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n28647), .I0(timer[17]), .I1(n1[17]), 
            .CO(n28648));
    SB_CARRY add_21_28 (.CI(n28452), .I0(bit_ctr[26]), .I1(GND_net), .CO(n28453));
    SB_LUT4 sub_14_add_2_18_lut (.I0(one_wire_N_513[15]), .I1(timer[16]), 
            .I2(n1[16]), .I3(n28646), .O(n29_adj_4202)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n28646), .I0(timer[16]), .I1(n1[16]), 
            .CO(n28647));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n28427));
    SB_CARRY mod_5_add_1607_9 (.CI(n29805), .I0(n2303), .I1(n2324), .CO(n29806));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n28645), .O(one_wire_N_513[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n29804), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n29804), .I0(n2304), .I1(n2324), .CO(n29805));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n29803), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n29803), .I0(n2305), .I1(n2324), .CO(n29804));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n29802), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n29802), .I0(n2306), .I1(n2324), .CO(n29803));
    SB_LUT4 add_21_27_lut (.I0(n19), .I1(bit_ctr[25]), .I2(GND_net), .I3(n28451), 
            .O(n41278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n29801), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n29801), .I0(n2307), .I1(n2324), .CO(n29802));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n29800), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n29800), .I0(n2308), .I1(n2324), .CO(n29801));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n44237), 
            .I3(n29799), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n29799), .I0(n2309), .I1(n44237), .CO(n29800));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n44237), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n44237), 
            .CO(n29799));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n29798), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n29797), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n29797), .I0(n2193), .I1(n2225), .CO(n29798));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n29796), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n29796), .I0(n2194), .I1(n2225), .CO(n29797));
    SB_CARRY sub_14_add_2_17 (.CI(n28645), .I0(timer[15]), .I1(n1[15]), 
            .CO(n28646));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n29795), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28807), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28806), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n29795), .I0(n2195), .I1(n2225), .CO(n29796));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n28644), .O(one_wire_N_513[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n29794), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28806), .I0(n1104), .I1(n1136), .CO(n28807));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28805), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28805), .I0(n1105), .I1(n1136), .CO(n28806));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28804), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n29794), .I0(n2196), .I1(n2225), .CO(n29795));
    SB_CARRY mod_5_add_803_6 (.CI(n28804), .I0(n1106), .I1(n1136), .CO(n28805));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28803), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28803), .I0(n1107), .I1(n1136), .CO(n28804));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n29793), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28802), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_16 (.CI(n28644), .I0(timer[14]), .I1(n1[14]), 
            .CO(n28645));
    SB_CARRY mod_5_add_803_4 (.CI(n28802), .I0(n1108), .I1(n1136), .CO(n28803));
    SB_CARRY mod_5_add_1540_15 (.CI(n29793), .I0(n2197), .I1(n2225), .CO(n29794));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n44239), 
            .I3(n28801), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n28801), .I0(n1109), .I1(n44239), .CO(n28802));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n44239), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n44239), 
            .CO(n28801));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n29792), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n29792), .I0(n2198), .I1(n2225), .CO(n29793));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n29791), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n28643), .O(one_wire_N_513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_13 (.CI(n29791), .I0(n2199), .I1(n2225), .CO(n29792));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n29790), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n29790), .I0(n2200), .I1(n2225), .CO(n29791));
    SB_CARRY sub_14_add_2_15 (.CI(n28643), .I0(timer[13]), .I1(n1[13]), 
            .CO(n28644));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n29789), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n29789), .I0(n2201), .I1(n2225), .CO(n29790));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n29788), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n29788), .I0(n2202), .I1(n2225), .CO(n29789));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n29787), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28792), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28791), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28791), .I0(n1203), .I1(n1235), .CO(n28792));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28790), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28790), .I0(n1204), .I1(n1235), .CO(n28791));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28789), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28789), .I0(n1205), .I1(n1235), .CO(n28790));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28788), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n29787), .I0(n2203), .I1(n2225), .CO(n29788));
    SB_CARRY mod_5_add_870_6 (.CI(n28788), .I0(n1206), .I1(n1235), .CO(n28789));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28787), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n29786), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n29786), .I0(n2204), .I1(n2225), .CO(n29787));
    SB_CARRY mod_5_add_870_5 (.CI(n28787), .I0(n1207), .I1(n1235), .CO(n28788));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n28642), .O(one_wire_N_513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n29785), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28786), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n28786), .I0(n1208), .I1(n1235), .CO(n28787));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n44240), 
            .I3(n28785), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_7 (.CI(n29785), .I0(n2205), .I1(n2225), .CO(n29786));
    SB_CARRY mod_5_add_870_3 (.CI(n28785), .I0(n1209), .I1(n44240), .CO(n28786));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n44240), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n29784), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n44240), 
            .CO(n28785));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28784), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28783), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28783), .I0(n1302), .I1(n1334), .CO(n28784));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28782), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28782), .I0(n1303), .I1(n1334), .CO(n28783));
    SB_CARRY mod_5_add_1540_6 (.CI(n29784), .I0(n2206), .I1(n2225), .CO(n29785));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n29783), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28781), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_27 (.CI(n28451), .I0(bit_ctr[25]), .I1(GND_net), .CO(n28452));
    SB_CARRY mod_5_add_937_8 (.CI(n28781), .I0(n1304), .I1(n1334), .CO(n28782));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28780), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n28780), .I0(n1305), .I1(n1334), .CO(n28781));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28779), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28779), .I0(n1306), .I1(n1334), .CO(n28780));
    SB_CARRY mod_5_add_1540_5 (.CI(n29783), .I0(n2207), .I1(n2225), .CO(n29784));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28778), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28778), .I0(n1307), .I1(n1334), .CO(n28779));
    SB_LUT4 add_21_26_lut (.I0(n19), .I1(bit_ctr[24]), .I2(GND_net), .I3(n28450), 
            .O(n41277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28777), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_26 (.CI(n28450), .I0(bit_ctr[24]), .I1(GND_net), .CO(n28451));
    SB_CARRY mod_5_add_937_4 (.CI(n28777), .I0(n1308), .I1(n1334), .CO(n28778));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n44241), 
            .I3(n28776), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n28776), .I0(n1309), .I1(n44241), .CO(n28777));
    SB_LUT4 add_21_25_lut (.I0(n19), .I1(bit_ctr[23]), .I2(GND_net), .I3(n28449), 
            .O(n41276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n44241), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n44241), 
            .CO(n28776));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n29782), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n29782), .I0(n2208), .I1(n2225), .CO(n29783));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n44238), 
            .I3(n29781), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n29781), .I0(n2209), .I1(n44238), .CO(n29782));
    SB_CARRY sub_14_add_2_14 (.CI(n28642), .I0(timer[12]), .I1(n1[12]), 
            .CO(n28643));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n28641), .O(\one_wire_N_513[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n44238), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n44238), 
            .CO(n29781));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n29780), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n29779), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n29779), .I0(n2094), .I1(n2126), .CO(n29780));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n29778), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n29778), .I0(n2095), .I1(n2126), .CO(n29779));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n29777), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n29777), .I0(n2096), .I1(n2126), .CO(n29778));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n29776), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n29776), .I0(n2097), .I1(n2126), .CO(n29777));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n29775), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n29775), .I0(n2098), .I1(n2126), .CO(n29776));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n29774), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n29774), .I0(n2099), .I1(n2126), .CO(n29775));
    SB_CARRY add_21_25 (.CI(n28449), .I0(bit_ctr[23]), .I1(GND_net), .CO(n28450));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n29773), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n29773), .I0(n2100), .I1(n2126), .CO(n29774));
    SB_CARRY sub_14_add_2_13 (.CI(n28641), .I0(timer[11]), .I1(n1[11]), 
            .CO(n28642));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n29772), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n29772), .I0(n2101), .I1(n2126), .CO(n29773));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n28640), .O(one_wire_N_513[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n28640), .I0(timer[10]), .I1(n1[10]), 
            .CO(n28641));
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n28448), 
            .O(n41275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n28639), .O(one_wire_N_513[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n28639), .I0(timer[9]), .I1(n1[9]), 
            .CO(n28640));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n28638), .O(\one_wire_N_513[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n29771), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n28638), .I0(timer[8]), .I1(n1[8]), 
            .CO(n28639));
    SB_CARRY add_21_8 (.CI(n28432), .I0(bit_ctr[6]), .I1(GND_net), .CO(n28433));
    SB_CARRY add_21_24 (.CI(n28448), .I0(bit_ctr[22]), .I1(GND_net), .CO(n28449));
    SB_CARRY mod_5_add_1473_10 (.CI(n29771), .I0(n2102), .I1(n2126), .CO(n29772));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n29770), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n29770), .I0(n2103), .I1(n2126), .CO(n29771));
    SB_LUT4 add_21_23_lut (.I0(n11), .I1(bit_ctr[21]), .I2(GND_net), .I3(n28447), 
            .O(n41270)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n29769), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n29769), .I0(n2104), .I1(n2126), .CO(n29770));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n30005), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n29768), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n29768), .I0(n2105), .I1(n2126), .CO(n29769));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n28637), .O(\one_wire_N_513[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n28447), .I0(bit_ctr[21]), .I1(GND_net), .CO(n28448));
    SB_CARRY sub_14_add_2_9 (.CI(n28637), .I0(timer[7]), .I1(n1[7]), .CO(n28638));
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n30004), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n29767), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n28636), .O(\one_wire_N_513[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_6 (.CI(n29767), .I0(n2106), .I1(n2126), .CO(n29768));
    SB_CARRY mod_5_add_2143_28 (.CI(n30004), .I0(n3084), .I1(n3116), .CO(n30005));
    SB_CARRY sub_14_add_2_8 (.CI(n28636), .I0(timer[6]), .I1(n1[6]), .CO(n28637));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n30003), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n29766), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n29766), .I0(n2107), .I1(n2126), .CO(n29767));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n28635), .O(\one_wire_N_513[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n30003), .I0(n3085), .I1(n3116), .CO(n30004));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n29765), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n29765), .I0(n2108), .I1(n2126), .CO(n29766));
    SB_LUT4 add_21_22_lut (.I0(n11), .I1(bit_ctr[20]), .I2(GND_net), .I3(n28446), 
            .O(n41269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n30002), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n44242), 
            .I3(n29764), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_26 (.CI(n30002), .I0(n3086), .I1(n3116), .CO(n30003));
    SB_CARRY add_21_22 (.CI(n28446), .I0(bit_ctr[20]), .I1(GND_net), .CO(n28447));
    SB_CARRY mod_5_add_1473_3 (.CI(n29764), .I0(n2109), .I1(n44242), .CO(n29765));
    SB_CARRY sub_14_add_2_7 (.CI(n28635), .I0(timer[5]), .I1(n1[5]), .CO(n28636));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n30001), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n44242), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_25 (.CI(n30001), .I0(n3087), .I1(n3116), .CO(n30002));
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n44242), 
            .CO(n29764));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n30000), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n29763), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n30000), .I0(n3088), .I1(n3116), .CO(n30001));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n29762), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n29762), .I0(n1995), .I1(n2027), .CO(n29763));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n29761), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(n11), .I1(bit_ctr[19]), .I2(GND_net), .I3(n28445), 
            .O(n41268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n29999), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n29999), .I0(n3089), .I1(n3116), .CO(n30000));
    SB_CARRY mod_5_add_1406_16 (.CI(n29761), .I0(n1996), .I1(n2027), .CO(n29762));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n29760), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n29760), .I0(n1997), .I1(n2027), .CO(n29761));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n29759), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_21 (.CI(n28445), .I0(bit_ctr[19]), .I1(GND_net), .CO(n28446));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n29998), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n29759), .I0(n1998), .I1(n2027), .CO(n29760));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n29758), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n28634), .O(one_wire_N_513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n29998), .I0(n3090), .I1(n3116), .CO(n29999));
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n28444), 
            .O(n41297)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1406_13 (.CI(n29758), .I0(n1999), .I1(n2027), .CO(n29759));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n29997), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n29997), .I0(n3091), .I1(n3116), .CO(n29998));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n29757), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n29996), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n29757), .I0(n2000), .I1(n2027), .CO(n29758));
    SB_CARRY mod_5_add_2143_20 (.CI(n29996), .I0(n3092), .I1(n3116), .CO(n29997));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n29995), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n29995), .I0(n3093), .I1(n3116), .CO(n29996));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n29756), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n29756), .I0(n2001), .I1(n2027), .CO(n29757));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n29755), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n29755), .I0(n2002), .I1(n2027), .CO(n29756));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n29994), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n29994), .I0(n3094), .I1(n3116), .CO(n29995));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n29754), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n29993), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n29754), .I0(n2003), .I1(n2027), .CO(n29755));
    SB_CARRY mod_5_add_2143_17 (.CI(n29993), .I0(n3095), .I1(n3116), .CO(n29994));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n29753), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n29992), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n29753), .I0(n2004), .I1(n2027), .CO(n29754));
    SB_CARRY mod_5_add_2143_16 (.CI(n29992), .I0(n3096), .I1(n3116), .CO(n29993));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n29991), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n29752), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n29991), .I0(n3097), .I1(n3116), .CO(n29992));
    SB_CARRY mod_5_add_1406_7 (.CI(n29752), .I0(n2005), .I1(n2027), .CO(n29753));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n29751), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n28444), .I0(bit_ctr[18]), .I1(GND_net), .CO(n28445));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n29990), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n29751), .I0(n2006), .I1(n2027), .CO(n29752));
    SB_CARRY mod_5_add_2143_14 (.CI(n29990), .I0(n3098), .I1(n3116), .CO(n29991));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n29989), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n29750), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut (.I0(n25771), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(\state[1] ), .O(n37679));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_4_lut (.I0(n30650), .I1(n15775), .I2(\neo_pixel_transmitter.done ), 
            .I3(start), .O(n1138));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff1f;
    SB_LUT4 i1_3_lut_4_lut (.I0(n15775), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n4_adj_4242), .O(n15887));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i37390_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44242));
    defparam i37390_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21046_2_lut_3_lut (.I0(n25553), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n25777));   // verilog/neopixel.v(22[26:36])
    defparam i21046_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i35085_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n36211), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17229));
    defparam i35085_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 i1_2_lut_3_lut (.I0(n25771), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n13454));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i29432_2_lut_3_lut (.I0(\state[0] ), .I1(n12), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n36197));
    defparam i29432_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i29424_2_lut_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n25553), .I2(n608), 
            .I3(bit_ctr[28]), .O(n36189));
    defparam i29424_2_lut_3_lut_4_lut.LUT_INIT = 16'h5600;
    SB_LUT4 i2794_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n36211), .I2(bit_ctr[27]), 
            .I3(n36154), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i2794_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31_2_lut_3_lut (.I0(\one_wire_N_513[11] ), .I1(n4), .I2(n15928), 
            .I3(GND_net), .O(n12));   // verilog/neopixel.v(6[16:24])
    defparam i31_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(n36154), .I1(n14417), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14417), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n36154), .O(n36288));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i35082_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n25777), .I2(n36211), 
            .I3(bit_ctr[28]), .O(n36154));
    defparam i35082_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 i20825_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n25553));   // verilog/neopixel.v(22[26:36])
    defparam i20825_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4244));
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'heeee;
    SB_LUT4 i20925_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n25655));
    defparam i20925_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1522 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4244), 
            .O(n30_adj_4245));
    defparam i13_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1523 (.I0(n2098), .I1(n25655), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4246));
    defparam i11_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1524 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4247));
    defparam i12_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1525 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4248));
    defparam i10_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1526 (.I0(n27_adj_4248), .I1(n29_adj_4247), .I2(n28_adj_4246), 
            .I3(n30_adj_4245), .O(n2126));
    defparam i16_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37386_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44238));
    defparam i37386_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37389_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44241));
    defparam i37389_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1527 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4249));
    defparam i1_2_lut_adj_1527.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4250));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1528 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4249), 
            .O(n16_adj_4251));
    defparam i7_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1529 (.I0(n1307), .I1(n16_adj_4251), .I2(n12_adj_4250), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i37388_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44240));
    defparam i37388_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1530 (.I0(n1205), .I1(n1202), .I2(n1206), .I3(n1208), 
            .O(n14_adj_4252));
    defparam i6_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1531 (.I0(bit_ctr[23]), .I1(n1207), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4253));
    defparam i1_3_lut_adj_1531.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1532 (.I0(n9_adj_4253), .I1(n14_adj_4252), .I2(n1203), 
            .I3(n1204), .O(n1235));
    defparam i7_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37387_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44239));
    defparam i37387_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20832_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n25561));
    defparam i20832_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n25561), .I3(n1108), 
            .O(n12_adj_4254));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1533 (.I0(n1107), .I1(n12_adj_4254), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1534 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4255));
    defparam i10_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1535 (.I0(n2203), .I1(n28_adj_4255), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4256));
    defparam i14_4_lut_adj_1535.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1536 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4257));
    defparam i12_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1537 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4258));
    defparam i13_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1538 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4259));
    defparam i11_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1539 (.I0(n29_adj_4259), .I1(n31_adj_4258), .I2(n30_adj_4257), 
            .I3(n32_adj_4256), .O(n2225));
    defparam i17_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i37385_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44237));
    defparam i37385_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4260));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1540 (.I0(bit_ctr[12]), .I1(n22_adj_4260), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4261));
    defparam i11_4_lut_adj_1540.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1541 (.I0(n2294), .I1(n30_adj_4261), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4262));
    defparam i15_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1542 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4263));
    defparam i13_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1543 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4264));
    defparam i14_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1544 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4265));
    defparam i12_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1545 (.I0(n31_adj_4265), .I1(n33_adj_4264), .I2(n32_adj_4263), 
            .I3(n34_adj_4262), .O(n2324));
    defparam i18_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i37384_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44236));
    defparam i37384_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37355_2_lut (.I0(n31958), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i37355_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37383_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44235));
    defparam i37383_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37357_2_lut (.I0(n31958), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i37357_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n31958), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32312_3_lut (.I0(n905), .I1(n906), .I2(n36288), .I3(GND_net), 
            .O(n39093));
    defparam i32312_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n39093), .I2(n17229), .I3(n14415), 
            .O(n31958));
    defparam i4_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n31958), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14415), .I1(n971[27]), .I2(n31958), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32320_3_lut (.I0(n971[31]), .I1(n971[28]), .I2(n971[29]), 
            .I3(GND_net), .O(n39101));
    defparam i32320_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6_adj_4266));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n31958), .I1(n6_adj_4266), .I2(n1005), .I3(n39101), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i37353_2_lut (.I0(n31958), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4228));   // verilog/neopixel.v(22[26:36])
    defparam i37353_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i34188_2_lut (.I0(bit_ctr[2]), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(GND_net), .O(n41043));
    defparam i34188_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i20915_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n25645));
    defparam i20915_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1546 (.I0(n3185), .I1(n3195), .I2(n3192), .I3(n3191), 
            .O(n48_adj_4267));
    defparam i20_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1547 (.I0(n3205), .I1(n3202), .I2(n3186), .I3(n3194), 
            .O(n46_adj_4268));
    defparam i18_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1548 (.I0(n3201), .I1(n3182), .I2(n3200), .I3(n3190), 
            .O(n47_adj_4269));
    defparam i19_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1549 (.I0(n3197), .I1(n3199), .I2(n3196), .I3(n3184), 
            .O(n45));
    defparam i17_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1550 (.I0(n3206), .I1(n3208), .I2(n3183), .I3(n3188), 
            .O(n44));
    defparam i16_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1551 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n25645), 
            .O(n43_adj_4270));
    defparam i15_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_4269), .I2(n46_adj_4268), 
            .I3(n48_adj_4267), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1552 (.I0(n3204), .I1(n3207), .I2(n3187), .I3(n3203), 
            .O(n49_adj_4271));
    defparam i21_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4271), .I1(n54), .I2(n43_adj_4270), 
            .I3(n44), .O(n25737));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i241_2_lut (.I0(n12), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n1141));   // verilog/neopixel.v(103[9] 111[12])
    defparam i241_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1553 (.I0(n8), .I1(n36197), .I2(\state[1] ), 
            .I3(n25771), .O(n17312));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1553.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1554 (.I0(\state[0] ), .I1(n13454), .I2(n1141), 
            .I3(\state[1] ), .O(n17058));
    defparam i1_4_lut_adj_1554.LUT_INIT = 16'haf33;
    SB_LUT4 i34779_3_lut (.I0(\color[20] ), .I1(bit_ctr[0]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41235));   // verilog/neopixel.v(22[26:36])
    defparam i34779_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i34465_3_lut (.I0(\color[4] ), .I1(bit_ctr[0]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41231));   // verilog/neopixel.v(22[26:36])
    defparam i34465_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 color_bit_I_0_i9_3_lut (.I0(\color[10] ), .I1(\color[11] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n9_adj_4273));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8366_rep_547_2_lut (.I0(bit_ctr[0]), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(GND_net), .O(n45277));   // verilog/neopixel.v(22[26:36])
    defparam i8366_rep_547_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35813_4_lut (.I0(\color[9] ), .I1(n9_adj_4273), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n42667));
    defparam i35813_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 color_bit_I_0_i18_4_lut (.I0(\color[17] ), .I1(n41235), .I2(bit_ctr[2]), 
            .I3(bit_ctr[0]), .O(n18_adj_4274));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i23749_rep_541_2_lut (.I0(bit_ctr[3]), .I1(n25737), .I2(GND_net), 
            .I3(GND_net), .O(n45271));   // verilog/neopixel.v(22[26:36])
    defparam i23749_rep_541_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 color_bit_I_0_i17_3_lut (.I0(\color[18] ), .I1(\color[19] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n17_adj_4275));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 color_bit_I_0_i3_4_lut (.I0(\color[1] ), .I1(n41231), .I2(bit_ctr[2]), 
            .I3(bit_ctr[0]), .O(n3_adj_4276));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i3_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 color_bit_I_0_i2_3_lut (.I0(\color[2] ), .I1(\color[3] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n2_adj_4277));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35608_4_lut (.I0(n42667), .I1(\color[12] ), .I2(bit_ctr[2]), 
            .I3(n45277), .O(n42462));
    defparam i35608_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32342_3_lut (.I0(n2_adj_4277), .I1(n3_adj_4276), .I2(n41043), 
            .I3(GND_net), .O(n39195));
    defparam i32342_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35024_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n25737), .I3(GND_net), 
            .O(color_bit_N_556[4]));
    defparam i35024_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i35591_4_lut (.I0(n17_adj_4275), .I1(n45271), .I2(n18_adj_4274), 
            .I3(n41043), .O(n41303));
    defparam i35591_4_lut.LUT_INIT = 16'h2230;
    SB_LUT4 i36203_4_lut (.I0(n39195), .I1(n42462), .I2(bit_ctr[3]), .I3(n25737), 
            .O(n43057));   // verilog/neopixel.v(22[26:36])
    defparam i36203_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i19969_4_lut (.I0(n43057), .I1(\state_3__N_362[1] ), .I2(n41303), 
            .I3(color_bit_N_556[4]), .O(state_3__N_362[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i19969_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14415));
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'h9999;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i20781_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i20781_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n25553), .I2(n36189), .I3(n608), 
            .O(n36211));
    defparam i2_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(bit_ctr[28]), .I1(n36211), .I2(GND_net), 
            .I3(GND_net), .O(n14417));
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'h9999;
    SB_LUT4 i32198_3_lut (.I0(n36211), .I1(n708), .I2(n36189), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i32198_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i2_2_lut (.I0(n2407), .I1(n2405), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4278));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1557 (.I0(n2390), .I1(n2400), .I2(n2393), .I3(n2394), 
            .O(n32_adj_4279));
    defparam i12_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i20941_2_lut (.I0(bit_ctr[11]), .I1(n2409), .I2(GND_net), 
            .I3(GND_net), .O(n25671));
    defparam i20941_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16_4_lut_adj_1558 (.I0(n2398), .I1(n32_adj_4279), .I2(n22_adj_4278), 
            .I3(n2403), .O(n36_adj_4280));
    defparam i16_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1559 (.I0(n2406), .I1(n2399), .I2(n2391), .I3(n2396), 
            .O(n34_adj_4281));
    defparam i14_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1560 (.I0(n2401), .I1(n2392), .I2(n2395), .I3(n25671), 
            .O(n35_adj_4282));
    defparam i15_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1561 (.I0(n2402), .I1(n2404), .I2(n2408), .I3(n2397), 
            .O(n33_adj_4283));
    defparam i13_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1562 (.I0(n33_adj_4283), .I1(n35_adj_4282), .I2(n34_adj_4281), 
            .I3(n36_adj_4280), .O(n2423));
    defparam i19_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37382_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44234));
    defparam i37382_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(bit_ctr[10]), .I1(n2506), .I2(n2509), .I3(GND_net), 
            .O(n26_adj_4284));
    defparam i5_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i12_4_lut_adj_1563 (.I0(n2496), .I1(n2502), .I2(n2498), .I3(n2489), 
            .O(n33_adj_4285));
    defparam i12_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(n2505), .I1(n2503), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4286));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1565 (.I0(n33_adj_4285), .I1(n2494), .I2(n26_adj_4284), 
            .I3(n2507), .O(n38_adj_4287));
    defparam i17_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1566 (.I0(n2501), .I1(n2497), .I2(n2490), .I3(n2491), 
            .O(n36_adj_4288));
    defparam i15_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1567 (.I0(n2504), .I1(n2508), .I2(n2493), .I3(n22_adj_4286), 
            .O(n37_adj_4289));
    defparam i16_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1568 (.I0(n2500), .I1(n2499), .I2(n2495), .I3(n2492), 
            .O(n35_adj_4290));
    defparam i14_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1569 (.I0(n35_adj_4290), .I1(n37_adj_4289), .I2(n36_adj_4288), 
            .I3(n38_adj_4287), .O(n2522));
    defparam i20_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37380_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44232));
    defparam i37380_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37379_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44231));
    defparam i37379_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1570 (.I0(bit_ctr[22]), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4291));
    defparam i2_2_lut_adj_1570.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1571 (.I0(bit_ctr[31]), .I1(bit_ctr[12]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[20]), .O(n48_adj_4292));
    defparam i20_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1572 (.I0(bit_ctr[26]), .I1(bit_ctr[5]), .I2(bit_ctr[17]), 
            .I3(bit_ctr[25]), .O(n46_adj_4293));
    defparam i18_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1573 (.I0(bit_ctr[14]), .I1(bit_ctr[28]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[21]), .O(n47_adj_4294));
    defparam i19_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1574 (.I0(bit_ctr[15]), .I1(bit_ctr[8]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[18]), .O(n45_adj_4295));
    defparam i17_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1575 (.I0(bit_ctr[6]), .I1(bit_ctr[9]), .I2(bit_ctr[10]), 
            .I3(bit_ctr[19]), .O(n44_adj_4296));
    defparam i16_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1576 (.I0(bit_ctr[3]), .I1(n30_adj_4291), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43_adj_4297));
    defparam i15_4_lut_adj_1576.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut_adj_1577 (.I0(n45_adj_4295), .I1(n47_adj_4294), .I2(n46_adj_4293), 
            .I3(n48_adj_4292), .O(n54_adj_4298));
    defparam i26_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1578 (.I0(bit_ctr[30]), .I1(bit_ctr[7]), .I2(bit_ctr[23]), 
            .I3(bit_ctr[24]), .O(n49_adj_4299));
    defparam i21_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1579 (.I0(n49_adj_4299), .I1(n54_adj_4298), .I2(n43_adj_4297), 
            .I3(n44_adj_4296), .O(\state_3__N_362[1] ));
    defparam i27_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i2063_3_lut (.I0(n15887), .I1(\state_3__N_362[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4443));
    defparam i2063_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_4_lut_adj_1580 (.I0(\state[1] ), .I1(n1138), .I2(n4443), 
            .I3(\state[0] ), .O(n4472));
    defparam i2_4_lut_adj_1580.LUT_INIT = 16'hf0ee;
    SB_LUT4 i5_3_lut_adj_1581 (.I0(n2986), .I1(bit_ctr[5]), .I2(n3009), 
            .I3(GND_net), .O(n31_adj_4300));
    defparam i5_3_lut_adj_1581.LUT_INIT = 16'heaea;
    SB_LUT4 i15_4_lut_adj_1582 (.I0(n2996), .I1(n3006), .I2(n3003), .I3(n2989), 
            .O(n41_adj_4301));
    defparam i15_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1583 (.I0(n2999), .I1(n2991), .I2(n2984), .I3(n2998), 
            .O(n40_adj_4302));
    defparam i14_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1584 (.I0(n3002), .I1(n2993), .I2(n3008), .I3(n3005), 
            .O(n45_adj_4303));
    defparam i19_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1585 (.I0(n3004), .I1(n2985), .I2(n2994), .I3(n2987), 
            .O(n44_adj_4304));
    defparam i18_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1586 (.I0(n2995), .I1(n3007), .I2(n2997), .I3(n3001), 
            .O(n43_adj_4305));
    defparam i17_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1587 (.I0(n41_adj_4301), .I1(n31_adj_4300), .I2(n2992), 
            .I3(n2990), .O(n47_adj_4306));
    defparam i21_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1588 (.I0(n45_adj_4303), .I1(n3000), .I2(n40_adj_4302), 
            .I3(n2988), .O(n49_adj_4307));
    defparam i23_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_adj_4307), .I1(n47_adj_4306), .I2(n43_adj_4305), 
            .I3(n44_adj_4304), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37365_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44217));
    defparam i37365_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1589 (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[4]), 
            .I2(one_wire_N_513[2]), .I3(GND_net), .O(n30650));
    defparam i2_3_lut_adj_1589.LUT_INIT = 16'h8080;
    SB_LUT4 i20981_2_lut (.I0(n30650), .I1(n15775), .I2(GND_net), .I3(GND_net), 
            .O(n25711));
    defparam i20981_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1590 (.I0(n30771), .I1(one_wire_N_513[4]), .I2(one_wire_N_513[3]), 
            .I3(GND_net), .O(n4_adj_4242));
    defparam i1_3_lut_adj_1590.LUT_INIT = 16'hecec;
    SB_LUT4 equal_342_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n8));
    defparam equal_342_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut_adj_1591 (.I0(n15928), .I1(\one_wire_N_513[11] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4308));   // verilog/neopixel.v(104[14:39])
    defparam i2_2_lut_adj_1591.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(one_wire_N_513[9]), .I1(\one_wire_N_513[5] ), 
            .I2(n6_adj_4308), .I3(\one_wire_N_513[6] ), .O(n6_adj_4309));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1593 (.I0(one_wire_N_513[10]), .I1(\one_wire_N_513[8] ), 
            .I2(\one_wire_N_513[7] ), .I3(n6_adj_4309), .O(n15775));   // verilog/neopixel.v(104[14:39])
    defparam i4_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i29434_2_lut (.I0(\state[1] ), .I1(n15887), .I2(GND_net), 
            .I3(GND_net), .O(n36199));
    defparam i29434_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1594 (.I0(n15928), .I1(n35266), .I2(n36306), 
            .I3(\state[1] ), .O(n17075));
    defparam i1_4_lut_adj_1594.LUT_INIT = 16'h0544;
    SB_LUT4 i104_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_576 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i104_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37377_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44229));
    defparam i37377_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29419_4_lut (.I0(n15775), .I1(n30650), .I2(n4_adj_4242), 
            .I3(\state[0] ), .O(n25771));   // verilog/neopixel.v(36[4] 116[11])
    defparam i29419_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i23_3_lut (.I0(n4_adj_4242), .I1(n30650), .I2(\state[0] ), 
            .I3(GND_net), .O(n36207));
    defparam i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1595 (.I0(n25417), .I1(\state[1] ), .I2(n15775), 
            .I3(n36207), .O(n37638));
    defparam i3_4_lut_adj_1595.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut_adj_1596 (.I0(\state[1] ), .I1(n37638), .I2(start), 
            .I3(n37679), .O(n36865));
    defparam i2_4_lut_adj_1596.LUT_INIT = 16'h8c00;
    SB_LUT4 mux_680_Mux_0_i3_3_lut_3_lut (.I0(\neo_pixel_transmitter.done ), 
            .I1(start), .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_680_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'ha1a1;
    SB_LUT4 i26_4_lut_adj_1597 (.I0(n47_adj_4226), .I1(n49), .I2(n48), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n18036, PWMLimit, clk32MHz, \data_out_frame[17] , GND_net, 
            n18035, n18034, n18033, n18032, n18031, n18030, \data_out_frame[15] , 
            \data_out_frame[19] , n18029, n18028, n18027, \data_in_frame[17] , 
            n17973, \data_in_frame[15] , n17902, \data_in_frame[6] , 
            n17972, \data_out_frame[16] , \data_out_frame[10] , \data_out_frame[14] , 
            \data_out_frame[13] , \data_out_frame[11] , n17933, \data_in_frame[10] , 
            n17932, n17901, n17931, n17930, \data_in_frame[9] , n17929, 
            n17928, n17927, \data_out_frame[8] , \data_out_frame[12] , 
            n17900, \data_out_frame[6] , \data_out_frame[9] , \data_out_frame[4][1] , 
            \data_out_frame[4][0] , n18153, setpoint, n18154, n18155, 
            n18156, n18157, n18158, n18142, n18143, n17515, n17548, 
            n17554, n17551, n17560, n17557, n17563, n18159, n18160, 
            n18144, n18145, n18146, n18147, n18148, n18149, n18150, 
            n18151, n18152, n18140, n18141, n18138, n18139, n17926, 
            n17925, n18108, VCC_net, \byte_transmit_counter[0] , n17899, 
            n18037, n18038, n18039, n18040, n18041, n18042, n17898, 
            \data_in_frame[5] , n17897, n17896, n17895, n44420, n44421, 
            n17971, n17970, \data_in_frame[14] , n17969, n17968, n17967, 
            n17966, n17894, n17893, n17892, n18048, n18049, n18046, 
            n18047, n17891, n18043, n18044, n18045, n17890, \data_in_frame[4] , 
            n17889, n17888, n17887, n17886, n17885, n17884, n17883, 
            n17882, \data_in_frame[3] , n17881, n17880, n17879, n17965, 
            n17878, n17877, n17876, n17875, n17964, n17874, \data_in_frame[2] , 
            n17873, n17872, n17871, n17870, n17924, n17869, n17923, 
            n17868, n17867, n17866, \data_in_frame[1] , n17922, \data_in_frame[8] , 
            n17921, \data_out_frame[5] , n17920, \data_out_frame[4][2] , 
            \data_out_frame[7] , n17919, n17918, n17917, n17916, n17915, 
            n17914, \data_in_frame[7] , n17913, n17912, n17911, n17910, 
            n17909, n17908, n17907, n17906, n17905, n17904, n17865, 
            \data_out_frame[18] , n17864, n17863, n17862, n17861, 
            n17860, n17859, n17963, n17858, \data_in_frame[0] , n17857, 
            n17856, n17855, n17854, n17853, n17852, n17851, control_mode, 
            n17850, n17849, n17848, n17962, \data_in_frame[13] , n17847, 
            n17846, n17845, n17844, \data_out_frame[20] , n17843, 
            n17842, n17841, n17840, n17839, n17838, n17837, rx_data_ready, 
            n17836, n17835, n17974, n17961, \data_out_frame[16][3] , 
            n17834, \data_out_frame[16][5] , n17833, n17832, n17831, 
            \FRAME_MATCHER.state[0] , n17513, n17546, n17549, n17552, 
            n17960, n17959, n17958, n17830, n17555, n17558, n17561, 
            n7821, n17829, n17828, n17827, n17826, n17825, n17824, 
            n17823, n17822, n17821, n17820, n17819, n13293, n17818, 
            n17817, n17816, n17815, n17814, n17813, n17812, n17811, 
            n17810, n17809, n17808, n17806, \data_out_frame[16][1] , 
            n17805, \data_out_frame[16][0] , n17804, n17803, n17802, 
            n17801, n17800, n17799, n17798, n17797, n17796, n17795, 
            n17794, n17793, n17792, n17791, n17790, n17789, n17788, 
            n17787, n17978, n17786, n17785, n17784, n17977, n17976, 
            n17783, n17782, n17781, n17780, n17779, n17778, n17777, 
            n17776, n17775, n17774, n17773, n17772, n17771, n17770, 
            n17769, n17768, n17767, n17766, n17765, n17764, n17763, 
            n17762, n17761, n17760, n17759, n17758, n17757, n17756, 
            \FRAME_MATCHER.i_31__N_2390 , n17755, n17754, n17753, n17752, 
            n17751, n17750, n17749, n17748, n17747, n17746, n17745, 
            n17744, n17743, ID1, ID0, n17742, n17741, n17740, 
            n17739, n17738, n17737, n17736, n17735, n17734, n17733, 
            n17732, ID2, n17731, n17730, n17729, \data_in_frame[12] , 
            n17728, n17727, n17726, n17725, \data_in_frame[11] , n17724, 
            n17723, n17722, n17721, n17720, n17719, n17718, n17717, 
            n17716, n17715, n17714, n17713, \data_in[3] , n17712, 
            n17711, n17710, n17709, n17708, n17707, n17706, n17705, 
            \data_in[2] , n17704, n17703, n17702, n17701, n17700, 
            n17699, n17698, n17697, \data_in[1] , n17696, n17695, 
            n17694, n17693, n17692, n17691, n17690, n17689, \data_in[0] , 
            n17688, n17687, n17686, n17685, n17684, n17683, n17682, 
            \Ki[7] , n17681, \Ki[6] , n17680, \Ki[5] , n17679, \Ki[4] , 
            n17678, \Ki[3] , n17677, \Ki[2] , n17676, \Ki[1] , n122, 
            n2855, n63, n5, n3741, \FRAME_MATCHER.state_31__N_2586[2] , 
            n17675, \Kp[7] , n17674, \Kp[6] , n17673, \Kp[5] , n17672, 
            \Kp[4] , n17671, \Kp[3] , n17670, \Kp[2] , n17669, \Kp[1] , 
            n17668, gearBoxRatio, n17667, n17666, n17665, n17664, 
            n17663, n17662, n17661, n17660, n17659, n17658, n17657, 
            n17656, n17655, n17654, n17653, n17652, n17651, n17650, 
            n17649, n17648, n17647, n17646, n17645, IntegralLimit, 
            n17644, n17643, n17642, n17641, n17640, n17639, n17638, 
            n17637, n17636, n17635, n17634, \FRAME_MATCHER.i_31__N_2388 , 
            n2778, n17633, n17632, n17631, n17630, n17629, n17628, 
            n17627, n17626, n17625, n17624, n17957, n737, \data_in_frame[18] , 
            \data_in_frame[19] , n17100, n17068, n17935, n17956, n17955, 
            n17623, n17954, n123, n10454, n17953, n17952, n17951, 
            n17950, n17949, n17948, n17947, n17946, n17945, n17944, 
            n17943, n17942, n17941, n17975, LED_c, n97, n16, n7, 
            n17934, \FRAME_MATCHER.state_31__N_2458[1] , n17940, n17939, 
            n17938, n17937, n17936, n17390, n17903, n4380, rx_data, 
            n4379, n4382, n4381, n17538, n34728, n17522, n17521, 
            n17520, n17519, n17518, \Ki[0] , n17517, \Kp[0] , n17516, 
            n61, n4393, n4392, n4391, n4390, n4389, n4388, n4387, 
            n4386, n4385, n4401, n4400, n35431, n35432, n35433, 
            n35430, n35434, n35429, n38107, \duty[10] , n35428, 
            n35435, n4378, n35419, n35423, n35420, n35416, n35417, 
            n4384, n4383, n35421, n35422, n35418, n4399, n4398, 
            n4397, n4396, n4395, n38059, n4394, tx_active, n17466, 
            \r_Clock_Count[6] , n17463, \r_Clock_Count[7] , n17481, 
            \r_Clock_Count[1] , n17512, r_Bit_Index, n17509, n18130, 
            r_SM_Main, n18105, tx_o, tx_enable, n19634, n17529, 
            n17528, n541, n314, n315, n320, o_Tx_Serial_N_3351, 
            n17108, n4683, n17186, n17330, n35270, r_Clock_Count, 
            n35268, n35273, n18165, n35086, n35088, n35090, n35000, 
            n34912, n34804, n34716, n17566, r_Bit_Index_adj_14, n17569, 
            n35004, n18111, n25741, r_SM_Main_adj_15, n35269, r_Rx_Data, 
            n35272, PIN_13_N_105, n35275, n35276, n35271, n35274, 
            n41248, n41247, n17576, n17575, n17574, n17573, n17572, 
            n17571, n17570, n17527, n17180, n17321, n4661, n35374, 
            n25555, n1, n24764, n4, n4_adj_12, n15912, n15917, 
            n4_adj_13, n6, n44844) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18036;
    output [23:0]PWMLimit;
    input clk32MHz;
    output [7:0]\data_out_frame[17] ;
    input GND_net;
    input n18035;
    input n18034;
    input n18033;
    input n18032;
    input n18031;
    input n18030;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[19] ;
    input n18029;
    input n18028;
    input n18027;
    output [7:0]\data_in_frame[17] ;
    input n17973;
    output [7:0]\data_in_frame[15] ;
    input n17902;
    output [7:0]\data_in_frame[6] ;
    input n17972;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[11] ;
    input n17933;
    output [7:0]\data_in_frame[10] ;
    input n17932;
    input n17901;
    input n17931;
    input n17930;
    output [7:0]\data_in_frame[9] ;
    input n17929;
    input n17928;
    input n17927;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[12] ;
    input n17900;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[9] ;
    output \data_out_frame[4][1] ;
    output \data_out_frame[4][0] ;
    input n18153;
    output [23:0]setpoint;
    input n18154;
    input n18155;
    input n18156;
    input n18157;
    input n18158;
    input n18142;
    input n18143;
    input n17515;
    input n17548;
    input n17554;
    input n17551;
    input n17560;
    input n17557;
    input n17563;
    input n18159;
    input n18160;
    input n18144;
    input n18145;
    input n18146;
    input n18147;
    input n18148;
    input n18149;
    input n18150;
    input n18151;
    input n18152;
    input n18140;
    input n18141;
    input n18138;
    input n18139;
    input n17926;
    input n17925;
    input n18108;
    input VCC_net;
    output \byte_transmit_counter[0] ;
    input n17899;
    input n18037;
    input n18038;
    input n18039;
    input n18040;
    input n18041;
    input n18042;
    input n17898;
    output [7:0]\data_in_frame[5] ;
    input n17897;
    input n17896;
    input n17895;
    input n44420;
    input n44421;
    input n17971;
    input n17970;
    output [7:0]\data_in_frame[14] ;
    input n17969;
    input n17968;
    input n17967;
    input n17966;
    input n17894;
    input n17893;
    input n17892;
    input n18048;
    input n18049;
    input n18046;
    input n18047;
    input n17891;
    input n18043;
    input n18044;
    input n18045;
    input n17890;
    output [7:0]\data_in_frame[4] ;
    input n17889;
    input n17888;
    input n17887;
    input n17886;
    input n17885;
    input n17884;
    input n17883;
    input n17882;
    output [7:0]\data_in_frame[3] ;
    input n17881;
    input n17880;
    input n17879;
    input n17965;
    input n17878;
    input n17877;
    input n17876;
    input n17875;
    input n17964;
    input n17874;
    output [7:0]\data_in_frame[2] ;
    input n17873;
    input n17872;
    input n17871;
    input n17870;
    input n17924;
    input n17869;
    input n17923;
    input n17868;
    input n17867;
    input n17866;
    output [7:0]\data_in_frame[1] ;
    input n17922;
    output [7:0]\data_in_frame[8] ;
    input n17921;
    output [7:0]\data_out_frame[5] ;
    input n17920;
    output \data_out_frame[4][2] ;
    output [7:0]\data_out_frame[7] ;
    input n17919;
    input n17918;
    input n17917;
    input n17916;
    input n17915;
    input n17914;
    output [7:0]\data_in_frame[7] ;
    input n17913;
    input n17912;
    input n17911;
    input n17910;
    input n17909;
    input n17908;
    input n17907;
    input n17906;
    input n17905;
    input n17904;
    input n17865;
    output [7:0]\data_out_frame[18] ;
    input n17864;
    input n17863;
    input n17862;
    input n17861;
    input n17860;
    input n17859;
    input n17963;
    input n17858;
    output [7:0]\data_in_frame[0] ;
    input n17857;
    input n17856;
    input n17855;
    input n17854;
    input n17853;
    input n17852;
    input n17851;
    output [7:0]control_mode;
    input n17850;
    input n17849;
    input n17848;
    input n17962;
    output [7:0]\data_in_frame[13] ;
    input n17847;
    input n17846;
    input n17845;
    input n17844;
    output [7:0]\data_out_frame[20] ;
    input n17843;
    input n17842;
    input n17841;
    input n17840;
    input n17839;
    input n17838;
    input n17837;
    output rx_data_ready;
    input n17836;
    input n17835;
    input n17974;
    input n17961;
    output \data_out_frame[16][3] ;
    input n17834;
    output \data_out_frame[16][5] ;
    input n17833;
    input n17832;
    input n17831;
    output \FRAME_MATCHER.state[0] ;
    output n17513;
    output n17546;
    output n17549;
    output n17552;
    input n17960;
    input n17959;
    input n17958;
    input n17830;
    output n17555;
    output n17558;
    output n17561;
    output n7821;
    input n17829;
    input n17828;
    input n17827;
    input n17826;
    input n17825;
    input n17824;
    input n17823;
    input n17822;
    input n17821;
    input n17820;
    input n17819;
    output n13293;
    input n17818;
    input n17817;
    input n17816;
    input n17815;
    input n17814;
    input n17813;
    input n17812;
    input n17811;
    input n17810;
    input n17809;
    input n17808;
    input n17806;
    output \data_out_frame[16][1] ;
    input n17805;
    output \data_out_frame[16][0] ;
    input n17804;
    input n17803;
    input n17802;
    input n17801;
    input n17800;
    input n17799;
    input n17798;
    input n17797;
    input n17796;
    input n17795;
    input n17794;
    input n17793;
    input n17792;
    input n17791;
    input n17790;
    input n17789;
    input n17788;
    input n17787;
    input n17978;
    input n17786;
    input n17785;
    input n17784;
    input n17977;
    input n17976;
    input n17783;
    input n17782;
    input n17781;
    input n17780;
    input n17779;
    input n17778;
    input n17777;
    input n17776;
    input n17775;
    input n17774;
    input n17773;
    input n17772;
    input n17771;
    input n17770;
    input n17769;
    input n17768;
    input n17767;
    input n17766;
    input n17765;
    input n17764;
    input n17763;
    input n17762;
    input n17761;
    input n17760;
    input n17759;
    input n17758;
    input n17757;
    input n17756;
    output \FRAME_MATCHER.i_31__N_2390 ;
    input n17755;
    input n17754;
    input n17753;
    input n17752;
    input n17751;
    input n17750;
    input n17749;
    input n17748;
    input n17747;
    input n17746;
    input n17745;
    input n17744;
    input n17743;
    input ID1;
    input ID0;
    input n17742;
    input n17741;
    input n17740;
    input n17739;
    input n17738;
    input n17737;
    input n17736;
    input n17735;
    input n17734;
    input n17733;
    input n17732;
    input ID2;
    input n17731;
    input n17730;
    input n17729;
    output [7:0]\data_in_frame[12] ;
    input n17728;
    input n17727;
    input n17726;
    input n17725;
    output [7:0]\data_in_frame[11] ;
    input n17724;
    input n17723;
    input n17722;
    input n17721;
    input n17720;
    input n17719;
    input n17718;
    input n17717;
    input n17716;
    input n17715;
    input n17714;
    input n17713;
    output [7:0]\data_in[3] ;
    input n17712;
    input n17711;
    input n17710;
    input n17709;
    input n17708;
    input n17707;
    input n17706;
    input n17705;
    output [7:0]\data_in[2] ;
    input n17704;
    input n17703;
    input n17702;
    input n17701;
    input n17700;
    input n17699;
    input n17698;
    input n17697;
    output [7:0]\data_in[1] ;
    input n17696;
    input n17695;
    input n17694;
    input n17693;
    input n17692;
    input n17691;
    input n17690;
    input n17689;
    output [7:0]\data_in[0] ;
    input n17688;
    input n17687;
    input n17686;
    input n17685;
    input n17684;
    input n17683;
    input n17682;
    output \Ki[7] ;
    input n17681;
    output \Ki[6] ;
    input n17680;
    output \Ki[5] ;
    input n17679;
    output \Ki[4] ;
    input n17678;
    output \Ki[3] ;
    input n17677;
    output \Ki[2] ;
    input n17676;
    output \Ki[1] ;
    output n122;
    output n2855;
    output n63;
    output n5;
    output n3741;
    output \FRAME_MATCHER.state_31__N_2586[2] ;
    input n17675;
    output \Kp[7] ;
    input n17674;
    output \Kp[6] ;
    input n17673;
    output \Kp[5] ;
    input n17672;
    output \Kp[4] ;
    input n17671;
    output \Kp[3] ;
    input n17670;
    output \Kp[2] ;
    input n17669;
    output \Kp[1] ;
    input n17668;
    output [23:0]gearBoxRatio;
    input n17667;
    input n17666;
    input n17665;
    input n17664;
    input n17663;
    input n17662;
    input n17661;
    input n17660;
    input n17659;
    input n17658;
    input n17657;
    input n17656;
    input n17655;
    input n17654;
    input n17653;
    input n17652;
    input n17651;
    input n17650;
    input n17649;
    input n17648;
    input n17647;
    input n17646;
    input n17645;
    output [23:0]IntegralLimit;
    input n17644;
    input n17643;
    input n17642;
    input n17641;
    input n17640;
    input n17639;
    input n17638;
    input n17637;
    input n17636;
    input n17635;
    input n17634;
    output \FRAME_MATCHER.i_31__N_2388 ;
    output n2778;
    input n17633;
    input n17632;
    input n17631;
    input n17630;
    input n17629;
    input n17628;
    input n17627;
    input n17626;
    input n17625;
    input n17624;
    input n17957;
    output n737;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[19] ;
    output n17100;
    output n17068;
    input n17935;
    input n17956;
    input n17955;
    input n17623;
    input n17954;
    output n123;
    output n10454;
    input n17953;
    input n17952;
    input n17951;
    input n17950;
    input n17949;
    input n17948;
    input n17947;
    input n17946;
    input n17945;
    input n17944;
    input n17943;
    input n17942;
    input n17941;
    input n17975;
    output LED_c;
    output n97;
    output n16;
    output n7;
    input n17934;
    output \FRAME_MATCHER.state_31__N_2458[1] ;
    input n17940;
    input n17939;
    input n17938;
    input n17937;
    input n17936;
    input n17390;
    input n17903;
    output n4380;
    output [7:0]rx_data;
    output n4379;
    output n4382;
    output n4381;
    input n17538;
    input n34728;
    input n17522;
    input n17521;
    input n17520;
    input n17519;
    input n17518;
    output \Ki[0] ;
    input n17517;
    output \Kp[0] ;
    input n17516;
    output n61;
    output n4393;
    output n4392;
    output n4391;
    output n4390;
    output n4389;
    output n4388;
    output n4387;
    output n4386;
    output n4385;
    output n4401;
    output n4400;
    output n35431;
    output n35432;
    output n35433;
    output n35430;
    output n35434;
    output n35429;
    output n38107;
    input \duty[10] ;
    output n35428;
    output n35435;
    output n4378;
    output n35419;
    output n35423;
    output n35420;
    output n35416;
    output n35417;
    output n4384;
    output n4383;
    output n35421;
    output n35422;
    output n35418;
    output n4399;
    output n4398;
    output n4397;
    output n4396;
    output n4395;
    output n38059;
    output n4394;
    output tx_active;
    input n17466;
    output \r_Clock_Count[6] ;
    input n17463;
    output \r_Clock_Count[7] ;
    input n17481;
    output \r_Clock_Count[1] ;
    input n17512;
    output [2:0]r_Bit_Index;
    input n17509;
    input n18130;
    output [2:0]r_SM_Main;
    input n18105;
    output tx_o;
    output tx_enable;
    output n19634;
    input n17529;
    input n17528;
    output n541;
    output n314;
    output n315;
    output n320;
    output o_Tx_Serial_N_3351;
    output n17108;
    output n4683;
    output n17186;
    output n17330;
    output n35270;
    output [7:0]r_Clock_Count;
    input n35268;
    output n35273;
    input n18165;
    input n35086;
    input n35088;
    input n35090;
    input n35000;
    input n34912;
    input n34804;
    input n34716;
    input n17566;
    output [2:0]r_Bit_Index_adj_14;
    input n17569;
    input n35004;
    input n18111;
    input n25741;
    output [2:0]r_SM_Main_adj_15;
    output n35269;
    output r_Rx_Data;
    output n35272;
    input PIN_13_N_105;
    output n35275;
    output n35276;
    output n35271;
    output n35274;
    output n41248;
    output n41247;
    input n17576;
    input n17575;
    input n17574;
    input n17573;
    input n17572;
    input n17571;
    input n17570;
    input n17527;
    output n17180;
    output n17321;
    output n4661;
    output n35374;
    output n25555;
    output n1;
    output n24764;
    output n4;
    output n4_adj_12;
    output n15912;
    output n15917;
    output n4_adj_13;
    output n6;
    output n44844;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n35619, n15522, n31104, n35673, n10, n28488;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n28489, n37402, n2, n2086, n17991, n31150, n35934, n10_adj_3893, 
        n2_adj_3894, n3, n18026;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n18025, n18024, n18023, n2_adj_3895, n28487, n18022, n7_c, 
        n35954, n35727, n37444, n1640, n36002, n36077, n35679, 
        n12, n36080, n16234, n35904, n35670, n35765, n35947, n31973, 
        n31142, n12_adj_3896, n16238, n31164, n36742, n35881, n1117, 
        n16_c, n35613, n36011, n16898, n17, n16042, n35918, n35547, 
        n36038, n35781, n10_adj_3897, n35864, n35826;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n35993, n30880;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n16403, n16698, n37377, n15502, n18, n30, n17990, n28, 
        n36008, n35823, n35870, n35542, n29, n36014, n36044, n35504, 
        n35937, n27, n1829, n35700, n2_adj_3898, n28486, n6_c, 
        n35571, n36035, n36068, n10_adj_3899, n35462, n35878, n10_adj_3900, 
        n31109, n16022, n35978, n28_adj_3901, n16394, n15489, n35691, 
        n43485, n16052, n30_adj_3902, n35684, n35478, n31, n35907, 
        n31090, n35604, n29_adj_3903, n32, n35753, n35657, n8, 
        n12_adj_3904, n1048, n12_adj_3905, n32044, n8_adj_3906, n35749, 
        n31802, n4_c, n36047, n6_adj_3907, n31168, n37260, n35846, 
        n16094, n32004, n35756, n30877, n35940, n14, n10_adj_3908, 
        n36725, n16535, n35558, n35513, n12_adj_3909, n13, n35913, 
        n16711, n31684, n35484, n32079, n35960, n6_adj_3910, n37263, 
        n39251, n39249, n39204, n2_adj_3911, n28485, n35833, n2_adj_3912, 
        n28484, n35487, n12_adj_3913, n12_adj_3914, n36029, n16_adj_3915, 
        n36083, n17_adj_3916, n18021, n14104, n35580, n36089, n35950, 
        n35465, n39242, n39240, n39201, n39232;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n19;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n39187, n39233, n39231, n44385, n44247, n42806, n32007, 
        n36937, n44337, n39188, n18020, n35507;
    wire [7:0]\data_out_frame[16]_c ;   // verilog/coms.v(95[12:26])
    
    wire n14_adj_3917, n8_adj_3918, n1238, n43499, n10_adj_3919, n35850, 
        n16704, n39198, n43063, n35778;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    wire [0:0]n3299;
    wire [2:0]r_SM_Main_2__N_3323;
    
    wire n3301, \FRAME_MATCHER.rx_data_ready_prev , n31226, n36056, 
        n35975, n10_adj_3920, n31124, n35910, n18019, n18018;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n17989, n1395, n35654, n35898, n17988, n1254, n35648, 
        n2_adj_3921, n2_adj_3922, n28483, n36032, n20, n36023, n19_adj_3923, 
        n18017, n18016, n21, n31288, n35577, n1173, n22, n16993, 
        n16_adj_3924, n24, n20_adj_3925, n16487, n14_adj_3926, n18_adj_3927, 
        n16_adj_3928, n20_adj_3929, n25693, n25503, n38973, n25687, 
        n35365, n17124, n12_adj_3930, n36731, n2783, n3_adj_3931, 
        n3_adj_3932, n3_adj_3933, n3_adj_3934, n3_adj_3935, n3_adj_3936, 
        n3_adj_3937, n3_adj_3938, n3_adj_3939, n3_adj_3940, n3_adj_3941, 
        n3_adj_3942, n3_adj_3943, n18015, n18014, n3_adj_3944, n18013, 
        n3_adj_3945, n3_adj_3946, n3_adj_3947, n3_adj_3948, n3_adj_3949, 
        n3_adj_3950, n3_adj_3951, n3_adj_3952, n3_adj_3953, n3_adj_3954, 
        n3_adj_3955, n3_adj_3956, n3_adj_3957, n3_adj_3958, n3_adj_3959, 
        n3_adj_3960, n17987, n2_adj_3961, n28482, n17986;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n2_adj_3962, n28481, n2_adj_3963, n28480, n15879, n99, 
        n96, n31898, tx_transmit_N_3220, n25775, n8_adj_3964, n2_adj_3965, 
        n28479, n2_adj_3966, n28478, n44226, n28518, n2_adj_3967, 
        n28477, n28517, n3_adj_3968, n2_adj_3969, n28476, n28516, 
        n17985, n28515, n17984, n17983, n17982, n2_adj_3970, n28475, 
        n2_adj_3971, n28474, n2_adj_3972, n28473, n2_adj_3973, n28472, 
        n28514, n28513, n9, n2_adj_3974, n28471, n28512, n17981, 
        n2_adj_3975, n28470, n17980, n37242, n35607, n35519, n35468, 
        Kp_23__N_839, n35610, n18_adj_3976, n39061, n30_adj_3977, 
        n5_c, n22_adj_3978, n4_adj_3979, n24_adj_3980, n35829, n32_adj_3981, 
        n27_adj_3982, n39063;
    wire [31:0]\FRAME_MATCHER.state_31__N_2490 ;
    
    wire n6_adj_3983, n161, n38135, n17807, n17979, n13_adj_3984, 
        n10_adj_3985, n14_adj_3986, n14_adj_3987, n15, n8_adj_3988, 
        n12_adj_3989, n35256, n91, n12_adj_3990, n10_adj_3991, n14_adj_3992, 
        n13455, Kp_23__N_760, n16514, n35645, n35966, n35892, n36071, 
        n35808, n74, n35814, n35494, n35639, n73, n16137, n35574, 
        n35996, n71, n48, Kp_23__N_1406, n35984, n70, n36059, 
        n80, n16630, n35987, n36098, n35491, n78, n16276, n76, 
        n36062, n16371, Kp_23__N_893, n77, n35737, n35568, n35633, 
        n35836, n75, n72, n86, n16919, n68, n16802, n85, n87, 
        n36065, n35500, n35843, n35820, n31231, n16496, n32001, 
        n35719, n36095, n16076, n35922, n31488, n31114, n35923, 
        n35963, n6_adj_3993, n31202, n63_c, n63_adj_3994, n41084, 
        n25745, n15862, n10_adj_3997, n15974, n36328, n38180, n15729, 
        n4_adj_3998, n42, n35990, n16173, n16592, n35856, Kp_23__N_1418, 
        n36020, n31987, n35733, n35928, n35805, n35969, n16197, 
        n16564, n40, n41, n39, n38, n37, n48_adj_3999, n43, 
        n35531, n35527, n6_adj_4000, n35497, n35787, n6_adj_4001, 
        n35839, n36107, n14_adj_4002, n36053, n31210, n15_adj_4003, 
        n36092, n35676, n6_adj_4004, n16306, n16557, n31156, n35772, 
        n35775, n31200, n14_adj_4005, n14_adj_4006, n15971, n15_adj_4007, 
        n15_adj_4008, n35630, n36050, n31964, n12_adj_4009, n35956, 
        n32016, n35999, n36074, n10_adj_4010, n6_adj_4011, n15769, 
        n16_adj_4012, n17_adj_4013, n6_adj_4014, n6_adj_4015, n35601, 
        n35688, n35481, n16192, n36967, n35901, n16808, n11, n35664, 
        n15859, n10_adj_4016, n6_adj_4017, n16748, n36101, n35762, 
        n35723, Kp_23__N_847, n35475, n31100, n31224, n31190, n4_adj_4018, 
        n16974, n31979, n16_adj_4019, n17_adj_4020, n31222, n35589, 
        n10_adj_4021, n35667, n35625, n16218, n12_adj_4022, n35798, 
        n16971, n31959, n35741, n12_adj_4023, n14_adj_4024, n15856, 
        n18_adj_4025, n20_adj_4026, n15_adj_4027, n16142, n16624, 
        Kp_23__N_946, n16532, n35972, n10_adj_4028, n16567, n16916, 
        n35595, n6_adj_4029, n35713, n35642, n16_adj_4030, n17_adj_4031, 
        n10_adj_4032, n31170, n35895, n15_adj_4033, n14_adj_4034, 
        n18_adj_4035, n24_adj_4036, n22_adj_4037, n26, n35888, n35801, 
        n16784, n35583, n10_adj_4038, n35784, n20_adj_4039, n19_adj_4040, 
        n39097, n35744, n18_adj_4041, n20_adj_4042, n36017, n15_adj_4043, 
        n35535, n35564, n24660, n25346, n35622, n35875, n20_adj_4044, 
        n35925, n19_adj_4045, n21_adj_4046, n37788, n35853, n12_adj_4047, 
        n15_adj_4048, n8_adj_4049, n35943, n6_adj_4050, n35884, n10_adj_4051, 
        n10_adj_4052, n16824, n24_adj_4053, n35730, n10_adj_4054, 
        n34, n25, n32_adj_4055, n36005, n35859, n31_adj_4056, n35, 
        n31962, n37_adj_4057, n37969, n10_adj_4058, n31794, n14_adj_4059, 
        n15_adj_4060, n15_adj_4061, n36026, n14_adj_4062, n35694, 
        n37640, n10_adj_4063, n37446, n18_adj_4064, n16_adj_4065, 
        n20_adj_4066, n35661, n19_adj_4067, n44816, n36896, n20_adj_4068, 
        n14_adj_4069, n15_adj_4070, n16_adj_4071, n17_adj_4072, n37311, 
        n4_adj_4073, n37705, n21_adj_4074, n12_adj_4075, n37238, n39065, 
        n37275, n27_adj_4076, n6_adj_4077, n36860, n18_adj_4078, n26_adj_4079, 
        n30_adj_4080, n17_adj_4081, n31_adj_4082, n104, n39023, n2_adj_4083, 
        n2_adj_4084, n2_adj_4085, n2_adj_4086, n2_adj_4087, n2_adj_4088, 
        n2_adj_4089, n2_adj_4090, n2_adj_4091, n2_adj_4092, n2_adj_4093, 
        n37040, n37659, n37704, n37148, n35540, n37006, n37420, 
        n35698, n37234, n35652, n34722, n34894, n35400, n34724, 
        n7_adj_4094, n8_adj_4095, n35403, n34798, n35397, n34796, 
        n35406, n34794, n35391, n34792, n35390, n34720, n35392, 
        n34790, n35407, n34788, n35398, n34786, n35404, n34784, 
        n35401, n34782, n35409, n34780, n35394, n34778, n7_adj_4096, 
        n8_adj_4097, n35395, n34776, n7_adj_4098, n8_adj_4099, n35393, 
        n34774, n24653, n25478, n35408, n34772, n7_adj_4100, n8_adj_4101, 
        n37102, n34680, n7_adj_4102, n8_adj_4103, n35399, n34732, 
        n35402, n34770, n35396, n34768, n35405, n34766, n35389, 
        n25470, n14_adj_4104, n28491, n28492, n18012, n28500, n28499, 
        n28498, n44382, n44376, n44379, n44370, n44373, n18011, 
        n18010, n18009, n18008, n18007, n18006, n18005, n18004, 
        n18003, n18002, n18001, n18000, n17291, n36732, n38154, 
        n44364, n28497, n28496, n44367, n44358, n44361, n28495, 
        n17999, Kp_23__N_1427, n4377, n28494, n8_adj_4107, n35439, 
        n17992, n28493, n17993, n17998, n17997, n17996, n17994, 
        n28490, n16348, n17995, n6_adj_4108, n31967, n37462, n35383, 
        n4_adj_4109, n35448, n131, n13197, n8_adj_4110, n24972, 
        n8_adj_4111, n12_adj_4112, n16_adj_4113, n2106, n14_adj_4114, 
        n35703, n16477, n32012, n30900, n16_adj_4115, n17_adj_4116, 
        n39270, n39271, n39274, n39273, n6_adj_4117, n35552, n35759, 
        n35867, n6_adj_4118, n35386, n38_adj_4119, n13142, n7_adj_4120, 
        n8_adj_4121, n8_adj_4122, n44352, n8_adj_4123, n44355, n44346, 
        n44349, n39185, n39184, n44340, n44343, n44334, n39182, 
        n39181, n39179, n44259, n44328, n44331, n44322, n44325, 
        n39209, n39208, n44316, n39212, n39211, n44319, n44310, 
        n44313, n44304, n44307, n8_adj_4124, n1_c, n44298, n44301, 
        n44292, n44295, n44286, n44289, n24745, n44280, n31208, 
        n19450, n31_adj_4125, n12969, n8_adj_4126, n28_adj_4127, n26_adj_4128, 
        n27_adj_4129, n25_adj_4130, n44283, n4_adj_4131, n38182, n36130, 
        n44274, n44277, n36104, n19_adj_4132, n41676, n5_adj_4133, 
        n39229, n39230, n39183, n19_adj_4134, n42389, n5_adj_4135, 
        n39226, n39227, n39180, n19_adj_4136, n39223, n41668, n5_adj_4137, 
        n39224, n39177, n19_adj_4138, n6_adj_4139, n5_adj_4140, n39220, 
        n39221, n39210, n19_adj_4141, n6_adj_4142, n5_adj_4143, n39217, 
        n39218, n39207, n39250, n44262, n19_adj_4144, n39193, n44265, 
        n42800, n39194, n43073, n44256, n19_adj_4145, n39190, n44253, 
        n42804, n39191, n43071, n44250, n43489, n44244, n35388, 
        n35449, n4_adj_4146, n7_adj_4147, n31228, n32092, n10_adj_4148, 
        n15497, n35561, n35539, n31140, n35817, n35553, n32094, 
        n35555, n35598, n35811, n14_adj_4149, n15_adj_4150, n37421, 
        n16723, n22_adj_4151, n21_adj_4152, n14_adj_4153, n23, n13_adj_4154, 
        n15_adj_4155, n52, n50, n51, n49, n46, n48_adj_4156, n47, 
        n58, n53, n15_adj_4157, n35616, n10_adj_4158;
    
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18036));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35619));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n35619), .I1(n15522), .I2(n31104), .I3(n35673), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_41_21 (.CI(n28488), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n28489));
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18035));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18034));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18033));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18032));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18031));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18030));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[15] [2]), .I1(n10), .I2(\data_out_frame[19] [4]), 
            .I3(GND_net), .O(n37402));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_22_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n28489), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_22_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18029));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18028));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18027));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n17991));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n17973));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[17] [2]), .I1(n15522), 
            .I2(GND_net), .I3(GND_net), .O(n31150));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17902));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n17972));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_865 (.I0(\data_out_frame[19] [3]), .I1(n35934), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[16] [7]), 
            .O(n10_adj_3893));
    defparam i4_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3894), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18026));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18025));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18023));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_20_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n28487), .O(n2_adj_3895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_20_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18022));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_866 (.I0(n7_c), .I1(\data_out_frame[17] [0]), .I2(n35954), 
            .I3(n35727), .O(n37444));
    defparam i4_4_lut_adj_866.LUT_INIT = 16'h9669;
    SB_CARRY add_41_20 (.CI(n28487), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n28488));
    SB_LUT4 i1_2_lut_adj_867 (.I0(\data_out_frame[15] [0]), .I1(n1640), 
            .I2(GND_net), .I3(GND_net), .O(n35673));
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(n36002), .I1(n36077), .I2(\data_out_frame[10] [3]), 
            .I3(n35679), .O(n12));   // verilog/coms.v(83[17:28])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[14] [7]), .I1(n12), .I2(n36080), 
            .I3(\data_out_frame[14] [6]), .O(n15522));   // verilog/coms.v(83[17:28])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[13] [4]), .I1(n16234), .I2(n35904), 
            .I3(n35670), .O(n35765));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(n35765), .I3(GND_net), .O(n35947));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_868 (.I0(n15522), .I1(n31973), .I2(n35954), .I3(n31142), 
            .O(n12_adj_3896));
    defparam i5_4_lut_adj_868.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n17933));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_869 (.I0(n16238), .I1(n12_adj_3896), .I2(n35947), 
            .I3(n31164), .O(n36742));
    defparam i6_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n17932));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17901));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n17931));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n17930));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n17929));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n17928));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n17927));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_870 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[12] [6]), 
            .I2(n35881), .I3(n1117), .O(n16_c));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17900));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[10] [4]), .I1(n35613), .I2(n36011), 
            .I3(n16898), .O(n17));   // verilog/coms.v(71[16:42])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_out_frame[13] [1]), .I2(n16_c), 
            .I3(n16042), .O(n1640));   // verilog/coms.v(71[16:42])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_871 (.I0(\data_out_frame[6] [6]), .I1(n35918), 
            .I2(n35547), .I3(\data_out_frame[11] [0]), .O(n36038));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_872 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n35781));
    defparam i2_3_lut_adj_872.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_873 (.I0(\data_out_frame[13] [2]), .I1(n36038), 
            .I2(\data_out_frame[9] [0]), .I3(\data_out_frame[4][1] ), .O(n10_adj_3897));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_874 (.I0(n35864), .I1(n10_adj_3897), .I2(\data_out_frame[4][0] ), 
            .I3(GND_net), .O(n35826));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n18153));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n18154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n18155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n18156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n18157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n18158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n18142));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n18143));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n17515));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n17548));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n17554));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n17551));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n17560));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n17557));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n17563));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n18159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n18160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n18144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n18145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n18146));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n18147));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n18148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n18149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n18150));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n18151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n18152));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n18140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n18141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n18138));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n18139));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_875 (.I0(\data_out_frame[12] [7]), .I1(n35993), 
            .I2(n35826), .I3(n35781), .O(n30880));
    defparam i3_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n17926));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n17925));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), .C(clk32MHz), 
            .E(VCC_net), .D(n18108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17899));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18037));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18038));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18042));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17898));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17897));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17896));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17895));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n44420));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n44421));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n17971));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n17970));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n17969));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n17968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n17967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n17966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17894));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17893));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17892));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18046));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18047));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17891));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18043));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18044));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18045));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17890));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17889));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17888));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17887));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17886));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17885));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17884));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17883));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17882));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17881));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17880));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17879));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n17965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17878));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17877));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17876));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17875));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n17964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17874));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17873));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_876 (.I0(n16403), .I1(n16698), .I2(\data_out_frame[12] [1]), 
            .I3(GND_net), .O(n37377));
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17872));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17871));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17870));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[14] [5]), 
            .I2(n15502), .I3(n18), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n17924));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n17869));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n17923));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n17868));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n17990));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n17867));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i11_4_lut (.I0(n35781), .I1(\data_out_frame[14] [1]), .I2(n37377), 
            .I3(n36038), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n36008), .I1(n35823), .I2(n35870), .I3(n35542), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n36014), .I1(n36044), .I2(n35504), .I3(n35937), 
            .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17866));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n31973));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n17922));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1073_2_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1829));   // verilog/coms.v(69[16:27])
    defparam i1073_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_877 (.I0(\data_out_frame[17] [1]), .I1(n31973), 
            .I2(n35700), .I3(n30880), .O(n35934));
    defparam i3_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_19_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n28486), .O(n2_adj_3898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_19 (.CI(n28486), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n28487));
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n17921));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_878 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_c));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_878.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_879 (.I0(\data_out_frame[5] [0]), .I1(n35571), 
            .I2(\data_out_frame[6] [4]), .I3(n6_c), .O(n35670));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n17920));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_880 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[4][2] ), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n35613));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_881 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36035));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_882 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35918));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_882.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_883 (.I0(n36035), .I1(n35613), .I2(\data_out_frame[7] [0]), 
            .I3(n36068), .O(n10_adj_3899));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n36008));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_out_frame[13] [3]), .I1(n15502), 
            .I2(GND_net), .I3(GND_net), .O(n35462));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_886 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35878));
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_887 (.I0(n35878), .I1(n35462), .I2(\data_out_frame[9] [2]), 
            .I3(n36008), .O(n10_adj_3900));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_888 (.I0(n35670), .I1(n10_adj_3900), .I2(\data_out_frame[7] [0]), 
            .I3(GND_net), .O(n31109));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_888.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_889 (.I0(n36011), .I1(n16898), .I2(\data_out_frame[10] [7]), 
            .I3(\data_out_frame[8] [5]), .O(n35993));   // verilog/coms.v(95[12:26])
    defparam i3_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_890 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[4][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n35571));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16022));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n17919));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n17918));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n17917));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17916));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_892 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n35978));
    defparam i2_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35547));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17915));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out_frame[4][2] ), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n36077));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17914));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17913));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17912));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10_4_lut_adj_895 (.I0(n36077), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[11] [1]), .I3(n35547), .O(n28_adj_3901));
    defparam i10_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i36631_3_lut (.I0(n16394), .I1(n15489), .I2(n35691), .I3(GND_net), 
            .O(n43485));
    defparam i36631_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17911));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17910));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17909));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17908));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12_4_lut_adj_896 (.I0(n16052), .I1(n36068), .I2(n43485), 
            .I3(n35978), .O(n30_adj_3902));
    defparam i12_4_lut_adj_896.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17907));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n17906));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17905));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13_4_lut_adj_897 (.I0(n35684), .I1(n35478), .I2(n35571), 
            .I3(\data_out_frame[11] [5]), .O(n31));
    defparam i13_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_898 (.I0(n35907), .I1(n35993), .I2(n31090), 
            .I3(n35604), .O(n29_adj_3903));
    defparam i11_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n29_adj_3903), .I1(n31), .I2(n30_adj_3902), 
            .I3(n32), .O(n35753));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n36014));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35881));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_901 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[4][0] ), .I3(n16022), .O(n36080));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_902 (.I0(n36080), .I1(n35657), .I2(GND_net), 
            .I3(GND_net), .O(n8));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_903 (.I0(n35881), .I1(n36014), .I2(\data_out_frame[12] [7]), 
            .I3(n35753), .O(n12_adj_3904));   // verilog/coms.v(83[17:70])
    defparam i5_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17904));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17865));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(n12_adj_3904), .I3(n8), .O(n35937));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_904 (.I0(n16042), .I1(n35937), .I2(\data_out_frame[8] [5]), 
            .I3(n1048), .O(n12_adj_3905));
    defparam i5_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_905 (.I0(\data_out_frame[12] [5]), .I1(n12_adj_3905), 
            .I2(\data_out_frame[15] [1]), .I3(n35753), .O(n32044));
    defparam i6_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_906 (.I0(n31109), .I1(\data_out_frame[15] [4]), 
            .I2(n8_adj_3906), .I3(\data_out_frame[15] [3]), .O(n35749));
    defparam i1_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_907 (.I0(n35749), .I1(n32044), .I2(GND_net), 
            .I3(GND_net), .O(n35954));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n16238), .I1(n31802), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[19] [2]), .I1(n35934), .I2(n1829), 
            .I3(n4_c), .O(n35727));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_909 (.I0(n35727), .I1(n36047), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3907));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_910 (.I0(n31168), .I1(\data_out_frame[19] [1]), 
            .I2(n35954), .I3(n6_adj_3907), .O(n37260));
    defparam i4_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i292_2_lut (.I0(\data_out_frame[4][1] ), .I1(\data_out_frame[4][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1048));   // verilog/coms.v(70[16:27])
    defparam i292_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_911 (.I0(\data_out_frame[10] [4]), .I1(n35657), 
            .I2(\data_out_frame[12] [5]), .I3(\data_out_frame[14] [6]), 
            .O(n35504));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_912 (.I0(\data_out_frame[6] [2]), .I1(n35846), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[12] [4]), 
            .O(n36002));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_913 (.I0(n16094), .I1(n36002), .I2(n35504), .I3(n1048), 
            .O(n16238));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_914 (.I0(\data_out_frame[19] [0]), .I1(n32004), 
            .I2(\data_out_frame[19] [1]), .I3(GND_net), .O(n35756));
    defparam i2_3_lut_adj_914.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_915 (.I0(n30877), .I1(n16238), .I2(GND_net), 
            .I3(GND_net), .O(n31168));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_916 (.I0(n35940), .I1(n31164), .I2(\data_out_frame[16] [6]), 
            .I3(n31168), .O(n14));
    defparam i6_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_917 (.I0(\data_out_frame[16] [7]), .I1(n14), .I2(n10_adj_3908), 
            .I3(\data_out_frame[16] [4]), .O(n36725));
    defparam i7_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16698));
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_919 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35691));
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_920 (.I0(n16535), .I1(n35558), .I2(n15489), .I3(n35513), 
            .O(n12_adj_3909));   // verilog/coms.v(95[12:26])
    defparam i4_4_lut_adj_920.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_921 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[8] [2]), 
            .I2(n35691), .I3(n16698), .O(n13));   // verilog/coms.v(95[12:26])
    defparam i5_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_922 (.I0(n13), .I1(n35913), .I2(n12_adj_3909), 
            .I3(n16711), .O(n31164));   // verilog/coms.v(95[12:26])
    defparam i7_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_923 (.I0(\data_out_frame[18] [5]), .I1(n31684), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n35484));
    defparam i2_3_lut_adj_923.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_924 (.I0(n35484), .I1(\data_out_frame[19] [0]), 
            .I2(n32079), .I3(GND_net), .O(n35960));
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_925 (.I0(\data_out_frame[16] [6]), .I1(n31802), 
            .I2(n35960), .I3(n6_adj_3910), .O(n37263));
    defparam i4_4_lut_adj_925.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17864));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17863));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17862));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17861));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17860));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17859));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n17963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17858));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17857));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17856));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17855));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17854));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17853));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17852));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n17851));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n17850));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n17849));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n17848));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i32351_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n39251), .I3(n39249), .O(n39204));
    defparam i32351_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n17962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n17847));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n17846));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n17845));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17844));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17843));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17842));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17841));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17840));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17839));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17838));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17837));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_18_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n28485), .O(n2_adj_3911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35657));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35833));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_CARRY add_41_18 (.CI(n28485), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n28486));
    SB_LUT4 add_41_17_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n28484), .O(n2_adj_3912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_928 (.I0(n35487), .I1(n35833), .I2(\data_out_frame[12] [3]), 
            .I3(\data_out_frame[5] [7]), .O(n12_adj_3913));   // verilog/coms.v(83[17:28])
    defparam i5_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_929 (.I0(\data_out_frame[12] [2]), .I1(n12_adj_3913), 
            .I2(n35846), .I3(n31090), .O(n31802));   // verilog/coms.v(83[17:28])
    defparam i6_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_930 (.I0(n15489), .I1(n12_adj_3914), .I2(n36029), 
            .I3(n16898), .O(n16_adj_3915));
    defparam i6_4_lut_adj_930.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_931 (.I0(\data_out_frame[14] [3]), .I1(n35907), 
            .I2(n36083), .I3(\data_out_frame[12] [1]), .O(n17_adj_3916));
    defparam i7_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18021));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_932 (.I0(n17_adj_3916), .I1(\data_out_frame[12] [2]), 
            .I2(n16_adj_3915), .I3(n14104), .O(n30877));
    defparam i9_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_933 (.I0(\data_out_frame[7] [0]), .I1(n35580), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [2]), .O(n35904));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n36089));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_935 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35950));
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_936 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35465));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_LUT4 i32348_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n39242), .I3(n39240), .O(n39201));
    defparam i32348_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i32379_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39232));
    defparam i32379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32334_4_lut (.I0(n19), .I1(\data_out_frame[22] [0]), .I2(byte_transmit_counter[1]), 
            .I3(\byte_transmit_counter[0] ), .O(n39187));
    defparam i32334_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32380_4_lut (.I0(n39232), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n39233));
    defparam i32380_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i32378_3_lut (.I0(\data_out_frame[4][0] ), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39231));
    defparam i32378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35952_3_lut (.I0(n44385), .I1(n44247), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n42806));
    defparam i35952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_937 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [1]), 
            .I2(n32007), .I3(GND_net), .O(n36937));
    defparam i2_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_LUT4 i32335_3_lut (.I0(n44337), .I1(n39187), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39188));
    defparam i32335_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18020));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_938 (.I0(n36089), .I1(n35507), .I2(n35904), .I3(\data_out_frame[16]_c [2]), 
            .O(n14_adj_3917));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i36645_4_lut (.I0(\data_out_frame[13] [7]), .I1(n36937), .I2(n8_adj_3918), 
            .I3(n1238), .O(n43499));
    defparam i36645_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_939 (.I0(n43499), .I1(n14_adj_3917), .I2(n10_adj_3919), 
            .I3(n35850), .O(n16704));   // verilog/coms.v(69[16:27])
    defparam i7_4_lut_adj_939.LUT_INIT = 16'h9669;
    SB_LUT4 i36209_3_lut (.I0(n39198), .I1(n42806), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n43063));   // verilog/coms.v(104[34:55])
    defparam i36209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_out_frame[20] [7]), .I1(n30877), 
            .I2(GND_net), .I3(GND_net), .O(n35778));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i36210_4_lut (.I0(n43063), .I1(n39188), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam i36210_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_3_lut_adj_941 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n35823));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_941.LUT_INIT = 16'h9696;
    SB_DFFSR tx_transmit_3205 (.Q(r_SM_Main_2__N_3323[0]), .C(clk32MHz), 
            .D(n3299[0]), .R(n3301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3206  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_942 (.I0(n35823), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n31226));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_942.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_943 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [2]), 
            .I2(n36056), .I3(n35975), .O(n10_adj_3920));   // verilog/coms.v(95[12:26])
    defparam i4_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_944 (.I0(n31124), .I1(n10_adj_3920), .I2(n35910), 
            .I3(GND_net), .O(n32007));   // verilog/coms.v(95[12:26])
    defparam i5_3_lut_adj_944.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_945 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35558));   // verilog/coms.v(95[12:26])
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_946 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35580));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_946.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_947 (.I0(\data_out_frame[9] [1]), .I1(n35580), 
            .I2(\data_out_frame[9] [4]), .I3(n16394), .O(n16052));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16898));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18019));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18018));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n17989));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17836));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35679));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_out_frame[9] [5]), .I1(n16052), 
            .I2(GND_net), .I3(GND_net), .O(n1395));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_out_frame[5] [4]), .I1(n35654), 
            .I2(GND_net), .I3(GND_net), .O(n15489));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16403));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35898));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35604));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35684));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n17988));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16394));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i498_2_lut (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1254));   // verilog/coms.v(83[17:28])
    defparam i498_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i364_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/coms.v(83[17:28])
    defparam i364_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35648));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17835));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n17974));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n17961));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_21_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n28488), .O(n2_adj_3921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_958 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[7] [3]), .O(n1238));
    defparam i3_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_959 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16094));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h6666;
    SB_CARRY add_41_17 (.CI(n28484), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n28485));
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35850));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 add_41_16_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n28483), .O(n2_adj_3922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_961 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n35864));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_962 (.I0(\data_out_frame[6] [7]), .I1(n35513), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n36032));
    defparam i2_3_lut_adj_962.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_out_frame[4][0] ), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35542));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(n35542), .I1(n36032), .I2(\data_out_frame[7] [0]), 
            .I3(n35864), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_964 (.I0(n35850), .I1(\data_out_frame[4][2] ), 
            .I2(n16094), .I3(n36023), .O(n19_adj_3923));
    defparam i7_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18017));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18016));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_965 (.I0(n35648), .I1(n1117), .I2(\data_out_frame[6] [0]), 
            .I3(n1254), .O(n21));
    defparam i9_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_966 (.I0(n31288), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36083));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_967 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[14] [3]), .I3(\data_out_frame[14] [2]), 
            .O(n35870));
    defparam i3_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_968 (.I0(n35898), .I1(n16403), .I2(n35577), .I3(n1173), 
            .O(n22));   // verilog/coms.v(95[12:26])
    defparam i9_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_969 (.I0(n16993), .I1(n22), .I2(n16_adj_3924), 
            .I3(n35870), .O(n24));   // verilog/coms.v(95[12:26])
    defparam i11_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_970 (.I0(n35910), .I1(n24), .I2(n20_adj_3925), 
            .I3(n35975), .O(n32079));   // verilog/coms.v(95[12:26])
    defparam i12_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_971 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16487));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_972 (.I0(n32079), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35940));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h9999;
    SB_LUT4 i3_2_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[16][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3926));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17834));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_973 (.I0(n15489), .I1(n14_adj_3926), .I2(n35558), 
            .I3(n32007), .O(n18_adj_3927));
    defparam i7_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3928));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_974 (.I0(n31226), .I1(n18_adj_3927), .I2(\data_out_frame[14] [2]), 
            .I3(n35898), .O(n20_adj_3929));
    defparam i9_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_975 (.I0(n35654), .I1(n20_adj_3929), .I2(n16_adj_3928), 
            .I3(n35465), .O(n31684));
    defparam i10_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i32193_2_lut (.I0(n25693), .I1(n25503), .I2(GND_net), .I3(GND_net), 
            .O(n38973));
    defparam i32193_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_976 (.I0(n38973), .I1(n25687), .I2(n35365), .I3(\FRAME_MATCHER.state [1]), 
            .O(n17124));
    defparam i3_4_lut_adj_976.LUT_INIT = 16'h0010;
    SB_LUT4 i5_4_lut_adj_977 (.I0(\data_out_frame[20] [6]), .I1(n35778), 
            .I2(\data_out_frame[16][5] ), .I3(n16704), .O(n12_adj_3930));
    defparam i5_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17833));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_978 (.I0(n31684), .I1(n12_adj_3930), .I2(n35940), 
            .I3(n16487), .O(n36731));
    defparam i6_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 select_353_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3931));
    defparam select_353_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3932));
    defparam select_353_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3933));
    defparam select_353_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3934));
    defparam select_353_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3935));
    defparam select_353_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3936));
    defparam select_353_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3937));
    defparam select_353_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3938));
    defparam select_353_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3939));
    defparam select_353_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3940));
    defparam select_353_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3941));
    defparam select_353_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3942));
    defparam select_353_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3943));
    defparam select_353_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18015));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18014));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_353_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3944));
    defparam select_353_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18013));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_353_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3945));
    defparam select_353_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3946));
    defparam select_353_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3947));
    defparam select_353_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3948));
    defparam select_353_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3949));
    defparam select_353_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3950));
    defparam select_353_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3951));
    defparam select_353_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3952));
    defparam select_353_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3953));
    defparam select_353_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3954));
    defparam select_353_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17832));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_353_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3955));
    defparam select_353_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3956));
    defparam select_353_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3957));
    defparam select_353_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3958));
    defparam select_353_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3959));
    defparam select_353_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_353_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3960));
    defparam select_353_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n17987));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_16 (.CI(n28483), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n28484));
    SB_LUT4 add_41_15_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n28482), .O(n2_adj_3961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_15_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17831));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_15 (.CI(n28482), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n28483));
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n17986));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_14_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n28481), .O(n2_adj_3962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_14 (.CI(n28481), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n28482));
    SB_LUT4 add_41_13_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n28480), .O(n2_adj_3963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_13 (.CI(n28480), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n28481));
    SB_LUT4 i1_2_lut_adj_979 (.I0(n15879), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n99));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_979.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_980 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n96));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_LUT4 i36652_2_lut (.I0(n31898), .I1(n15879), .I2(GND_net), .I3(GND_net), 
            .O(n3301));
    defparam i36652_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 select_353_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_353_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_775_i1_4_lut (.I0(tx_transmit_N_3220), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n25775), .I3(n8_adj_3964), .O(n3299[0]));   // verilog/coms.v(144[4] 288[11])
    defparam mux_775_i1_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 add_41_12_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n28479), .O(n2_adj_3965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_12 (.CI(n28479), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n28480));
    SB_LUT4 add_41_11_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n28478), .O(n2_adj_3966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3279_9_lut (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[7]), 
            .I2(n44226), .I3(n28518), .O(n17513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_41_11 (.CI(n28478), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n28479));
    SB_LUT4 add_41_10_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n28477), .O(n2_adj_3967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3279_8_lut (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[6]), 
            .I2(n44226), .I3(n28517), .O(n17546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 select_353_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2783), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3968));
    defparam select_353_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_41_10 (.CI(n28477), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n28478));
    SB_CARRY add_3279_8 (.CI(n28517), .I0(byte_transmit_counter[6]), .I1(n44226), 
            .CO(n28518));
    SB_LUT4 add_41_9_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n28476), .O(n2_adj_3969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3279_7_lut (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[5]), 
            .I2(n44226), .I3(n28516), .O(n17549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_7_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n17985));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_3279_7 (.CI(n28516), .I0(byte_transmit_counter[5]), .I1(n44226), 
            .CO(n28517));
    SB_LUT4 add_3279_6_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[4]), 
            .I2(n44226), .I3(n28515), .O(n17552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_41_9 (.CI(n28476), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n28477));
    SB_CARRY add_3279_6 (.CI(n28515), .I0(byte_transmit_counter[4]), .I1(n44226), 
            .CO(n28516));
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n17984));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n17960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n17983));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n17982));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n17959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n17958));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_8_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n28475), .O(n2_adj_3970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_8 (.CI(n28475), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n28476));
    SB_LUT4 add_41_7_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n28474), .O(n2_adj_3971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_7 (.CI(n28474), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n28475));
    SB_LUT4 add_41_6_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n28473), .O(n2_adj_3972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_6 (.CI(n28473), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n28474));
    SB_LUT4 add_41_5_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n28472), .O(n2_adj_3973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17830));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_3279_5_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[3]), 
            .I2(n44226), .I3(n28514), .O(n17555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_3279_5 (.CI(n28514), .I0(byte_transmit_counter[3]), .I1(n44226), 
            .CO(n28515));
    SB_CARRY add_41_5 (.CI(n28472), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n28473));
    SB_LUT4 add_3279_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[2]), 
            .I2(n44226), .I3(n28513), .O(n17558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 equal_122_i9_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/coms.v(151[7:23])
    defparam equal_122_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_41_4_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n28471), .O(n2_adj_3974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3279_4 (.CI(n28513), .I0(byte_transmit_counter[2]), .I1(n44226), 
            .CO(n28514));
    SB_CARRY add_41_4 (.CI(n28471), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n28472));
    SB_LUT4 add_3279_3_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[1]), 
            .I2(n44226), .I3(n28512), .O(n17561)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_3279_3 (.CI(n28512), .I0(byte_transmit_counter[1]), .I1(n44226), 
            .CO(n28513));
    SB_LUT4 add_3279_2_lut (.I0(GND_net), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3220), .I3(GND_net), .O(n7821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3220), .CO(n28512));
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n17981));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_3_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n28470), .O(n2_adj_3975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17829));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17828));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17827));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17826));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n17980));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17825));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17824));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17823));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17822));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17821));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17820));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17819));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n15879), .I3(\FRAME_MATCHER.state[0] ), .O(n37242));   // verilog/coms.v(126[12] 289[6])
    defparam i2_4_lut_4_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35607));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_982 (.I0(\data_in_frame[0] [5]), .I1(n35607), .I2(n35519), 
            .I3(n35468), .O(Kp_23__N_839));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_983 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_839), 
            .I2(GND_net), .I3(GND_net), .O(n35610));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n18_adj_3976));
    defparam i1_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i13_4_lut_adj_984 (.I0(n39061), .I1(\data_in_frame[2] [0]), 
            .I2(n18_adj_3976), .I3(n35610), .O(n30_adj_3977));
    defparam i13_4_lut_adj_984.LUT_INIT = 16'h4010;
    SB_LUT4 i5_3_lut_adj_985 (.I0(n5_c), .I1(Kp_23__N_839), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22_adj_3978));
    defparam i5_3_lut_adj_985.LUT_INIT = 16'h1414;
    SB_LUT4 i15_4_lut (.I0(n4_adj_3979), .I1(n30_adj_3977), .I2(n24_adj_3980), 
            .I3(n35829), .O(n32_adj_3981));
    defparam i15_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i10_4_lut_adj_986 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [6]), .O(n27_adj_3982));
    defparam i10_4_lut_adj_986.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_987 (.I0(n27_adj_3982), .I1(n32_adj_3981), .I2(n39063), 
            .I3(n22_adj_3978), .O(\FRAME_MATCHER.state_31__N_2490 [3]));
    defparam i16_4_lut_adj_987.LUT_INIT = 16'h0800;
    SB_LUT4 i2_2_lut (.I0(n15879), .I1(\FRAME_MATCHER.state_31__N_2490 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3983));   // verilog/coms.v(126[12] 289[6])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(150[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_988 (.I0(n38135), .I1(n6_adj_3983), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n35365), .O(n13293));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_988.LUT_INIT = 16'hc080;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17818));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17817));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17816));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17815));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17814));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17813));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17812));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17811));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16][5] ), .C(clk32MHz), 
           .D(n17810));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17809));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16][3] ), .C(clk32MHz), 
           .D(n17808));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16]_c [2]), .C(clk32MHz), 
           .D(n17807));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16][1] ), .C(clk32MHz), 
           .D(n17806));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16][0] ), .C(clk32MHz), 
           .D(n17805));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17804));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17803));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17802));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17801));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17800));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17799));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17798));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17797));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17796));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17795));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17794));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17793));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17792));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17791));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17790));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17789));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17788));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17787));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n17979));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n17978));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17786));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17785));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17784));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n17977));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n17976));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17783));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17782));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17781));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17780));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17779));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17778));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17777));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17776));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17775));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17774));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17773));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17772));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17771));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17770));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17769));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17768));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17767));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17766));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17765));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17764));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17763));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17762));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17761));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_3 (.CI(n28470), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n28471));
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17760));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17759));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17758));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17757));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17756));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i32345_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n39233), .I3(n39231), .O(n39198));
    defparam i32345_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_41_2_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_3894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n28470));
    SB_LUT4 i1_3_lut_adj_989 (.I0(n15879), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n13_adj_3984));
    defparam i1_3_lut_adj_989.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_adj_990 (.I0(\FRAME_MATCHER.i_31__N_2390 ), .I1(n13_adj_3984), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n2086));
    defparam i2_3_lut_adj_990.LUT_INIT = 16'habab;
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17755));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_2_lut_adj_991 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3985));
    defparam i2_2_lut_adj_991.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_992 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [11]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [15]), 
            .O(n14_adj_3986));
    defparam i6_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_993 (.I0(\FRAME_MATCHER.state [14]), .I1(n14_adj_3986), 
            .I2(n10_adj_3985), .I3(\FRAME_MATCHER.state [9]), .O(n25687));
    defparam i7_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_994 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [28]), 
            .I2(\FRAME_MATCHER.state [24]), .I3(GND_net), .O(n14_adj_3987));
    defparam i5_3_lut_adj_994.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17754));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17753));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17752));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_995 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [18]), 
            .O(n15));
    defparam i6_4_lut_adj_995.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17751));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_996 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3988));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17750));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_997 (.I0(\FRAME_MATCHER.state [25]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(\FRAME_MATCHER.state [29]), 
            .O(n12_adj_3989));
    defparam i5_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17749));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_4_lut_adj_998 (.I0(n15), .I1(\FRAME_MATCHER.state [16]), 
            .I2(n14_adj_3987), .I3(\FRAME_MATCHER.state [19]), .O(n35256));
    defparam i8_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17748));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut_adj_999 (.I0(\FRAME_MATCHER.state [27]), .I1(n35256), 
            .I2(n12_adj_3989), .I3(n8_adj_3988), .O(n25693));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17747));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [4]), 
            .I2(\FRAME_MATCHER.state [6]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n25503));
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17746));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n91));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17745));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17744));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1002 (.I0(n25503), .I1(n25693), .I2(n25687), 
            .I3(GND_net), .O(n15879));
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17743));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_1003 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(ID1), .I3(ID0), .O(n12_adj_3990));   // verilog/coms.v(230[12:32])
    defparam i4_4_lut_adj_1003.LUT_INIT = 16'h7bde;
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17742));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17741));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17740));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17739));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17738));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17737));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17736));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17735));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17734));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17733));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17732));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1004 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [2]), 
            .I2(ID2), .I3(GND_net), .O(n10_adj_3991));   // verilog/coms.v(230[12:32])
    defparam i2_3_lut_adj_1004.LUT_INIT = 16'hbebe;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17731));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[0] [6]), .I1(n12_adj_3990), .I2(\data_in_frame[0] [4]), 
            .I3(GND_net), .O(n14_adj_3992));   // verilog/coms.v(230[12:32])
    defparam i6_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17730));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_1005 (.I0(\data_in_frame[0] [3]), .I1(n14_adj_3992), 
            .I2(n10_adj_3991), .I3(\data_in_frame[0] [7]), .O(n13455));   // verilog/coms.v(230[12:32])
    defparam i7_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17729));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 data_in_frame_12__7__I_0_3226_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_760));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_12__7__I_0_3226_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17728));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17727));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1006 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16514));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17726));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35645));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17725));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35966));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17724));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17723));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i29_4_lut (.I0(\data_in_frame[12] [5]), .I1(n35892), .I2(n36071), 
            .I3(n35808), .O(n74));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17722));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17721));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17720));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17719));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17718));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17717));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4][2] ), .C(clk32MHz), 
           .D(n17716));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4][1] ), .C(clk32MHz), 
           .D(n17715));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i28_4_lut (.I0(n35814), .I1(n35494), .I2(n35639), .I3(\data_in_frame[8] [1]), 
            .O(n73));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(\data_in_frame[13] [2]), .I1(n16137), .I2(n35574), 
            .I3(n35996), .O(n71));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1009 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n48));
    defparam i3_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_LUT4 i25_4_lut (.I0(Kp_23__N_1406), .I1(n35645), .I2(n35984), .I3(\data_in_frame[13] [3]), 
            .O(n70));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(\data_in_frame[14] [0]), .I1(n70), .I2(n48), 
            .I3(n36059), .O(n80));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n16630), .I1(n35987), .I2(n36098), .I3(n35491), 
            .O(n78));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n16276), .I1(\data_in_frame[12] [1]), .I2(\data_in_frame[9] [5]), 
            .I3(Kp_23__N_760), .O(n76));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(\data_in_frame[6] [4]), .I1(n36062), .I2(n16371), 
            .I3(Kp_23__N_893), .O(n77));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n35737), .I1(n35568), .I2(n35633), .I3(n35836), 
            .O(n75));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i41_4_lut (.I0(n71), .I1(n73), .I2(n72), .I3(n74), .O(n86));
    defparam i41_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i40_4_lut (.I0(n16919), .I1(n80), .I2(n68), .I3(n16802), 
            .O(n85));
    defparam i40_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i42_4_lut (.I0(n75), .I1(n77), .I2(n76), .I3(n78), .O(n87));
    defparam i42_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1010 (.I0(\data_in_frame[15] [1]), .I1(n87), .I2(n85), 
            .I3(n86), .O(n36065));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(n35500), .I1(n36065), .I2(\data_in_frame[15] [0]), 
            .I3(GND_net), .O(n35843));
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1012 (.I0(\data_in_frame[16] [0]), .I1(n35843), 
            .I2(n35820), .I3(\data_in_frame[15] [7]), .O(n31231));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1013 (.I0(\data_in_frame[13] [4]), .I1(n16496), 
            .I2(n32001), .I3(\data_in_frame[11] [3]), .O(n35719));
    defparam i3_4_lut_adj_1013.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1014 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[8] [5]), .I3(GND_net), .O(n36095));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1014.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1015 (.I0(\data_in_frame[8] [6]), .I1(n36095), 
            .I2(n16076), .I3(\data_in_frame[10] [7]), .O(n35494));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(\data_in_frame[13] [3]), .I1(n35719), 
            .I2(GND_net), .I3(GND_net), .O(n35922));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1017 (.I0(n31488), .I1(n31114), .I2(n35923), 
            .I3(n31231), .O(n35963));
    defparam i3_4_lut_adj_1017.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[15] [6]), .I1(n35963), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3993));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1019 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(n35843), .I3(n6_adj_3993), .O(n31202));
    defparam i4_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4][0] ), .C(clk32MHz), 
           .D(n17714));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17713));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17712));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17711));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17710));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17709));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17708));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17707));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17706));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17705));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17704));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17703));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17702));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17701));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17700));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17699));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17698));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17697));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17696));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17695));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17694));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17693));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17692));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17691));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17690));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n17689));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n17688));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n17687));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n17686));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n17685));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17684));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n17683));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17682));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17681));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17680));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17679));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17678));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17677));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17676));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20239_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), .I2(n63_adj_3994), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(138[4] 140[7])
    defparam i20239_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_381_Select_2_i5_4_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2390 ), 
            .I2(n2855), .I3(n63), .O(n5));
    defparam select_381_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i19971_3_lut (.I0(n122), .I1(n3741), .I2(n63), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2586[2] ));   // verilog/coms.v(248[6] 250[9])
    defparam i19971_3_lut.LUT_INIT = 16'hecec;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17675));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17674));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17673));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17672));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17671));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20390_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n41084));
    defparam i20390_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36658_4_lut (.I0(byte_transmit_counter[7]), .I1(n25745), .I2(byte_transmit_counter[6]), 
            .I3(byte_transmit_counter[5]), .O(tx_transmit_N_3220));
    defparam i36658_4_lut.LUT_INIT = 16'h0001;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17670));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17669));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n17668));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n17667));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n17666));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n17665));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n17664));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n17663));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n17662));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n17661));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15862));   // verilog/coms.v(158[5:29])
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'hbbbb;
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n17660));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n17659));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n17658));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n17657));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n17656));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n17655));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n17654));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n17653));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20140_4_lut (.I0(n10_adj_3997), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n15974), .O(n3741));   // verilog/coms.v(248[9:58])
    defparam i20140_4_lut.LUT_INIT = 16'h3332;
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n17652));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n17651));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n17650));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n17649));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n17648));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n17647));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n17646));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17645));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17644));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i29559_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36328));   // verilog/coms.v(110[11:16])
    defparam i29559_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1021 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n15879), .I3(n36328), .O(n38180));
    defparam i3_4_lut_adj_1021.LUT_INIT = 16'h0002;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17643));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17642));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17641));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17640));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17639));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17638));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17637));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17636));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17635));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17634));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1022 (.I0(n2086), .I1(n37242), .I2(\FRAME_MATCHER.i_31__N_2388 ), 
            .I3(n38180), .O(n2778));
    defparam i3_4_lut_adj_1022.LUT_INIT = 16'h0004;
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17633));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17632));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17631));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17630));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17629));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17628));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17627));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17626));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17625));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17624));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n17957));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1023 (.I0(n15729), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3998));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i20135_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3998), .I3(\FRAME_MATCHER.i [1]), .O(n737));   // verilog/coms.v(154[9:60])
    defparam i20135_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i17_4_lut_adj_1024 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i17_4_lut_adj_1024.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(n31202), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35990));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_in_frame[15] [6]), .I1(n16173), 
            .I2(GND_net), .I3(GND_net), .O(n35820));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1027 (.I0(n16592), .I1(n35856), .I2(\data_in_frame[8] [5]), 
            .I3(\data_in_frame[12] [7]), .O(Kp_23__N_1418));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\data_in_frame[17] [1]), .I1(Kp_23__N_1418), 
            .I2(GND_net), .I3(GND_net), .O(n36020));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[16] [4]), .I1(n31987), 
            .I2(GND_net), .I3(GND_net), .O(n35733));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1030 (.I0(\data_in_frame[18] [4]), .I1(n35733), 
            .I2(\data_in_frame[18] [5]), .I3(n35928), .O(n35805));
    defparam i3_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1031 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[17] [2]), .I3(GND_net), .O(n35969));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1031.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[8] [4]), .I1(n16197), 
            .I2(GND_net), .I3(GND_net), .O(n16564));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_1033 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [16]), .O(n40));
    defparam i15_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1034 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n48_adj_3999));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [27]), .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1035 (.I0(\data_in_frame[10] [7]), .I1(n35531), 
            .I2(n35527), .I3(n6_adj_4000), .O(n35856));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(n35497), .I1(n35787), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4001));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1037 (.I0(n35839), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[14] [7]), .I3(n6_adj_4001), .O(n36107));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1038 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n14_adj_4002));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_1038.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1039 (.I0(n36107), .I1(n36053), .I2(n35856), 
            .I3(n31210), .O(n15_adj_4003));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1040 (.I0(n15_adj_4003), .I1(n36092), .I2(n14_adj_4002), 
            .I3(n35969), .O(n35676));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1041 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(n4_adj_3979), .I3(n6_adj_4004), .O(n16306));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(n16306), .I1(n16557), .I2(GND_net), 
            .I3(GND_net), .O(n35836));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n31156), .I1(n35772), .I2(n35775), 
            .I3(\data_in_frame[11] [4]), .O(n31114));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(n31200), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35772));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1045 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n14_adj_4005));
    defparam i5_3_lut_adj_1045.LUT_INIT = 16'h9696;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48_adj_3999), .I2(n37), .I3(n38), 
            .O(n15974));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1046 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4006));
    defparam i5_3_lut_adj_1046.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1047 (.I0(\data_in[0] [6]), .I1(n15971), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4007));
    defparam i6_4_lut_adj_1047.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1048 (.I0(\data_in_frame[12] [0]), .I1(n31114), 
            .I2(n35836), .I3(n35996), .O(n15_adj_4008));
    defparam i6_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1049 (.I0(n15_adj_4008), .I1(n35630), .I2(n14_adj_4005), 
            .I3(\data_in_frame[11] [7]), .O(n35928));
    defparam i8_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(n35928), .I1(n36050), .I2(n35772), 
            .I3(GND_net), .O(n31964));
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1406));   // verilog/coms.v(68[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1051 (.I0(n16496), .I1(n35775), .I2(\data_in_frame[15] [6]), 
            .I3(\data_in_frame[13] [4]), .O(n12_adj_4009));
    defparam i5_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1052 (.I0(\data_in_frame[16] [0]), .I1(n12_adj_4009), 
            .I2(n35956), .I3(\data_in_frame[13] [5]), .O(n32016));
    defparam i6_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35999));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1054 (.I0(n35999), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[12] [2]), .I3(n36074), .O(n10_adj_4010));
    defparam i4_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1055 (.I0(n35839), .I1(n10_adj_4010), .I2(\data_in_frame[12] [0]), 
            .I3(GND_net), .O(n35808));
    defparam i5_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35468));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\data_in_frame[3] [2]), .I1(n35829), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4011));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1058 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(n6_adj_4011), .O(n16557));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16630));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1060 (.I0(n15_adj_4007), .I1(\data_in[2] [2]), 
            .I2(n14_adj_4006), .I3(\data_in[0] [3]), .O(n15769));
    defparam i8_4_lut_adj_1060.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1061 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4012));
    defparam i6_4_lut_adj_1061.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1062 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4013));
    defparam i7_4_lut_adj_1062.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_4_lut_adj_1063 (.I0(\data_in_frame[10] [3]), .I1(\data_in_frame[10] [2]), 
            .I2(\data_in_frame[8] [2]), .I3(\data_in_frame[12] [4]), .O(n36071));
    defparam i3_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1064 (.I0(n16197), .I1(n36071), .I2(n16630), 
            .I3(n16557), .O(n35497));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35984));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1066 (.I0(n16557), .I1(\data_in_frame[9] [4]), 
            .I2(n35808), .I3(n6_adj_4014), .O(n31987));
    defparam i4_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4015));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(n35601), .I1(n35497), .I2(n35688), 
            .I3(n6_adj_4015), .O(n35481));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16192));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1070 (.I0(n16192), .I1(n35481), .I2(\data_in_frame[18] [6]), 
            .I3(n31987), .O(n36967));
    defparam i3_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(n16919), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35901));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35531));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[7] [0]), .I1(n35568), 
            .I2(GND_net), .I3(GND_net), .O(n16808));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16076));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\data_in_frame[6] [4]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n35664));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1076 (.I0(n17_adj_4013), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4012), .I3(\data_in[3] [7]), .O(n15859));
    defparam i9_4_lut_adj_1076.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1077 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4016));
    defparam i4_4_lut_adj_1077.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1078 (.I0(\data_in[2] [7]), .I1(n10_adj_4016), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n15971));
    defparam i5_3_lut_adj_1078.LUT_INIT = 16'hdfdf;
    SB_LUT4 i4_4_lut_adj_1079 (.I0(\data_in_frame[9] [0]), .I1(n35531), 
            .I2(n35901), .I3(n6_adj_4017), .O(n16496));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(\data_in_frame[14] [7]), .I1(n16496), 
            .I2(GND_net), .I3(GND_net), .O(n16748));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1081 (.I0(\data_in_frame[15] [1]), .I1(n16748), 
            .I2(\data_in_frame[15] [3]), .I3(\data_in_frame[19] [5]), .O(n36101));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1082 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n35762), .I3(n16371), .O(n35630));
    defparam i3_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35723));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_0__1__I_0_2_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_847));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_0__1__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(\data_in_frame[5] [1]), .I1(n35475), 
            .I2(n35723), .I3(n31100), .O(n31224));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(n31190), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[4] [6]), .I3(n31224), .O(n35987));
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1086 (.I0(\data_in_frame[4] [4]), .I1(n4_adj_4018), 
            .I2(Kp_23__N_847), .I3(\data_in_frame[2] [2]), .O(n16974));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_in_frame[7] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35814));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1088 (.I0(n31979), .I1(\data_in_frame[9] [2]), 
            .I2(n35814), .I3(\data_in_frame[6] [7]), .O(n16_adj_4019));
    defparam i6_4_lut_adj_1088.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1089 (.I0(\data_in_frame[6] [6]), .I1(n16974), 
            .I2(n35987), .I3(\data_in_frame[4] [6]), .O(n17_adj_4020));
    defparam i7_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1090 (.I0(n17_adj_4020), .I1(\data_in_frame[7] [0]), 
            .I2(n16_adj_4019), .I3(n31222), .O(n31156));
    defparam i9_4_lut_adj_1090.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35589));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1092 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4021));
    defparam i2_2_lut_adj_1092.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1093 (.I0(n35667), .I1(\data_in_frame[5] [0]), 
            .I2(n4_adj_3979), .I3(GND_net), .O(n31222));
    defparam i2_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(\data_in_frame[6] [6]), .I1(n31222), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n36098));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35625));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1096 (.I0(\data_in_frame[4] [3]), .I1(n35625), 
            .I2(\data_in_frame[0] [1]), .I3(\data_in_frame[1] [7]), .O(n16218));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1097 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[6] [5]), .O(n12_adj_4022));
    defparam i5_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1098 (.I0(n16218), .I1(n12_adj_4022), .I2(n35798), 
            .I3(\data_in_frame[7] [1]), .O(n32001));
    defparam i6_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1099 (.I0(\data_in_frame[11] [4]), .I1(n31156), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n35737));
    defparam i2_3_lut_adj_1099.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1100 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35956));
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(n31488), .I1(n35956), .I2(n16173), 
            .I3(\data_in_frame[15] [7]), .O(n36050));
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35519));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1103 (.I0(n4_adj_4018), .I1(n5_c), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n16919));
    defparam i2_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_in_frame[6] [7]), .I1(n16919), 
            .I2(GND_net), .I3(GND_net), .O(n16971));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1105 (.I0(n31959), .I1(n35741), .I2(n16971), 
            .I3(\data_in_frame[9] [3]), .O(n12_adj_4023));
    defparam i5_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1106 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4024));
    defparam i6_4_lut_adj_1106.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1107 (.I0(\data_in[3] [6]), .I1(n14_adj_4024), 
            .I2(n10_adj_4021), .I3(\data_in[2] [1]), .O(n15856));
    defparam i7_4_lut_adj_1107.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1108 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n15856), .I3(\data_in[1] [0]), .O(n18_adj_4025));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1109 (.I0(\data_in[1] [4]), .I1(n18_adj_4025), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n20_adj_4026));
    defparam i9_4_lut_adj_1109.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_1110 (.I0(n15_adj_4027), .I1(n20_adj_4026), .I2(n15859), 
            .I3(\data_in[0] [6]), .O(n63_c));
    defparam i10_4_lut_adj_1110.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1111 (.I0(\data_in_frame[9] [4]), .I1(n12_adj_4023), 
            .I2(\data_in_frame[11] [5]), .I3(\data_in_frame[7] [1]), .O(n31200));
    defparam i6_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16142));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_in_frame[5] [7]), .I1(n16624), 
            .I2(GND_net), .I3(GND_net), .O(n16802));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35633));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(Kp_23__N_946), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16532));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1116 (.I0(n16532), .I1(n35633), .I2(n16802), 
            .I3(GND_net), .O(n35972));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1116.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[6] [2]), .I1(n10_adj_4028), 
            .I2(GND_net), .I3(GND_net), .O(n16567));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(n16197), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16916));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1119 (.I0(\data_in_frame[1] [5]), .I1(n35595), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[4] [1]), .O(n10_adj_4028));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4029));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1121 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[1] [6]), .I3(n6_adj_4029), .O(n11));   // verilog/coms.v(228[9:81])
    defparam i4_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1122 (.I0(\data_in_frame[4] [0]), .I1(n35713), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[1] [4]), .O(n16197));   // verilog/coms.v(228[9:81])
    defparam i3_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1123 (.I0(n11), .I1(\data_in_frame[6] [3]), .I2(n10_adj_4028), 
            .I3(GND_net), .O(n35527));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(Kp_23__N_946), .I1(n35527), .I2(n16197), 
            .I3(GND_net), .O(n35491));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35892));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1126 (.I0(\data_in_frame[8] [3]), .I1(n35892), 
            .I2(n35642), .I3(n35491), .O(n16592));   // verilog/coms.v(70[16:41])
    defparam i3_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n35839));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1128 (.I0(n15769), .I1(\data_in[0] [7]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_4030));
    defparam i6_4_lut_adj_1128.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1129 (.I0(n15859), .I1(\data_in[3] [1]), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n17_adj_4031));
    defparam i7_4_lut_adj_1129.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1130 (.I0(n17_adj_4031), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4030), .I3(\data_in[0] [2]), .O(n63_adj_3994));
    defparam i9_4_lut_adj_1130.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(\data_in_frame[7] [4]), .I1(n16306), 
            .I2(\data_in_frame[10] [0]), .I3(n16624), .O(n10_adj_4032));
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1132 (.I0(n36020), .I1(\data_in_frame[14] [5]), 
            .I2(n31170), .I3(n35895), .O(n15_adj_4033));
    defparam i6_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1133 (.I0(n15_adj_4033), .I1(n16748), .I2(n14_adj_4034), 
            .I3(\data_in_frame[15] [1]), .O(n31210));
    defparam i8_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4035));   // verilog/coms.v(74[16:43])
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1134 (.I0(\data_in_frame[14] [7]), .I1(n35601), 
            .I2(\data_in_frame[16] [6]), .I3(n35839), .O(n24_adj_4036));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1135 (.I0(\data_in_frame[19] [2]), .I1(n35688), 
            .I2(\data_in_frame[12] [6]), .I3(\data_in_frame[15] [0]), .O(n22_adj_4037));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1136 (.I0(n16592), .I1(n24_adj_4036), .I2(n18_adj_4035), 
            .I3(\data_in_frame[14] [6]), .O(n26));   // verilog/coms.v(74[16:43])
    defparam i12_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1137 (.I0(n16916), .I1(n26), .I2(n22_adj_4037), 
            .I3(n35888), .O(n35801));   // verilog/coms.v(74[16:43])
    defparam i13_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16784));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1139 (.I0(\data_in_frame[3] [4]), .I1(n35583), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[5] [6]), .O(n16624));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35642));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1141 (.I0(\data_in_frame[10] [3]), .I1(n16624), 
            .I2(n16784), .I3(Kp_23__N_946), .O(n10_adj_4038));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_in_frame[7] [3]), .I1(n31224), 
            .I2(GND_net), .I3(GND_net), .O(n31959));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16137));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[16] [5]), .I3(GND_net), .O(n35784));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1145 (.I0(n15856), .I1(\data_in[3] [7]), .I2(n15769), 
            .I3(\data_in[1] [6]), .O(n20_adj_4039));
    defparam i8_4_lut_adj_1145.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1146 (.I0(\data_in[1] [3]), .I1(\data_in[2] [6]), 
            .I2(\data_in[0] [5]), .I3(\data_in[1] [2]), .O(n19_adj_4040));
    defparam i7_4_lut_adj_1146.LUT_INIT = 16'hdfff;
    SB_LUT4 i32316_4_lut (.I0(\data_in[3] [2]), .I1(\data_in[2] [5]), .I2(\data_in[0] [1]), 
            .I3(\data_in[2] [0]), .O(n39097));
    defparam i32316_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n39097), .I1(n19_adj_4040), .I2(n20_adj_4039), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1147 (.I0(n35888), .I1(n35744), .I2(\data_in_frame[18] [7]), 
            .I3(\data_in_frame[14] [6]), .O(n18_adj_4041));
    defparam i7_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1148 (.I0(n16137), .I1(n18_adj_4041), .I2(\data_in_frame[19] [1]), 
            .I3(n31959), .O(n20_adj_4042));
    defparam i9_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1149 (.I0(n36017), .I1(n35784), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4043));
    defparam i4_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1150 (.I0(n15_adj_4043), .I1(n20_adj_4042), .I2(n35535), 
            .I3(n31979), .O(n35564));
    defparam i10_4_lut_adj_1150.LUT_INIT = 16'h9669;
    SB_LUT4 i3_2_lut_3_lut (.I0(n24660), .I1(n25346), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n8_adj_3964));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35622));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35583));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35713));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1154 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[1] [5]), 
            .I2(n35875), .I3(\data_in_frame[1] [7]), .O(n35475));   // verilog/coms.v(71[16:34])
    defparam i3_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1155 (.I0(\data_in_frame[2] [7]), .I1(Kp_23__N_893), 
            .I2(n35595), .I3(n35875), .O(n20_adj_4044));   // verilog/coms.v(163[9:87])
    defparam i8_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(n35925), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [6]), .I3(n35829), .O(n19_adj_4045));   // verilog/coms.v(163[9:87])
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1157 (.I0(n35625), .I1(\data_in_frame[2] [3]), 
            .I2(n35589), .I3(Kp_23__N_847), .O(n21_adj_4046));   // verilog/coms.v(163[9:87])
    defparam i9_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1158 (.I0(n21_adj_4046), .I1(n19_adj_4045), .I2(n20_adj_4044), 
            .I3(GND_net), .O(n37788));   // verilog/coms.v(163[9:87])
    defparam i11_3_lut_adj_1158.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1159 (.I0(n37788), .I1(n35853), .I2(n35583), 
            .I3(n35622), .O(n12_adj_4047));   // verilog/coms.v(71[16:34])
    defparam i5_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1160 (.I0(\data_in_frame[1] [7]), .I1(n12_adj_4047), 
            .I2(\data_in_frame[1] [0]), .I3(n35713), .O(n31100));   // verilog/coms.v(71[16:34])
    defparam i6_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1161 (.I0(n31100), .I1(\data_in_frame[3] [0]), 
            .I2(n35475), .I3(\data_in_frame[0] [6]), .O(n35667));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1162 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_c));   // verilog/coms.v(163[9:87])
    defparam i2_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(n24660), .I1(n25346), .I2(n13_adj_3984), 
            .I3(\FRAME_MATCHER.i_31__N_2388 ), .O(n17100));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff02;
    SB_LUT4 equal_1197_i15_2_lut (.I0(Kp_23__N_893), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4048));   // verilog/coms.v(228[9:81])
    defparam equal_1197_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(n16306), .I1(n31222), .I2(GND_net), 
            .I3(GND_net), .O(n35741));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(n31190), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n31979));
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1165 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[7] [3]), 
            .I2(n8_adj_4049), .I3(n15_adj_4048), .O(n36074));
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1166 (.I0(n35999), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[12] [1]), .I3(\data_in_frame[7] [6]), .O(n35744));
    defparam i3_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1167 (.I0(\data_in_frame[0] [7]), .I1(n35853), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n16276));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(n31200), .I1(\data_in_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36059));
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(n16276), .I1(n35744), .I2(GND_net), 
            .I3(GND_net), .O(n35943));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1170 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(n6_adj_4050), .I3(n35723), .O(n16371));
    defparam i1_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[9] [4]), .I1(n36074), 
            .I2(GND_net), .I3(GND_net), .O(n35884));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1172 (.I0(n35943), .I1(\data_in_frame[7] [5]), 
            .I2(\data_in_frame[14] [2]), .I3(n36059), .O(n10_adj_4051));
    defparam i4_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1173 (.I0(n35884), .I1(\data_in_frame[16] [3]), 
            .I2(n10_adj_4051), .I3(n16371), .O(n10_adj_4052));
    defparam i3_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(Kp_23__N_1418), .I1(\data_in_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16824));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35787));
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i4_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n24_adj_4053));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35730));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1177 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[16] [2]), 
            .I2(n35784), .I3(n16192), .O(n10_adj_4054));
    defparam i4_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1178 (.I0(n32016), .I1(\data_in_frame[18] [3]), 
            .I2(n16514), .I3(n35969), .O(n34));
    defparam i14_4_lut_adj_1178.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1179 (.I0(n31231), .I1(n35805), .I2(n10_adj_4054), 
            .I3(\data_in_frame[16] [3]), .O(n25));
    defparam i5_4_lut_adj_1179.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1180 (.I0(n35564), .I1(n24_adj_4053), .I2(n16916), 
            .I3(n35801), .O(n32_adj_4055));
    defparam i12_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1181 (.I0(n36005), .I1(n35676), .I2(n35859), 
            .I3(n31964), .O(n31_adj_4056));
    defparam i11_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1182 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[18] [7]), 
            .I2(n35730), .I3(n35733), .O(n35));
    defparam i15_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1183 (.I0(n25), .I1(n34), .I2(n31962), .I3(n36020), 
            .O(n37_adj_4057));
    defparam i17_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n37_adj_4057), .I1(n35), .I2(n31_adj_4056), 
            .I3(n32_adj_4055), .O(n37969));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1184 (.I0(n35943), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[16] [5]), .I3(n36017), .O(n10_adj_4058));
    defparam i4_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1185 (.I0(n35762), .I1(n10_adj_4058), .I2(n31170), 
            .I3(GND_net), .O(n31794));
    defparam i5_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1186 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n14_adj_4059));
    defparam i5_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1187 (.I0(n35922), .I1(n31962), .I2(n35895), 
            .I3(\data_in_frame[20] [2]), .O(n15_adj_4060));
    defparam i6_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1188 (.I0(\data_in_frame[17] [2]), .I1(n35888), 
            .I2(n35859), .I3(n35966), .O(n15_adj_4061));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1189 (.I0(n15_adj_4061), .I1(n36026), .I2(n14_adj_4062), 
            .I3(n35694), .O(n37640));   // verilog/coms.v(73[16:43])
    defparam i8_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1190 (.I0(n36062), .I1(n36107), .I2(n37640), 
            .I3(\data_in_frame[21] [6]), .O(n10_adj_4063));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_in_frame[20] [3]), .I1(n35730), 
            .I2(n32016), .I3(n31202), .O(n37446));
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1192 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(n35719), .I3(n16916), .O(n18_adj_4064));   // verilog/coms.v(71[16:42])
    defparam i7_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1193 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4065));   // verilog/coms.v(71[16:42])
    defparam i5_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1194 (.I0(\data_in_frame[13] [0]), .I1(n18_adj_4064), 
            .I2(n35500), .I3(n35972), .O(n20_adj_4066));   // verilog/coms.v(71[16:42])
    defparam i9_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1195 (.I0(\data_in_frame[17] [4]), .I1(n16_adj_4065), 
            .I2(n35661), .I3(\data_in_frame[17] [6]), .O(n19_adj_4067));   // verilog/coms.v(71[16:42])
    defparam i8_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_86_2_lut (.I0(n35564), .I1(n35801), .I2(GND_net), .I3(GND_net), 
            .O(n44816));
    defparam i1_rep_86_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1196 (.I0(\data_in_frame[21] [7]), .I1(n36005), 
            .I2(n35859), .I3(n16916), .O(n36896));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1197 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[21] [1]), 
            .I2(n44816), .I3(n37969), .O(n20_adj_4068));
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'hde7b;
    SB_LUT4 i5_3_lut_adj_1198 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[20] [1]), 
            .I2(n35963), .I3(GND_net), .O(n14_adj_4069));
    defparam i5_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1199 (.I0(n36065), .I1(\data_in_frame[13] [1]), 
            .I2(n16173), .I3(n35990), .O(n15_adj_4070));
    defparam i6_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1200 (.I0(n35481), .I1(\data_in_frame[20] [7]), 
            .I2(n35733), .I3(\data_in_frame[16] [6]), .O(n16_adj_4071));
    defparam i6_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1201 (.I0(n31794), .I1(\data_in_frame[13] [7]), 
            .I2(n37969), .I3(\data_in_frame[18] [5]), .O(n17_adj_4072));
    defparam i7_4_lut_adj_1201.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1202 (.I0(n15_adj_4070), .I1(n35787), .I2(n14_adj_4069), 
            .I3(n16824), .O(n37311));
    defparam i8_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(n35564), .I1(\data_in_frame[21] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4073));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1204 (.I0(n15_adj_4060), .I1(\data_in_frame[13] [2]), 
            .I2(n14_adj_4059), .I3(\data_in_frame[17] [7]), .O(n37705));
    defparam i8_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1205 (.I0(n37311), .I1(n17_adj_4072), .I2(n10_adj_4052), 
            .I3(n16_adj_4071), .O(n21_adj_4074));
    defparam i5_4_lut_adj_1205.LUT_INIT = 16'hebbe;
    SB_LUT4 i5_3_lut_adj_1206 (.I0(n31200), .I1(n10_adj_4052), .I2(\data_in_frame[18] [4]), 
            .I3(GND_net), .O(n12_adj_4075));
    defparam i5_3_lut_adj_1206.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1207 (.I0(\data_in_frame[21] [4]), .I1(n35801), 
            .I2(\data_in_frame[19] [3]), .I3(n31210), .O(n37238));
    defparam i3_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i32285_4_lut (.I0(n36101), .I1(n37446), .I2(n10_adj_4063), 
            .I3(\data_in_frame[19] [4]), .O(n39065));
    defparam i32285_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i6_4_lut_adj_1208 (.I0(\data_in_frame[20] [5]), .I1(n12_adj_4075), 
            .I2(n36050), .I3(\data_in_frame[18] [3]), .O(n37275));
    defparam i6_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1209 (.I0(n21_adj_4074), .I1(n36967), .I2(n37705), 
            .I3(n4_adj_4073), .O(n27_adj_4076));
    defparam i11_4_lut_adj_1209.LUT_INIT = 16'hfbfe;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(n32016), .I1(\data_in_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4077));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1211 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[20] [4]), 
            .I2(n31964), .I3(n6_adj_4077), .O(n36860));
    defparam i4_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1212 (.I0(\data_in_frame[20] [6]), .I1(n19_adj_4067), 
            .I2(n35805), .I3(n20_adj_4066), .O(n18_adj_4078));
    defparam i2_4_lut_adj_1212.LUT_INIT = 16'hde7b;
    SB_LUT4 i10_4_lut_adj_1213 (.I0(\data_in_frame[21] [5]), .I1(n20_adj_4068), 
            .I2(n36896), .I3(n35676), .O(n26_adj_4079));
    defparam i10_4_lut_adj_1213.LUT_INIT = 16'hdfef;
    SB_LUT4 i14_4_lut_adj_1214 (.I0(n27_adj_4076), .I1(n37275), .I2(n39065), 
            .I3(n37238), .O(n30_adj_4080));
    defparam i14_4_lut_adj_1214.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(\data_in_frame[21] [0]), .I1(n36860), 
            .I2(n36967), .I3(n37969), .O(n17_adj_4081));
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'hedde;
    SB_LUT4 i15_4_lut_adj_1216 (.I0(n17_adj_4081), .I1(n30_adj_4080), .I2(n26_adj_4079), 
            .I3(n18_adj_4078), .O(n31_adj_4082));
    defparam i15_4_lut_adj_1216.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[16][5] ), .I1(n31164), .I2(\data_out_frame[17] [0]), 
            .I3(GND_net), .O(n32004));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i120_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));
    defparam i120_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1217 (.I0(n13455), .I1(n15879), .I2(n91), .I3(n39023), 
            .O(n17068));
    defparam i4_4_lut_adj_1217.LUT_INIT = 16'h0010;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3975), .S(n3_adj_3968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n17935));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n17956));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3974), .S(n3_adj_3960));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3973), .S(n3_adj_3959));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3972), .S(n3_adj_3958));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3971), .S(n3_adj_3957));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3970), .S(n3_adj_3956));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3969), .S(n3_adj_3955));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3967), .S(n3_adj_3954));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3966), .S(n3_adj_3953));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3965), .S(n3_adj_3952));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3963), .S(n3_adj_3951));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3962), .S(n3_adj_3950));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3961), .S(n3_adj_3949));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3922), .S(n3_adj_3948));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3912), .S(n3_adj_3947));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3911), .S(n3_adj_3946));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3898), .S(n3_adj_3945));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3895), .S(n3_adj_3944));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3921), .S(n3_adj_3943));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3942));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4083), .S(n3_adj_3941));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4084), .S(n3_adj_3940));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4085), .S(n3_adj_3939));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4086), .S(n3_adj_3938));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4087), .S(n3_adj_3937));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4088), .S(n3_adj_3936));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4089), .S(n3_adj_3935));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4090), .S(n3_adj_3934));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4091), .S(n3_adj_3933));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4092), .S(n3_adj_3932));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4093), .S(n3_adj_3931));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n17955));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n17124), .D(n36731));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n17124), .D(n37263));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n17124), .D(n36725));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n17124), .D(n37260));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n17124), .D(n37444));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n17124), .D(n37402));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n17124), .D(n37040));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n17124), .D(n37659));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n17124), .D(n37704));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n17124), .D(n37148));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n17124), .D(n35540));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n17124), .D(n37006));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n17124), .D(n37420));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n17124), .D(n35698));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n17124), .D(n37234));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n17124), .D(n35652));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n34722), .S(n34894));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[3] [3]), .O(n35853));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n35400), .S(n34724));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n7_adj_4094), .S(n8_adj_4095));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n35403), .S(n34798));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n35397), .S(n34796));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n35406), .S(n34794));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n35391), .S(n34792));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n35390), .S(n34720));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n35392), .S(n34790));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n35407), .S(n34788));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n35398), .S(n34786));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n35404), .S(n34784));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n35401), .S(n34782));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n35409), .S(n34780));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n35394), .S(n34778));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_4096), .S(n8_adj_4097));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n35395), .S(n34776));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n7_adj_4098), .S(n8_adj_4099));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n35393), .S(n34774));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n24653), .S(n25478));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n35408), .S(n34772));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n7_adj_4100), .S(n8_adj_4101));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n37102), .S(n34680));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n7_adj_4102), .S(n8_adj_4103));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n35399), .S(n34732));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n35402), .S(n34770));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n35396), .S(n34768));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n35405), .S(n34766));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n35389), .S(n25470));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17623));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n17954));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1218 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [6]), .I3(n35583), .O(n35875));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i19939_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n24660));
    defparam i19939_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(n35607), .I2(n35610), 
            .I3(\data_in_frame[1] [7]), .O(n24_adj_3980));   // verilog/coms.v(163[9:87])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0990;
    SB_LUT4 i1_2_lut_3_lut_adj_1219 (.I0(\data_out_frame[16][5] ), .I1(n31164), 
            .I2(\data_out_frame[18] [7]), .I3(GND_net), .O(n36047));
    defparam i1_2_lut_3_lut_adj_1219.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1220 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n35996));
    defparam i1_2_lut_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1221 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[14] [3]), .O(n36017));
    defparam i2_3_lut_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i20086_2_lut_3_lut (.I0(n63_adj_3994), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));
    defparam i20086_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1222 (.I0(n63_adj_3994), .I1(n63_c), .I2(n63), 
            .I3(GND_net), .O(n10454));
    defparam i1_2_lut_3_lut_adj_1222.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1223 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n14_adj_4104));
    defparam i1_2_lut_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i23_3_lut_4_lut (.I0(n35737), .I1(n32001), .I2(\data_in_frame[13] [1]), 
            .I3(\data_in_frame[6] [2]), .O(n68));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_41_24 (.CI(n28491), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n28492));
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n17953));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n17952));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n17951));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n17950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n17949));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n17948));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n17947));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n17946));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(n35737), .I1(n32001), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n16173));
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n17945));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18012));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(n16218), .I1(n16974), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(n36062));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_33_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n28500), .O(n2_adj_4093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_32_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n28499), .O(n2_adj_4092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_32 (.CI(n28499), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n28500));
    SB_LUT4 add_41_31_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n28498), .O(n2_adj_4091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n44382));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n44382_bdd_4_lut (.I0(n44382), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n44385));
    defparam n44382_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37507 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n44376));
    defparam byte_transmit_counter_0__bdd_4_lut_37507.LUT_INIT = 16'he4aa;
    SB_LUT4 n44376_bdd_4_lut (.I0(n44376), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n44379));
    defparam n44376_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37502 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n44370));
    defparam byte_transmit_counter_0__bdd_4_lut_37502.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(n16218), .I1(n16974), .I2(\data_in_frame[11] [0]), 
            .I3(GND_net), .O(n6_adj_4000));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'h9696;
    SB_LUT4 n44370_bdd_4_lut (.I0(n44370), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n44373));
    defparam n44370_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18011));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(n16218), .I1(n35664), .I2(\data_in_frame[17] [4]), 
            .I3(\data_in_frame[13] [2]), .O(n14_adj_4062));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18010));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18009));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18008));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18007));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18006));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18005));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18004));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18003));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18002));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18001));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18000));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n17944));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n17943));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n17942));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n17941));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n17975));   // verilog/coms.v(126[12] 289[6])
    SB_DFFESR LED_3208 (.Q(LED_c), .C(clk32MHz), .E(n36732), .D(n17291), 
            .R(n38154));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37497 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n44364));
    defparam byte_transmit_counter_0__bdd_4_lut_37497.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut_4_lut (.I0(n63), .I1(n737), .I2(n97), .I3(n16), 
            .O(n7));   // verilog/coms.v(154[6] 156[9])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'haa02;
    SB_CARRY add_41_31 (.CI(n28498), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n28499));
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n17934));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20228_2_lut_3_lut (.I0(n63), .I1(n737), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2458[1] ));   // verilog/coms.v(154[6] 156[9])
    defparam i20228_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n24660), .I1(n13_adj_3984), .I2(tx_transmit_N_3220), 
            .I3(n25346), .O(n16));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h2220;
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n17940));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_30_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n28497), .O(n2_adj_4090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_30_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n17939));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n17938));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n17937));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n17936));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_30 (.CI(n28497), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n28498));
    SB_LUT4 i1_2_lut_4_lut (.I0(n35494), .I1(n35527), .I2(n16808), .I3(n35922), 
            .O(n35923));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_29_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n28496), .O(n2_adj_4089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n44364_bdd_4_lut (.I0(n44364), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16][5] ), .I3(byte_transmit_counter[1]), 
            .O(n44367));
    defparam n44364_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37492 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n44358));
    defparam byte_transmit_counter_0__bdd_4_lut_37492.LUT_INIT = 16'he4aa;
    SB_CARRY add_41_29 (.CI(n28496), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n28497));
    SB_LUT4 n44358_bdd_4_lut (.I0(n44358), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n44361));
    defparam n44358_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_41_28_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n28495), .O(n2_adj_4088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_28_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n17390));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[15] [2]), .I3(\data_out_frame[15] [5]), 
            .O(n8_adj_3906));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17903));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n17999));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_28 (.CI(n28495), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n28496));
    SB_LUT4 i1_2_lut_4_lut_adj_1227 (.I0(n35494), .I1(n35527), .I2(n16808), 
            .I3(Kp_23__N_1427), .O(n35895));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1068_i3_3_lut (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4377), .I3(GND_net), .O(n4380));
    defparam mux_1068_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_27_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n28494), .O(n2_adj_4087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13247_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n17992));
    defparam i13247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_27 (.CI(n28494), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n28495));
    SB_LUT4 mux_1068_i2_3_lut (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4377), .I3(GND_net), .O(n4379));
    defparam mux_1068_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i5_3_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4377), .I3(GND_net), .O(n4382));
    defparam mux_1068_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_26_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n28493), .O(n2_adj_4086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13248_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n17993));
    defparam i13248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n17998));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n17997));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n17996));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1068_i4_3_lut (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4377), .I3(GND_net), .O(n4381));
    defparam mux_1068_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13249_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n17994));
    defparam i13249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17538));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n34728));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17522));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17521));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17520));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n17519));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n17518));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17517));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n17516));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_26 (.CI(n28493), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n28494));
    SB_LUT4 add_41_25_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n28492), .O(n2_adj_4085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_25 (.CI(n28492), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n28493));
    SB_LUT4 add_41_24_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n28491), .O(n2_adj_4084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13242_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n17987));
    defparam i13242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_22 (.CI(n28489), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n28490));
    SB_LUT4 i13243_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n17988));
    defparam i13243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13244_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n17989));
    defparam i13244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13245_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n17990));
    defparam i13245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_23_lut (.I0(n2086), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n28490), .O(n2_adj_4083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_23 (.CI(n28490), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n28491));
    SB_LUT4 i1_2_lut_3_lut_adj_1228 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(n16348), .I3(GND_net), .O(n35652));
    defparam i1_2_lut_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n17995));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [4]), .I3(GND_net), .O(n6_adj_4108));
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n17994));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1230 (.I0(\data_out_frame[20] [3]), .I1(n31967), 
            .I2(n37462), .I3(\data_out_frame[20] [2]), .O(n37420));
    defparam i2_3_lut_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n17993));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(n737), .I1(n10454), .I2(n13_adj_3984), 
            .I3(GND_net), .O(n35383));   // verilog/coms.v(154[6] 156[9])
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'h0404;
    SB_LUT4 i13246_3_lut_4_lut (.I0(n8_adj_4107), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n17991));
    defparam i13246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(n737), .I1(n10454), .I2(n97), 
            .I3(GND_net), .O(n4_adj_4109));   // verilog/coms.v(154[6] 156[9])
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h0404;
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n17992));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1233 (.I0(n96), .I1(n35448), .I2(n35383), 
            .I3(\FRAME_MATCHER.state [30]), .O(n34766));
    defparam i1_2_lut_4_lut_adj_1233.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1234 (.I0(n96), .I1(n35448), .I2(n35383), 
            .I3(\FRAME_MATCHER.state [27]), .O(n34732));
    defparam i1_2_lut_4_lut_adj_1234.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1235 (.I0(n96), .I1(n35448), .I2(n35383), 
            .I3(\FRAME_MATCHER.state [23]), .O(n34772));
    defparam i1_2_lut_4_lut_adj_1235.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1236 (.I0(n96), .I1(n35448), .I2(n35383), 
            .I3(\FRAME_MATCHER.state [4]), .O(n34724));
    defparam i1_2_lut_4_lut_adj_1236.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1237 (.I0(n131), .I1(n61), .I2(n13197), 
            .I3(\FRAME_MATCHER.state [26]), .O(n7_adj_4102));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_4_lut_adj_1237.LUT_INIT = 16'hba00;
    SB_LUT4 equal_113_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4110));   // verilog/coms.v(151[7:23])
    defparam equal_113_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1238 (.I0(n131), .I1(n61), .I2(n13197), 
            .I3(\FRAME_MATCHER.state [24]), .O(n7_adj_4100));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_4_lut_adj_1238.LUT_INIT = 16'hba00;
    SB_LUT4 i19932_2_lut_4_lut (.I0(n131), .I1(n61), .I2(n13197), .I3(\FRAME_MATCHER.state [22]), 
            .O(n24653));   // verilog/coms.v(113[11:12])
    defparam i19932_2_lut_4_lut.LUT_INIT = 16'hba00;
    SB_LUT4 mux_1068_i16_3_lut (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4377), .I3(GND_net), .O(n4393));
    defparam mux_1068_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1239 (.I0(n131), .I1(n61), .I2(n13197), 
            .I3(\FRAME_MATCHER.state [20]), .O(n7_adj_4098));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_4_lut_adj_1239.LUT_INIT = 16'hba00;
    SB_LUT4 mux_1068_i15_3_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4377), .I3(GND_net), .O(n4392));
    defparam mux_1068_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1240 (.I0(n131), .I1(n61), .I2(n13197), 
            .I3(\FRAME_MATCHER.state [18]), .O(n7_adj_4096));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_4_lut_adj_1240.LUT_INIT = 16'hba00;
    SB_LUT4 equal_112_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4107));   // verilog/coms.v(151[7:23])
    defparam equal_112_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1241 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n15974), .I3(\FRAME_MATCHER.i [4]), .O(n15729));   // verilog/coms.v(151[7:23])
    defparam i2_3_lut_4_lut_adj_1241.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1242 (.I0(n131), .I1(n61), .I2(n13197), 
            .I3(\FRAME_MATCHER.state [5]), .O(n7_adj_4094));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_4_lut_adj_1242.LUT_INIT = 16'hba00;
    SB_LUT4 mux_1068_i14_3_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4377), .I3(GND_net), .O(n4391));
    defparam mux_1068_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i13_3_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4377), .I3(GND_net), .O(n4390));
    defparam mux_1068_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1243 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n24972), .O(n35439));   // verilog/coms.v(151[7:23])
    defparam i2_3_lut_4_lut_adj_1243.LUT_INIT = 16'hefff;
    SB_LUT4 mux_1068_i12_3_lut (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4377), .I3(GND_net), .O(n4389));
    defparam mux_1068_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i11_3_lut (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4377), .I3(GND_net), .O(n4388));
    defparam mux_1068_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i10_3_lut (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4377), .I3(GND_net), .O(n4387));
    defparam mux_1068_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i9_3_lut (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4377), .I3(GND_net), .O(n4386));
    defparam mux_1068_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i8_3_lut (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4377), .I3(GND_net), .O(n4385));
    defparam mux_1068_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i24_3_lut (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4377), .I3(GND_net), .O(n4401));
    defparam mux_1068_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i23_3_lut (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4377), .I3(GND_net), .O(n4400));
    defparam mux_1068_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35595));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35925));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1246 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4111), .O(n35431));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1246.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35639));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_LUT4 i3_2_lut_adj_1248 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4112));
    defparam i3_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1249 (.I0(n16532), .I1(n16142), .I2(\data_in_frame[5] [7]), 
            .I3(n16371), .O(n16_adj_4113));
    defparam i7_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1250 (.I0(n35639), .I1(n16_adj_4113), .I2(n12_adj_4112), 
            .I3(n16784), .O(n31170));
    defparam i8_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(n36053), .I1(n36095), .I2(GND_net), 
            .I3(GND_net), .O(n35694));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1252 (.I0(n16564), .I1(n36092), .I2(\data_in_frame[8] [5]), 
            .I3(Kp_23__N_760), .O(n35661));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1253 (.I0(\data_in_frame[8] [6]), .I1(n35901), 
            .I2(n35694), .I3(n35574), .O(Kp_23__N_1427));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(n16276), .I1(n35535), .I2(GND_net), 
            .I3(GND_net), .O(n35859));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1255 (.I0(\data_out_frame[20] [0]), .I1(n2106), 
            .I2(\data_out_frame[19] [4]), .I3(n32044), .O(n14_adj_4114));
    defparam i5_3_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1256 (.I0(n35703), .I1(n16477), .I2(\data_out_frame[17] [6]), 
            .I3(n32012), .O(n30900));
    defparam i2_3_lut_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1257 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[15] [4]), .I3(\data_in_frame[17] [3]), .O(n16_adj_4115));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1258 (.I0(n36101), .I1(Kp_23__N_1427), .I2(n16824), 
            .I3(n35661), .O(n17_adj_4116));   // verilog/coms.v(71[16:42])
    defparam i7_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1259 (.I0(n17_adj_4116), .I1(\data_in_frame[15] [2]), 
            .I2(n16_adj_4115), .I3(n16567), .O(n36005));   // verilog/coms.v(71[16:42])
    defparam i9_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i32417_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39270));
    defparam i32417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32418_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39271));
    defparam i32418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1260 (.I0(\data_out_frame[13] [3]), .I1(n15502), 
            .I2(n35826), .I3(\data_out_frame[15] [4]), .O(n16477));
    defparam i2_3_lut_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i32421_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39274));
    defparam i32421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32420_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39273));
    defparam i32420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1261 (.I0(\data_out_frame[15] [6]), .I1(n36742), 
            .I2(n35703), .I3(GND_net), .O(n6_adj_4117));
    defparam i1_2_lut_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1262 (.I0(\data_out_frame[15] [5]), .I1(n35670), 
            .I2(n10_adj_3900), .I3(\data_out_frame[7] [0]), .O(n35552));
    defparam i1_2_lut_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1263 (.I0(n35703), .I1(n35759), .I2(n32012), 
            .I3(n35867), .O(n6_adj_4118));
    defparam i1_2_lut_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1264 (.I0(n3741), .I1(n10454), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state [1]), .O(n35386));
    defparam i1_2_lut_4_lut_adj_1264.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_adj_1265 (.I0(n10454), .I1(n2778), .I2(n38_adj_4119), 
            .I3(GND_net), .O(n35448));
    defparam i1_2_lut_3_lut_adj_1265.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_3_lut_adj_1266 (.I0(n13142), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n7_adj_4120));
    defparam i1_2_lut_3_lut_adj_1266.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1267 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[8] [1]), .O(n35913));   // verilog/coms.v(95[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1268 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4121), .O(n35432));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1268.LUT_INIT = 16'hffbf;
    SB_LUT4 i27_3_lut_3_lut_4_lut (.I0(\data_in_frame[7] [3]), .I1(n31190), 
            .I2(\data_in_frame[4] [7]), .I3(n36098), .O(n72));
    defparam i27_3_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [7]), .O(n6_adj_4004));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1270 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[9] [5]), .I3(n16052), .O(n35975));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1271 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(n35577), .I3(n35478), .O(n31124));
    defparam i1_2_lut_3_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1272 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4122), .O(n35433));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1272.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_1273 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4110), .O(n35430));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1273.LUT_INIT = 16'hffbf;
    SB_LUT4 i37349_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n17291));
    defparam i37349_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37487 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n44352));
    defparam byte_transmit_counter_0__bdd_4_lut_37487.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1274 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4123), .O(n35434));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1274.LUT_INIT = 16'hffbf;
    SB_LUT4 n44352_bdd_4_lut (.I0(n44352), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16][3] ), .I3(byte_transmit_counter[1]), 
            .O(n44355));
    defparam n44352_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37482 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n44346));
    defparam byte_transmit_counter_0__bdd_4_lut_37482.LUT_INIT = 16'he4aa;
    SB_LUT4 n44346_bdd_4_lut (.I0(n44346), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16]_c [2]), .I3(byte_transmit_counter[1]), 
            .O(n44349));
    defparam n44346_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n39185), .I3(n39184), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37477 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n44340));
    defparam byte_transmit_counter_0__bdd_4_lut_37477.LUT_INIT = 16'he4aa;
    SB_LUT4 n44340_bdd_4_lut (.I0(n44340), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16][1] ), .I3(byte_transmit_counter[1]), 
            .O(n44343));
    defparam n44340_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37472 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n44334));
    defparam byte_transmit_counter_0__bdd_4_lut_37472.LUT_INIT = 16'he4aa;
    SB_LUT4 n44334_bdd_4_lut (.I0(n44334), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16][0] ), .I3(byte_transmit_counter[1]), 
            .O(n44337));
    defparam n44334_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n39182), .I3(n39181), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n39179), .I3(n44259), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37467 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n44328));
    defparam byte_transmit_counter_0__bdd_4_lut_37467.LUT_INIT = 16'he4aa;
    SB_LUT4 n44328_bdd_4_lut (.I0(n44328), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n44331));
    defparam n44328_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37462 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n44322));
    defparam byte_transmit_counter_0__bdd_4_lut_37462.LUT_INIT = 16'he4aa;
    SB_LUT4 n44322_bdd_4_lut (.I0(n44322), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n44325));
    defparam n44322_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n39209), .I3(n39208), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37457 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n44316));
    defparam byte_transmit_counter_0__bdd_4_lut_37457.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n39212), .I3(n39211), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 n44316_bdd_4_lut (.I0(n44316), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n44319));
    defparam n44316_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37452 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n44310));
    defparam byte_transmit_counter_0__bdd_4_lut_37452.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1275 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4107), .O(n35429));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1275.LUT_INIT = 16'hffbf;
    SB_LUT4 n44310_bdd_4_lut (.I0(n44310), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n44313));
    defparam n44310_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37447 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n44304));
    defparam byte_transmit_counter_0__bdd_4_lut_37447.LUT_INIT = 16'he4aa;
    SB_LUT4 n44304_bdd_4_lut (.I0(n44304), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n44307));
    defparam n44304_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_127_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4124));   // verilog/coms.v(151[7:23])
    defparam equal_127_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_126_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4111));   // verilog/coms.v(151[7:23])
    defparam equal_126_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n96), .I3(n15879), .O(n38107));
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h0004;
    SB_LUT4 i22827_3_lut (.I0(\data_out_frame[16]_c [2]), .I1(\duty[10] ), 
            .I2(n13293), .I3(GND_net), .O(n17807));
    defparam i22827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1277 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [5]), .O(n8_adj_4095));
    defparam i1_2_lut_3_lut_4_lut_adj_1277.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1278 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [6]), .O(n34798));
    defparam i1_2_lut_3_lut_4_lut_adj_1278.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1279 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [7]), .O(n34796));
    defparam i1_2_lut_3_lut_4_lut_adj_1279.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1280 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [8]), .O(n34794));
    defparam i1_2_lut_3_lut_4_lut_adj_1280.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1281 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [9]), .O(n34792));
    defparam i1_2_lut_3_lut_4_lut_adj_1281.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1282 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [11]), .O(n34790));
    defparam i1_2_lut_3_lut_4_lut_adj_1282.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37442 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n44298));
    defparam byte_transmit_counter_0__bdd_4_lut_37442.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1283 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [12]), .O(n34788));
    defparam i1_2_lut_3_lut_4_lut_adj_1283.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1284 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [13]), .O(n34786));
    defparam i1_2_lut_3_lut_4_lut_adj_1284.LUT_INIT = 16'hfe00;
    SB_LUT4 n44298_bdd_4_lut (.I0(n44298), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n44301));
    defparam n44298_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1285 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [14]), .O(n34784));
    defparam i1_2_lut_3_lut_4_lut_adj_1285.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37437 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n44292));
    defparam byte_transmit_counter_0__bdd_4_lut_37437.LUT_INIT = 16'he4aa;
    SB_LUT4 n44292_bdd_4_lut (.I0(n44292), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n44295));
    defparam n44292_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13258_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18003));
    defparam i13258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37432 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n44286));
    defparam byte_transmit_counter_0__bdd_4_lut_37432.LUT_INIT = 16'he4aa;
    SB_LUT4 i13259_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18004));
    defparam i13259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n44286_bdd_4_lut (.I0(n44286), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n44289));
    defparam n44286_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13260_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18005));
    defparam i13260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [15]), .O(n34782));
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1287 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n35365));
    defparam i1_2_lut_3_lut_4_lut_adj_1287.LUT_INIT = 16'h0100;
    SB_LUT4 i13261_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18006));
    defparam i13261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13262_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18007));
    defparam i13262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13263_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18008));
    defparam i13263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_4_lut_4_lut_adj_1288 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n31898));
    defparam i2_4_lut_4_lut_4_lut_adj_1288.LUT_INIT = 16'h01ff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1289 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [16]), .O(n34780));
    defparam i1_2_lut_3_lut_4_lut_adj_1289.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1290 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4124), .O(n35428));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1290.LUT_INIT = 16'hffbf;
    SB_LUT4 i13264_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18009));
    defparam i13264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13265_3_lut_4_lut (.I0(n8_adj_4111), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18010));
    defparam i13265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13250_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n17995));
    defparam i13250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n24745), .O(n35435));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'hbfff;
    SB_LUT4 i13251_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n17996));
    defparam i13251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13252_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n17997));
    defparam i13252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2060_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3997));
    defparam i2060_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i13253_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n17998));
    defparam i13253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13254_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n17999));
    defparam i13254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1292 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [17]), .O(n34778));
    defparam i1_2_lut_3_lut_4_lut_adj_1292.LUT_INIT = 16'hfe00;
    SB_LUT4 i13255_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18000));
    defparam i13255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13256_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18001));
    defparam i13256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13257_3_lut_4_lut (.I0(n8_adj_4124), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18002));
    defparam i13257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20139_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15729), .I3(\FRAME_MATCHER.i [31]), .O(n2855));
    defparam i20139_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 mux_1068_i1_3_lut (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4377), .I3(GND_net), .O(n4378));
    defparam mux_1068_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1293 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [18]), .O(n8_adj_4097));
    defparam i1_2_lut_3_lut_4_lut_adj_1293.LUT_INIT = 16'hfe00;
    SB_LUT4 equal_123_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4123));
    defparam equal_123_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i21044_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n15879), .O(n25775));
    defparam i21044_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1294 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [19]), .O(n34776));
    defparam i1_2_lut_3_lut_4_lut_adj_1294.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1295 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [20]), .O(n8_adj_4099));
    defparam i1_2_lut_3_lut_4_lut_adj_1295.LUT_INIT = 16'hfe00;
    SB_LUT4 i20024_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24745));
    defparam i20024_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1296 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [21]), .O(n34774));
    defparam i1_2_lut_3_lut_4_lut_adj_1296.LUT_INIT = 16'hfe00;
    SB_LUT4 i20753_2_lut_3_lut_4_lut (.I0(n4_adj_4109), .I1(n1_c), .I2(n38_adj_4119), 
            .I3(\FRAME_MATCHER.state [22]), .O(n25478));
    defparam i20753_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1297 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [24]), .O(n8_adj_4101));
    defparam i1_2_lut_3_lut_4_lut_adj_1297.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1298 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [26]), .O(n8_adj_4103));
    defparam i1_2_lut_3_lut_4_lut_adj_1298.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1299 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [28]), .O(n34770));
    defparam i1_2_lut_3_lut_4_lut_adj_1299.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1300 (.I0(n4_adj_4109), .I1(n1_c), 
            .I2(n38_adj_4119), .I3(\FRAME_MATCHER.state [29]), .O(n34768));
    defparam i1_2_lut_3_lut_4_lut_adj_1300.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1301 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4110), .O(n35419));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1301.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1302 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n24745), .O(n35423));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1302.LUT_INIT = 16'hfbff;
    SB_LUT4 i20746_2_lut_3_lut_4_lut (.I0(n4_adj_4109), .I1(n1_c), .I2(n38_adj_4119), 
            .I3(\FRAME_MATCHER.state [31]), .O(n25470));
    defparam i20746_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1303 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4107), .O(n35420));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1303.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1304 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4124), .O(n35416));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1304.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1305 (.I0(n36742), .I1(n35947), .I2(\data_out_frame[17] [7]), 
            .I3(GND_net), .O(n35703));
    defparam i1_2_lut_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1306 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4111), .O(n35417));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1306.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_1068_i7_3_lut (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4377), .I3(GND_net), .O(n4384));
    defparam mux_1068_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i6_3_lut (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4377), .I3(GND_net), .O(n4383));
    defparam mux_1068_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1307 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4121), .O(n35421));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1307.LUT_INIT = 16'hfffb;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37427 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n44280));
    defparam byte_transmit_counter_0__bdd_4_lut_37427.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1308 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4122), .O(n35422));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1308.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1309 (.I0(n9), .I1(n24972), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n8_adj_4123), .O(n35418));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_4_lut_adj_1309.LUT_INIT = 16'hfffb;
    SB_LUT4 i5_3_lut_4_lut_adj_1310 (.I0(n35749), .I1(n10_adj_3893), .I2(\data_out_frame[17] [2]), 
            .I3(n15522), .O(n31104));
    defparam i5_3_lut_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1068_i22_3_lut (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4377), .I3(GND_net), .O(n4399));
    defparam mux_1068_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i21_3_lut (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4377), .I3(GND_net), .O(n4398));
    defparam mux_1068_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i20_3_lut (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4377), .I3(GND_net), .O(n4397));
    defparam mux_1068_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1311 (.I0(\data_out_frame[20] [3]), .I1(n31967), 
            .I2(n31208), .I3(\data_out_frame[20] [4]), .O(n35698));
    defparam i1_2_lut_3_lut_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1312 (.I0(n96), .I1(n99), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2388 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1312.LUT_INIT = 16'h1010;
    SB_LUT4 i13241_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n17986));
    defparam i13241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1068_i19_3_lut (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4377), .I3(GND_net), .O(n4396));
    defparam mux_1068_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i18_3_lut (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4377), .I3(GND_net), .O(n4395));
    defparam mux_1068_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1313 (.I0(n96), .I1(n99), .I2(n2086), .I3(\FRAME_MATCHER.state [3]), 
            .O(n2783));   // verilog/coms.v(126[12] 289[6])
    defparam i1_3_lut_4_lut_adj_1313.LUT_INIT = 16'h0f0e;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n19450));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2064_3_lut (.I0(n31_adj_4082), .I1(n31_adj_4125), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n12969));
    defparam i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_1197_i8_2_lut (.I0(Kp_23__N_946), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4126));   // verilog/coms.v(228[9:81])
    defparam equal_1197_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1315 (.I0(n16306), .I1(n8_adj_4126), .I2(n31979), 
            .I3(n16276), .O(n28_adj_4127));   // verilog/coms.v(228[9:81])
    defparam i12_4_lut_adj_1315.LUT_INIT = 16'hfdff;
    SB_LUT4 i10_4_lut_adj_1316 (.I0(n16919), .I1(n10_adj_4028), .I2(n16624), 
            .I3(n16974), .O(n26_adj_4128));   // verilog/coms.v(228[9:81])
    defparam i10_4_lut_adj_1316.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1317 (.I0(n16371), .I1(n31224), .I2(n16197), 
            .I3(n31222), .O(n27_adj_4129));   // verilog/coms.v(228[9:81])
    defparam i11_4_lut_adj_1317.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1318 (.I0(n11), .I1(n16557), .I2(n15_adj_4048), 
            .I3(n16218), .O(n25_adj_4130));   // verilog/coms.v(228[9:81])
    defparam i9_4_lut_adj_1318.LUT_INIT = 16'hfffe;
    SB_LUT4 i13274_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n18019));
    defparam i13274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1319 (.I0(n25_adj_4130), .I1(n27_adj_4129), .I2(n26_adj_4128), 
            .I3(n28_adj_4127), .O(n31_adj_4125));   // verilog/coms.v(228[9:81])
    defparam i15_4_lut_adj_1319.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1320 (.I0(\FRAME_MATCHER.state [1]), .I1(n31_adj_4125), 
            .I2(n13455), .I3(GND_net), .O(n4377));
    defparam i2_3_lut_adj_1320.LUT_INIT = 16'h0202;
    SB_LUT4 i4_4_lut_adj_1321 (.I0(n99), .I1(n12969), .I2(n13455), .I3(n19450), 
            .O(n38059));
    defparam i4_4_lut_adj_1321.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1068_i17_3_lut (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4377), .I3(GND_net), .O(n4394));
    defparam mux_1068_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n44280_bdd_4_lut (.I0(n44280), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n44283));
    defparam n44280_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13275_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n18020));
    defparam i13275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1322 (.I0(tx_active), .I1(r_SM_Main_2__N_3323[0]), 
            .I2(tx_transmit_N_3220), .I3(n10454), .O(n13142));
    defparam i1_2_lut_3_lut_4_lut_adj_1322.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n25775), .I2(n31898), 
            .I3(GND_net), .O(n38154));
    defparam i3_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\FRAME_MATCHER.state[0] ), .I1(n13455), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4131));
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1324 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state_31__N_2490 [3]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n38182));
    defparam i2_3_lut_adj_1324.LUT_INIT = 16'h0808;
    SB_LUT4 i2_4_lut_adj_1325 (.I0(\FRAME_MATCHER.state [2]), .I1(n12969), 
            .I2(n38182), .I3(n4_adj_4131), .O(n36130));
    defparam i2_4_lut_adj_1325.LUT_INIT = 16'h5072;
    SB_LUT4 i2_4_lut_adj_1326 (.I0(n3301), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n36130), .I3(n25775), .O(n36732));
    defparam i2_4_lut_adj_1326.LUT_INIT = 16'h5011;
    SB_LUT4 i13276_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n18021));
    defparam i13276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1327 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n13_adj_3984), .I3(n13142), 
            .O(n131));
    defparam i1_2_lut_3_lut_4_lut_adj_1327.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1328 (.I0(n16218), .I1(\data_in_frame[6] [4]), 
            .I2(n11), .I3(\data_in_frame[10] [6]), .O(n36092));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1329 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(n5_c), .O(Kp_23__N_893));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1330 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(n35667), .O(n31190));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i32243_2_lut_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n31_adj_4082), .I3(GND_net), .O(n39023));
    defparam i32243_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13277_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n18022));
    defparam i13277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [7]), .O(n6_adj_4050));   // verilog/coms.v(69[16:69])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1331 (.I0(\data_in_frame[7] [2]), .I1(n31190), 
            .I2(\data_in_frame[4] [7]), .I3(n35741), .O(n8_adj_4049));
    defparam i3_3_lut_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1332 (.I0(n13_adj_3984), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n97));
    defparam i1_2_lut_3_lut_adj_1332.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut_4_lut_adj_1333 (.I0(\data_in_frame[12] [5]), .I1(n10_adj_4038), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[6] [1]), .O(n35535));   // verilog/coms.v(70[16:41])
    defparam i5_3_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1334 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[1] [3]), .O(Kp_23__N_946));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1335 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[13] [0]), .O(n14_adj_4034));
    defparam i5_3_lut_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1336 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[10] [1]), 
            .I2(n10_adj_4032), .I3(\data_in_frame[9] [6]), .O(n35601));
    defparam i5_3_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1337 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[14] [5]), 
            .I2(\data_in_frame[14] [4]), .I3(GND_net), .O(n35688));
    defparam i1_2_lut_3_lut_adj_1337.LUT_INIT = 16'h9696;
    SB_LUT4 i13278_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n18023));
    defparam i13278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(\data_in_frame[6] [2]), .I1(n10_adj_4028), 
            .I2(n35972), .I3(GND_net), .O(n35888));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_LUT4 i13279_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n18024));
    defparam i13279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13280_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n18025));
    defparam i13280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13281_3_lut_4_lut (.I0(n8_adj_4122), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n18026));
    defparam i13281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_124_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4122));   // verilog/coms.v(151[7:23])
    defparam equal_124_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(n36742), .I1(n35947), .I2(n1640), 
            .I3(GND_net), .O(n35700));
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 equal_125_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4121));   // verilog/coms.v(151[7:23])
    defparam equal_125_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in[2] [7]), .I1(n10_adj_4016), .I2(\data_in[3] [4]), 
            .I3(\data_in[3] [0]), .O(n15_adj_4027));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_4_lut_adj_1340 (.I0(n16394), .I1(n35577), .I2(\data_out_frame[10] [2]), 
            .I3(\data_out_frame[10] [0]), .O(n31090));
    defparam i2_3_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_adj_4018));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n35630), .I1(\data_in_frame[9] [4]), 
            .I2(n36074), .I3(GND_net), .O(n31488));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(n31190), .I1(\data_in_frame[4] [7]), 
            .I2(n36098), .I3(GND_net), .O(n35798));
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_LUT4 i13234_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n17979));
    defparam i13234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37422 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n44274));
    defparam byte_transmit_counter_0__bdd_4_lut_37422.LUT_INIT = 16'he4aa;
    SB_LUT4 n44274_bdd_4_lut (.I0(n44274), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n44277));
    defparam n44274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13235_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n17980));
    defparam i13235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1344 (.I0(n21), .I1(n19_adj_3923), .I2(n20), 
            .I3(n16898), .O(n36104));
    defparam i1_2_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i13236_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n17981));
    defparam i13236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1345 (.I0(n21), .I1(n19_adj_3923), .I2(n20), 
            .I3(\data_out_frame[11] [7]), .O(n35478));
    defparam i1_2_lut_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4132));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34822_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41676));   // verilog/coms.v(104[34:55])
    defparam i34822_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4133));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32376_4_lut (.I0(n19_adj_4132), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39229));
    defparam i32376_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32377_3_lut (.I0(n44379), .I1(n39229), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39230));
    defparam i32377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32330_4_lut (.I0(n5_adj_4133), .I1(n41676), .I2(n41084), 
            .I3(\byte_transmit_counter[0] ), .O(n39183));
    defparam i32330_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i32332_4_lut (.I0(n39183), .I1(n39230), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n39185));
    defparam i32332_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32331_3_lut (.I0(n44283), .I1(n44277), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39184));
    defparam i32331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n4_adj_3979));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4134));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35535_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42389));   // verilog/coms.v(104[34:55])
    defparam i35535_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4135));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32373_4_lut (.I0(n19_adj_4134), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39226));
    defparam i32373_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32374_3_lut (.I0(n44373), .I1(n39226), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39227));
    defparam i32374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32327_4_lut (.I0(n5_adj_4135), .I1(n42389), .I2(n41084), 
            .I3(\byte_transmit_counter[0] ), .O(n39180));
    defparam i32327_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i32329_4_lut (.I0(n39180), .I1(n39227), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n39182));
    defparam i32329_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32328_3_lut (.I0(n44295), .I1(n44289), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39181));
    defparam i32328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1347 (.I0(n31190), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [3]), .I3(n31224), .O(n35762));
    defparam i1_2_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4136));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32370_4_lut (.I0(n19_adj_4136), .I1(\data_out_frame[22] [5]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39223));
    defparam i32370_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n41668));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4137));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32371_3_lut (.I0(n44367), .I1(n39223), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39224));
    defparam i32371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32324_4_lut (.I0(n5_adj_4137), .I1(\byte_transmit_counter[0] ), 
            .I2(n41084), .I3(n41668), .O(n39177));
    defparam i32324_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i32326_4_lut (.I0(n39177), .I1(n39224), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n39179));
    defparam i32326_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(\data_in_frame[6] [4]), .I1(n11), 
            .I2(n36026), .I3(GND_net), .O(n6_adj_4017));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4138));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4139));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4140));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32367_4_lut (.I0(n19_adj_4138), .I1(\data_out_frame[22] [4]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39220));
    defparam i32367_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1349 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[7] [0]), .I3(n35568), .O(n36026));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i32368_3_lut (.I0(n44361), .I1(n39220), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39221));
    defparam i32368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32357_3_lut (.I0(n5_adj_4140), .I1(n6_adj_4139), .I2(n41084), 
            .I3(GND_net), .O(n39210));
    defparam i32357_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32359_4_lut (.I0(n39210), .I1(n39221), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n39212));
    defparam i32359_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32358_3_lut (.I0(n44307), .I1(n44301), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39211));
    defparam i32358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1350 (.I0(\data_in_frame[6] [7]), .I1(n16919), 
            .I2(Kp_23__N_893), .I3(\data_in_frame[4] [6]), .O(n35568));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(n16624), .I1(\data_in_frame[14] [3]), 
            .I2(\data_in_frame[14] [2]), .I3(GND_net), .O(n6_adj_4014));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n35829));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4141));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4142));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(n31802), .I3(GND_net), .O(n12_adj_3914));   // verilog/coms.v(73[16:27])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4143));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32364_4_lut (.I0(n19_adj_4141), .I1(\data_out_frame[22] [3]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39217));
    defparam i32364_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n35513));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i32365_3_lut (.I0(n44355), .I1(n39217), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39218));
    defparam i32365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32354_3_lut (.I0(n5_adj_4143), .I1(n6_adj_4142), .I2(n41084), 
            .I3(GND_net), .O(n39207));
    defparam i32354_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32356_4_lut (.I0(n39207), .I1(n39218), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n39209));
    defparam i32356_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32355_3_lut (.I0(n44319), .I1(n44313), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39208));
    defparam i32355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(n35630), .I1(n35884), .I2(\data_in_frame[13] [7]), 
            .I3(\data_in_frame[13] [6]), .O(n35775));
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i32397_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39250));
    defparam i32397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37417 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n44262));
    defparam byte_transmit_counter_0__bdd_4_lut_37417.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4144));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32340_4_lut (.I0(n19_adj_4144), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39193));
    defparam i32340_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n44262_bdd_4_lut (.I0(n44262), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n44265));
    defparam n44262_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i32398_4_lut (.I0(n39250), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n39251));
    defparam i32398_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i32396_3_lut (.I0(\data_out_frame[4][2] ), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39249));
    defparam i32396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35946_3_lut (.I0(n44325), .I1(n44265), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n42800));
    defparam i35946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32341_3_lut (.I0(n44349), .I1(n39193), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39194));
    defparam i32341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36219_3_lut (.I0(n39204), .I1(n42800), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n43073));   // verilog/coms.v(104[34:55])
    defparam i36219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36220_4_lut (.I0(n43073), .I1(n39194), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam i36220_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n39273), .I2(n39274), .I3(byte_transmit_counter[2]), .O(n44256));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4][1] ), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n36068));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4145));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32337_4_lut (.I0(n19_adj_4145), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n39190));
    defparam i32337_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32389_4_lut (.I0(\data_out_frame[6] [1]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n39242));
    defparam i32389_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i32387_3_lut (.I0(\data_out_frame[4][1] ), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n39240));
    defparam i32387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35950_3_lut (.I0(n44331), .I1(n44253), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n42804));
    defparam i35950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n44256_bdd_4_lut (.I0(n44256), .I1(n39271), .I2(n39270), .I3(byte_transmit_counter[2]), 
            .O(n44259));
    defparam n44256_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1356 (.I0(\data_in_frame[6] [2]), .I1(n10_adj_4028), 
            .I2(\data_in_frame[8] [4]), .I3(n16197), .O(n36053));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i32338_3_lut (.I0(n44343), .I1(n39190), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39191));
    defparam i32338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36217_3_lut (.I0(n39201), .I1(n42804), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n43071));   // verilog/coms.v(104[34:55])
    defparam i36217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36218_4_lut (.I0(n43071), .I1(n39191), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam i36218_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1357 (.I0(\data_in_frame[15] [6]), .I1(n16173), 
            .I2(n31202), .I3(\data_in_frame[18] [0]), .O(n31962));
    defparam i1_2_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37408 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n44250));
    defparam byte_transmit_counter_0__bdd_4_lut_37408.LUT_INIT = 16'he4aa;
    SB_LUT4 i37374_1_lut_4_lut (.I0(n24660), .I1(n25346), .I2(n13_adj_3984), 
            .I3(\FRAME_MATCHER.i_31__N_2388 ), .O(n44226));
    defparam i37374_1_lut_4_lut.LUT_INIT = 16'h00fd;
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n13_adj_3984), .I3(GND_net), .O(n61));
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'hfbfb;
    SB_LUT4 i21015_3_lut_4_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[3]), 
            .O(n25745));
    defparam i21015_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 n44250_bdd_4_lut (.I0(n44250), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n44253));
    defparam n44250_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[15] [3]), .I3(GND_net), .O(n35500));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4][1] ), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n1173));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(n43489), .I1(n35507), .I2(\data_out_frame[9] [5]), 
            .I3(GND_net), .O(n35907));   // verilog/coms.v(95[12:26])
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37399 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n44244));
    defparam byte_transmit_counter_0__bdd_4_lut_37399.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(n43489), .I1(n35507), .I2(n36029), 
            .I3(GND_net), .O(n35910));   // verilog/coms.v(95[12:26])
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n35507));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(n16974), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[9] [0]), .O(n35574));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\FRAME_MATCHER.state [31]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35389));
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n13_adj_3984), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2390 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\FRAME_MATCHER.state [30]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35405));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h8888;
    SB_LUT4 i20249_2_lut_3_lut (.I0(n2086), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n24972));
    defparam i20249_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_1368 (.I0(\FRAME_MATCHER.state [29]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35396));
    defparam i1_2_lut_adj_1368.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1369 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n38135));
    defparam i2_3_lut_4_lut_adj_1369.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\FRAME_MATCHER.state [28]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35402));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h8888;
    SB_LUT4 i32283_3_lut_4_lut (.I0(n13455), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[2] [2]), .O(n39063));
    defparam i32283_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\FRAME_MATCHER.state [27]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35399));
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h8888;
    SB_LUT4 i32281_3_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [3]), 
            .I2(n35519), .I3(n35723), .O(n39061));
    defparam i32281_3_lut_4_lut.LUT_INIT = 16'h7dbe;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\FRAME_MATCHER.state [25]), .I1(n35449), 
            .I2(GND_net), .I3(GND_net), .O(n34680));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1373 (.I0(n13_adj_3984), .I1(n35386), .I2(\FRAME_MATCHER.state [25]), 
            .I3(n7_adj_4120), .O(n37102));
    defparam i2_4_lut_adj_1373.LUT_INIT = 16'h5040;
    SB_LUT4 i1_2_lut_adj_1374 (.I0(\FRAME_MATCHER.state [23]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35408));
    defparam i1_2_lut_adj_1374.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1375 (.I0(\FRAME_MATCHER.state [21]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35393));
    defparam i1_2_lut_adj_1375.LUT_INIT = 16'h8888;
    SB_LUT4 i7_3_lut_4_lut_adj_1376 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[5] [4]), 
            .I2(n35654), .I3(n36023), .O(n20_adj_3925));   // verilog/coms.v(95[12:26])
    defparam i7_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_adj_1377 (.I0(\data_out_frame[9] [5]), .I1(n31288), 
            .I2(\data_out_frame[10] [1]), .I3(GND_net), .O(n16_adj_3924));   // verilog/coms.v(95[12:26])
    defparam i3_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1378 (.I0(\FRAME_MATCHER.state [19]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35395));
    defparam i1_2_lut_adj_1378.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1379 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[9] [1]), .I3(\data_out_frame[9] [2]), .O(n16993));
    defparam i1_2_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1380 (.I0(n16394), .I1(n35577), .I2(n35478), 
            .I3(\data_out_frame[8] [1]), .O(n31288));
    defparam i1_2_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1381 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n35846));
    defparam i1_2_lut_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(n1238), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4][1] ), .I3(\data_out_frame[6] [4]), .O(n36023));
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(\FRAME_MATCHER.state [17]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35394));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h8888;
    SB_LUT4 i13266_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18011));
    defparam i13266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1384 (.I0(\FRAME_MATCHER.state [16]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35409));
    defparam i1_2_lut_adj_1384.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1385 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(n16535), .I3(\data_out_frame[5] [3]), .O(n35577));
    defparam i2_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\FRAME_MATCHER.state [15]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35401));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n16535));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1388 (.I0(\FRAME_MATCHER.state [14]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35404));
    defparam i1_2_lut_adj_1388.LUT_INIT = 16'h8888;
    SB_LUT4 n44244_bdd_4_lut (.I0(n44244), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n44247));
    defparam n44244_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13267_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18012));
    defparam i13267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n35654));
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(n36104), .I3(GND_net), .O(n36029));
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(\FRAME_MATCHER.state [13]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35398));
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h8888;
    SB_LUT4 i36635_2_lut_3_lut (.I0(\data_out_frame[5] [4]), .I1(n35654), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n43489));   // verilog/coms.v(95[12:26])
    defparam i36635_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1392 (.I0(\FRAME_MATCHER.state [12]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35407));
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\FRAME_MATCHER.state [11]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35392));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1394 (.I0(\FRAME_MATCHER.state [2]), .I1(n35448), 
            .I2(n35383), .I3(\FRAME_MATCHER.state [1]), .O(n35449));
    defparam i1_4_lut_adj_1394.LUT_INIT = 16'hccdc;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\FRAME_MATCHER.state [10]), .I1(n35449), 
            .I2(GND_net), .I3(GND_net), .O(n34720));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1396 (.I0(\FRAME_MATCHER.state [10]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35390));
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_4_lut_adj_1397 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[13] [6]), .I3(\data_out_frame[11] [6]), 
            .O(n10_adj_3919));   // verilog/coms.v(69[16:27])
    defparam i2_2_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1398 (.I0(\FRAME_MATCHER.state [9]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35391));
    defparam i1_2_lut_adj_1398.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_4_lut_adj_1399 (.I0(\data_out_frame[9] [4]), .I1(n14104), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[14] [1]), .O(n8_adj_3918));   // verilog/coms.v(83[17:28])
    defparam i3_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i13268_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18013));
    defparam i13268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(\FRAME_MATCHER.state [8]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35406));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [3]), .O(n14104));
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i13269_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18014));
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\FRAME_MATCHER.state [7]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35397));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[13] [6]), .I3(GND_net), .O(n36044));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i13270_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18015));
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\FRAME_MATCHER.state [6]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35403));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n35487));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_out_frame[20] [7]), .I1(n30877), 
            .I2(n36047), .I3(GND_net), .O(n6_adj_3910));
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1407 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4][0] ), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n16711));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_1407.LUT_INIT = 16'h9696;
    SB_LUT4 i13237_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n17982));
    defparam i13237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1408 (.I0(\data_out_frame[19] [0]), .I1(n32004), 
            .I2(\data_out_frame[19] [1]), .I3(n31802), .O(n10_adj_3908));
    defparam i2_2_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4146));
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1410 (.I0(n13_adj_3984), .I1(n13197), .I2(n7_adj_4120), 
            .I3(n4_adj_4146), .O(n35388));
    defparam i1_4_lut_adj_1410.LUT_INIT = 16'h5450;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n16042));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\FRAME_MATCHER.state [4]), .I1(n35388), 
            .I2(GND_net), .I3(GND_net), .O(n35400));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h8888;
    SB_LUT4 i13271_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18016));
    defparam i13271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1413 (.I0(n3741), .I1(n10454), .I2(GND_net), 
            .I3(GND_net), .O(n13197));   // verilog/coms.v(248[6] 250[9])
    defparam i1_2_lut_adj_1413.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1414 (.I0(n10454), .I1(n2778), .I2(GND_net), 
            .I3(GND_net), .O(n1_c));
    defparam i1_2_lut_adj_1414.LUT_INIT = 16'h8888;
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(n28_adj_3901), .I3(\data_out_frame[8] [3]), .O(n32));
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1415 (.I0(\FRAME_MATCHER.i_31__N_2390 ), .I1(n10454), 
            .I2(n2855), .I3(GND_net), .O(n38_adj_4119));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1415.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_adj_1416 (.I0(\FRAME_MATCHER.state [3]), .I1(n38_adj_4119), 
            .I2(n4_adj_4109), .I3(n131), .O(n7_adj_4147));
    defparam i1_4_lut_adj_1416.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_1417 (.I0(n6_adj_3983), .I1(n7_adj_4147), .I2(n15862), 
            .I3(n104), .O(n34894));
    defparam i1_4_lut_adj_1417.LUT_INIT = 16'hccce;
    SB_LUT4 i1_4_lut_adj_1418 (.I0(\FRAME_MATCHER.state [3]), .I1(n1_c), 
            .I2(n13_adj_3984), .I3(n35386), .O(n34722));
    defparam i1_4_lut_adj_1418.LUT_INIT = 16'h8a88;
    SB_LUT4 i13272_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18017));
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[5] [7]), .I3(n35542), .O(n36011));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1420 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(n31228), .I3(n32092), .O(n10_adj_4148));
    defparam i4_4_lut_adj_1420.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1421 (.I0(n31684), .I1(n10_adj_4148), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n37234));
    defparam i5_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1422 (.I0(n31208), .I1(\data_out_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n31228));
    defparam i1_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1423 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(n10_adj_3899), .I3(\data_out_frame[9] [1]), .O(n15502));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(n16234), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n18));
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1425 (.I0(n15497), .I1(n35561), .I2(n37462), 
            .I3(GND_net), .O(n37006));
    defparam i2_3_lut_adj_1425.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1426 (.I0(\data_out_frame[20] [1]), .I1(n35539), 
            .I2(GND_net), .I3(GND_net), .O(n35540));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1426.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1427 (.I0(\data_out_frame[19] [7]), .I1(n31140), 
            .I2(n35552), .I3(n6_adj_4118), .O(n15497));
    defparam i4_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1428 (.I0(n15497), .I1(n35817), .I2(n31967), 
            .I3(GND_net), .O(n37148));
    defparam i2_3_lut_adj_1428.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1429 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[18] [0]), .I3(GND_net), .O(n35867));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1430 (.I0(n35553), .I1(n35759), .I2(n32094), 
            .I3(\data_out_frame[18] [0]), .O(n37462));
    defparam i3_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1431 (.I0(n32079), .I1(n35555), .I2(n35484), 
            .I3(n32092), .O(n16348));
    defparam i3_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i13238_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n17983));
    defparam i13238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13273_3_lut_4_lut (.I0(n8_adj_4121), .I1(n35439), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18018));
    defparam i13273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\data_out_frame[18] [1]), .I1(n35552), 
            .I2(GND_net), .I3(GND_net), .O(n35553));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1433 (.I0(n35553), .I1(n32092), .I2(\data_out_frame[18] [2]), 
            .I3(n6_adj_4117), .O(n31967));
    defparam i4_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i13239_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n17984));
    defparam i13239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n35598));
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n16234));
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1436 (.I0(\data_out_frame[19] [5]), .I1(n2106), 
            .I2(n35811), .I3(GND_net), .O(n14_adj_4149));
    defparam i5_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1437 (.I0(n16348), .I1(n32004), .I2(n37462), 
            .I3(\data_out_frame[19] [4]), .O(n15_adj_4150));
    defparam i6_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i13240_3_lut_4_lut (.I0(n8_adj_4110), .I1(n35439), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n17985));
    defparam i13240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1438 (.I0(n15_adj_4150), .I1(n35960), .I2(n14_adj_4149), 
            .I3(\data_out_frame[19] [1]), .O(n35817));
    defparam i8_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1439 (.I0(n35700), .I1(n32012), .I2(\data_out_frame[19] [6]), 
            .I3(\data_out_frame[17] [7]), .O(n37421));
    defparam i3_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1440 (.I0(n37421), .I1(\data_out_frame[20] [0]), 
            .I2(n35867), .I3(n16723), .O(n35539));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1441 (.I0(n35539), .I1(n35817), .I2(n31967), 
            .I3(GND_net), .O(n37704));
    defparam i2_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_out_frame[18] [3]), .I1(n16704), 
            .I2(GND_net), .I3(GND_net), .O(n35555));
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1443 (.I0(\data_out_frame[11] [3]), .I1(n31226), 
            .I2(n1238), .I3(n35598), .O(n22_adj_4151));   // verilog/coms.v(69[16:27])
    defparam i9_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1444 (.I0(n35950), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[11] [5]), .I3(n35765), .O(n21_adj_4152));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[15] [7]), .I3(n14104), .O(n14_adj_4153));
    defparam i5_3_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1446 (.I0(n35878), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[5] [0]), .I3(n14_adj_4104), .O(n23));   // verilog/coms.v(69[16:27])
    defparam i10_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(\data_out_frame[16][0] ), .I1(n23), .I2(n21_adj_4152), 
            .I3(n22_adj_4151), .O(n32094));
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1448 (.I0(n32094), .I1(n35555), .I2(\data_out_frame[18] [2]), 
            .I3(GND_net), .O(n31208));
    defparam i2_3_lut_adj_1448.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35561));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(n30880), .I1(\data_out_frame[15] [0]), 
            .I2(n1640), .I3(GND_net), .O(n31142));
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1451 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [3]), 
            .I2(n35561), .I3(n6_adj_4108), .O(n2106));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(\data_out_frame[15] [6]), .I1(n36742), 
            .I2(GND_net), .I3(GND_net), .O(n32012));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(n16477), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35759));
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[13] [7]), 
            .I2(n16993), .I3(GND_net), .O(n36056));
    defparam i1_2_lut_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1455 (.I0(\data_out_frame[16] [7]), .I1(n35749), 
            .I2(n10_adj_3893), .I3(n31150), .O(n7_c));
    defparam i2_2_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1456 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4154));
    defparam i4_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1457 (.I0(n36035), .I1(n16234), .I2(\data_out_frame[14] [0]), 
            .I3(n35978), .O(n15_adj_4155));
    defparam i6_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(\data_out_frame[16][1] ), .I1(n15_adj_4155), 
            .I2(n13_adj_4154), .I3(n14_adj_4153), .O(n32092));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(n30880), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n31140));
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[17] [4]), 
            .I2(n31288), .I3(\data_out_frame[18] [5]), .O(n52));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n16487), .I1(n32092), .I2(n36742), .I3(n30900), 
            .O(n50));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n36089), .I1(n35684), .I2(n36032), .I3(n43489), 
            .O(n51));
    defparam i21_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1460 (.I0(n35619), .I1(n36104), .I2(\data_out_frame[16][3] ), 
            .I3(n35913), .O(n49));
    defparam i19_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1461 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[19] [3]), 
            .I2(n1395), .I3(\data_out_frame[19] [7]), .O(n46));
    defparam i16_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1462 (.I0(\data_out_frame[19] [6]), .I1(n36056), 
            .I2(n16477), .I3(\data_out_frame[18] [1]), .O(n48_adj_4156));
    defparam i18_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1463 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[18] [7]), 
            .I2(n1829), .I3(\data_out_frame[18] [6]), .O(n47));
    defparam i17_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut_adj_1464 (.I0(n49), .I1(n51), .I2(n50), .I3(n52), 
            .O(n58));
    defparam i28_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut (.I0(\data_out_frame[18] [0]), .I1(n46), .I2(\data_out_frame[17] [1]), 
            .I3(GND_net), .O(n53));
    defparam i23_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i29_4_lut_adj_1465 (.I0(n53), .I1(n58), .I2(n47), .I3(n48_adj_4156), 
            .O(n35811));
    defparam i29_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1466 (.I0(n35811), .I1(n31140), .I2(\data_out_frame[17] [4]), 
            .I3(n35756), .O(n15_adj_4157));
    defparam i6_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1467 (.I0(n15_adj_4157), .I1(n31208), .I2(n14_adj_4114), 
            .I3(\data_out_frame[17] [3]), .O(n37659));
    defparam i8_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(\data_out_frame[19] [4]), .I1(n32044), 
            .I2(GND_net), .I3(GND_net), .O(n35616));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16723));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1470 (.I0(n31150), .I1(n16723), .I2(\data_out_frame[15] [3]), 
            .I3(n35616), .O(n10_adj_4158));
    defparam i4_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1471 (.I0(n31142), .I1(n10_adj_4158), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n37040));
    defparam i5_3_lut_adj_1471.LUT_INIT = 16'h9696;
    uart_tx tx (.VCC_net(VCC_net), .GND_net(GND_net), .clk32MHz(clk32MHz), 
            .n17466(n17466), .\r_Clock_Count[6] (\r_Clock_Count[6] ), .n17463(n17463), 
            .\r_Clock_Count[7] (\r_Clock_Count[7] ), .n17481(n17481), .\r_Clock_Count[1] (\r_Clock_Count[1] ), 
            .n17512(n17512), .r_Bit_Index({r_Bit_Index}), .n17509(n17509), 
            .n18130(n18130), .r_SM_Main({r_SM_Main}), .n18105(n18105), 
            .tx_data({tx_data}), .tx_o(tx_o), .tx_enable(tx_enable), .tx_active(tx_active), 
            .\r_SM_Main_2__N_3323[0] (r_SM_Main_2__N_3323[0]), .n25346(n25346), 
            .n19634(n19634), .n17529(n17529), .n17528(n17528), .n541(n541), 
            .n314(n314), .n315(n315), .n320(n320), .o_Tx_Serial_N_3351(o_Tx_Serial_N_3351), 
            .n17108(n17108), .n4683(n4683), .n17186(n17186), .n17330(n17330)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.n35270(n35270), .r_Clock_Count({r_Clock_Count}), .GND_net(GND_net), 
            .n35268(n35268), .n35273(n35273), .VCC_net(VCC_net), .rx_data_ready(rx_data_ready), 
            .clk32MHz(clk32MHz), .n18165(n18165), .rx_data({rx_data}), 
            .n35086(n35086), .n35088(n35088), .n35090(n35090), .n35000(n35000), 
            .n34912(n34912), .n34804(n34804), .n34716(n34716), .n17566(n17566), 
            .r_Bit_Index({r_Bit_Index_adj_14}), .n17569(n17569), .n35004(n35004), 
            .n18111(n18111), .n25741(n25741), .r_SM_Main({r_SM_Main_adj_15}), 
            .n35269(n35269), .r_Rx_Data(r_Rx_Data), .n35272(n35272), .PIN_13_N_105(PIN_13_N_105), 
            .n35275(n35275), .n35276(n35276), .n35271(n35271), .n35274(n35274), 
            .n41248(n41248), .n41247(n41247), .n17576(n17576), .n17575(n17575), 
            .n17574(n17574), .n17573(n17573), .n17572(n17572), .n17571(n17571), 
            .n17570(n17570), .n17527(n17527), .n17180(n17180), .n17321(n17321), 
            .n4661(n4661), .n35374(n35374), .n25555(n25555), .n1(n1), 
            .n24764(n24764), .n4(n4), .n4_adj_1(n4_adj_12), .n15912(n15912), 
            .n15917(n15917), .n4_adj_2(n4_adj_13), .n6(n6), .n44844(n44844)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (VCC_net, GND_net, clk32MHz, n17466, \r_Clock_Count[6] , 
            n17463, \r_Clock_Count[7] , n17481, \r_Clock_Count[1] , 
            n17512, r_Bit_Index, n17509, n18130, r_SM_Main, n18105, 
            tx_data, tx_o, tx_enable, tx_active, \r_SM_Main_2__N_3323[0] , 
            n25346, n19634, n17529, n17528, n541, n314, n315, 
            n320, o_Tx_Serial_N_3351, n17108, n4683, n17186, n17330) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input VCC_net;
    input GND_net;
    input clk32MHz;
    input n17466;
    output \r_Clock_Count[6] ;
    input n17463;
    output \r_Clock_Count[7] ;
    input n17481;
    output \r_Clock_Count[1] ;
    input n17512;
    output [2:0]r_Bit_Index;
    input n17509;
    input n18130;
    output [2:0]r_SM_Main;
    input n18105;
    input [7:0]tx_data;
    output tx_o;
    output tx_enable;
    output tx_active;
    input \r_SM_Main_2__N_3323[0] ;
    output n25346;
    output n19634;
    input n17529;
    input n17528;
    output n541;
    output n314;
    output n315;
    output n320;
    output o_Tx_Serial_N_3351;
    output n17108;
    output n4683;
    output n17186;
    output n17330;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n28526, n17472, n17469, n17460, n17478, n17475, n18168, 
        n13276;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n44388, n44391, n19635, n35074, n44764, n41252, n28533, 
        n28532, n28531, n41250, n28530, n41251, n28529, n41253, 
        n28528;
    wire [8:0]n312;
    
    wire n28527, n41254, n44271, n8896, n25512, n12, n10, n38070, 
        n44268;
    
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n28526));
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n17472));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n17469));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(clk32MHz), .D(n17466));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(\r_Clock_Count[7] ), .C(clk32MHz), .D(n17463));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n17460));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(\r_Clock_Count[1] ), .C(clk32MHz), .D(n17481));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17478));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n17475));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17512));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17509));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n18168));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n18130));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18105));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i18193_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(tx_enable));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i18193_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20623_2_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n25346));
    defparam i20623_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13276), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n44388));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n44388_bdd_4_lut (.I0(n44388), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n44391));
    defparam n44388_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n19634), .I2(GND_net), .I3(GND_net), 
            .O(n19635));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n35074));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n17529));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n17528));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n44764));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(n541), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n28533), .O(n41252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(\r_Clock_Count[7] ), .I2(GND_net), 
            .I3(n28532), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_9 (.CI(n28532), .I0(\r_Clock_Count[7] ), .I1(GND_net), 
            .CO(n28533));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(\r_Clock_Count[6] ), .I2(GND_net), 
            .I3(n28531), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n28531), .I0(\r_Clock_Count[6] ), .I1(GND_net), 
            .CO(n28532));
    SB_LUT4 add_59_7_lut (.I0(n541), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n28530), .O(n41250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_7 (.CI(n28530), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n28531));
    SB_LUT4 add_59_6_lut (.I0(n541), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n28529), .O(n41251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_6 (.CI(n28529), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n28530));
    SB_LUT4 add_59_5_lut (.I0(n541), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n28528), .O(n41253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_5 (.CI(n28528), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n28529));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n28527), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n28527), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n28528));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(\r_Clock_Count[1] ), .I2(GND_net), 
            .I3(n28526), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n28526), .I0(\r_Clock_Count[1] ), .I1(GND_net), 
            .CO(n28527));
    SB_LUT4 add_59_2_lut (.I0(n541), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n41254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i22470_3_lut (.I0(r_Clock_Count[0]), .I1(n41254), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n18168));
    defparam i22470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3323[0] ), 
            .I3(r_SM_Main[2]), .O(n13276));   // verilog/uart_tx.v(31[16:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(n19634), 
            .I3(r_SM_Main[2]), .O(n541));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff0e;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(n19634), .O(n44764));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i2108940_i1_3_lut (.I0(n44391), .I1(n44271), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3351));
    defparam i2108940_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_860 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n8896));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n8896), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n19635), .O(n17108));
    defparam i2_4_lut.LUT_INIT = 16'h3202;
    SB_LUT4 i29_4_lut (.I0(\r_SM_Main_2__N_3323[0] ), .I1(n25512), .I2(r_SM_Main[1]), 
            .I3(n19634), .O(n12));   // verilog/uart_tx.v(31[16:25])
    defparam i29_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n12), .I2(n19634), .I3(r_SM_Main[0]), 
            .O(n35074));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1304_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4683));   // verilog/uart_tx.v(98[36:51])
    defparam i1304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n25512));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_861 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n19634), .O(n17186));
    defparam i2_4_lut_adj_861.LUT_INIT = 16'h1101;
    SB_LUT4 i12585_3_lut (.I0(n17186), .I1(r_SM_Main[1]), .I2(n25512), 
            .I3(GND_net), .O(n17330));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12585_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i22456_3_lut (.I0(r_Clock_Count[3]), .I1(n41253), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17475));
    defparam i22456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_862 (.I0(n541), .I1(r_Clock_Count[2]), .I2(n312[2]), 
            .I3(r_SM_Main[2]), .O(n17478));
    defparam i1_4_lut_adj_862.LUT_INIT = 16'h88a0;
    SB_LUT4 i22443_3_lut (.I0(r_Clock_Count[8]), .I1(n41252), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17460));
    defparam i22443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(\r_Clock_Count[1] ), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[5]), 
            .I3(r_Clock_Count[2]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[4]), .I1(n10), .I2(r_Clock_Count[0]), 
            .I3(GND_net), .O(n38070));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut_adj_863 (.I0(r_Clock_Count[8]), .I1(\r_Clock_Count[6] ), 
            .I2(\r_Clock_Count[7] ), .I3(n38070), .O(n19634));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut_adj_863.LUT_INIT = 16'hfffe;
    SB_LUT4 i22396_3_lut (.I0(r_Clock_Count[5]), .I1(n41250), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17469));
    defparam i22396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22409_3_lut (.I0(r_Clock_Count[4]), .I1(n41251), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17472));
    defparam i22409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_37512 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n44268));
    defparam r_Bit_Index_0__bdd_4_lut_37512.LUT_INIT = 16'he4aa;
    SB_LUT4 n44268_bdd_4_lut (.I0(n44268), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n44271));
    defparam n44268_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n35270, r_Clock_Count, GND_net, n35268, n35273, VCC_net, 
            rx_data_ready, clk32MHz, n18165, rx_data, n35086, n35088, 
            n35090, n35000, n34912, n34804, n34716, n17566, r_Bit_Index, 
            n17569, n35004, n18111, n25741, r_SM_Main, n35269, r_Rx_Data, 
            n35272, PIN_13_N_105, n35275, n35276, n35271, n35274, 
            n41248, n41247, n17576, n17575, n17574, n17573, n17572, 
            n17571, n17570, n17527, n17180, n17321, n4661, n35374, 
            n25555, n1, n24764, n4, n4_adj_1, n15912, n15917, 
            n4_adj_2, n6, n44844) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n35270;
    output [7:0]r_Clock_Count;
    input GND_net;
    input n35268;
    output n35273;
    input VCC_net;
    output rx_data_ready;
    input clk32MHz;
    input n18165;
    output [7:0]rx_data;
    input n35086;
    input n35088;
    input n35090;
    input n35000;
    input n34912;
    input n34804;
    input n34716;
    input n17566;
    output [2:0]r_Bit_Index;
    input n17569;
    input n35004;
    input n18111;
    input n25741;
    output [2:0]r_SM_Main;
    output n35269;
    output r_Rx_Data;
    output n35272;
    input PIN_13_N_105;
    output n35275;
    output n35276;
    output n35271;
    output n35274;
    output n41248;
    output n41247;
    input n17576;
    input n17575;
    input n17574;
    input n17573;
    input n17572;
    input n17571;
    input n17570;
    input n17527;
    output n17180;
    output n17321;
    output n4661;
    output n35374;
    output n25555;
    output n1;
    output n24764;
    output n4;
    output n4_adj_1;
    output n15912;
    output n15917;
    output n4_adj_2;
    output n6;
    output n44844;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n28525, n28524, n34812, n28523, r_Rx_Data_R, n28522, n28521, 
        n28520, n28519;
    wire [2:0]r_SM_Main_2__N_3249;
    
    wire n35368;
    wire [2:0]r_SM_Main_2__N_3255;
    
    wire n25413, n17094, n15738, n6_adj_3892;
    
    SB_LUT4 add_62_9_lut (.I0(n35268), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n28525), .O(n35270)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n35268), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n28524), .O(n35273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n34812));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18165));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n35086));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n35088));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n35090));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n35000));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n34912));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n34804));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n34716));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17566));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17569));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n35004));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18111));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n25741));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_8 (.CI(n28524), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n28525));
    SB_LUT4 add_62_7_lut (.I0(n35268), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n28523), .O(n35269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n28523), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n28524));
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 add_62_6_lut (.I0(n35268), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n28522), .O(n35272)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_CARRY add_62_6 (.CI(n28522), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n28523));
    SB_LUT4 add_62_5_lut (.I0(n35268), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n28521), .O(n35275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n28521), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n28522));
    SB_LUT4 add_62_4_lut (.I0(n35268), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n28520), .O(n35276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n28520), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n28521));
    SB_LUT4 add_62_3_lut (.I0(n35268), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n28519), .O(n35271)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n28519), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n28520));
    SB_LUT4 add_62_2_lut (.I0(n35268), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n35274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n28519));
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3249[2]), 
            .R(n35368));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i34870_2_lut (.I0(r_SM_Main_2__N_3249[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n41248));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34870_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34820_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3255[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n41247));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34820_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17576));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17575));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17574));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17573));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17572));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17571));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17570));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n17527));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n25413));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3249[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n17180));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i12576_3_lut (.I0(n17180), .I1(n25413), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17321));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12576_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1282_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4661));   // verilog/uart_rx.v(102[36:51])
    defparam i1282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n35374), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3249[2]));   // verilog/uart_rx.v(68[17:52])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n35374), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3255[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n25413), .I1(r_SM_Main_2__N_3249[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n25555));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i37346_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n35368));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i37346_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3249[2]), 
            .I3(r_SM_Main[0]), .O(n17094));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3255[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n17094), 
            .I3(rx_data_ready), .O(n34812));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i20043_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n24764));
    defparam i20043_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_140_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_140_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_142_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_142_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n15738), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n15912));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_3249[2]), .O(n15738));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_858 (.I0(r_Bit_Index[0]), .I1(n15738), .I2(GND_net), 
            .I3(GND_net), .O(n15917));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_858.LUT_INIT = 16'heeee;
    SB_LUT4 equal_145_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_145_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3255[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_adj_859 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3892));
    defparam i2_2_lut_adj_859.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(n6_adj_3892), 
            .I3(r_Clock_Count[4]), .O(n35374));
    defparam i1_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_rep_114_2_lut (.I0(r_Clock_Count[5]), .I1(n35374), .I2(GND_net), 
            .I3(GND_net), .O(n44844));
    defparam i1_rep_114_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n18067, encoder0_position, clk32MHz, 
            n18068, n18069, n18070, n18071, n18072, n18056, n18057, 
            n18058, n18059, n18060, n18061, n18062, n18063, n18064, 
            n18065, n18066, n18054, n18055, n18052, n18053, n18050, 
            n18051, data_o, n2998, GND_net, n17523, count_enable, 
            n18101, reg_B, n37457, PIN_2_c_0, n17526, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18067;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n18068;
    input n18069;
    input n18070;
    input n18071;
    input n18072;
    input n18056;
    input n18057;
    input n18058;
    input n18059;
    input n18060;
    input n18061;
    input n18062;
    input n18063;
    input n18064;
    input n18065;
    input n18066;
    input n18054;
    input n18055;
    input n18052;
    input n18053;
    input n18050;
    input n18051;
    output [1:0]data_o;
    output [23:0]n2998;
    input GND_net;
    input n17523;
    output count_enable;
    input n18101;
    output [1:0]reg_B;
    output n37457;
    input PIN_2_c_0;
    input n17526;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2994, n28596, n28595, n28594, n28593, 
        n28592, n28591, n28590, n28589, n28588, n28587, n28586, 
        n28585, n28584, n28583, n28582, n28581, n28580, n28579, 
        n28578, n28577, n28576, n28575, n28574, count_direction, 
        n28573;
    
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n18067));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n18068));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n18069));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n18070));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n18071));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n18072));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n18056));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n18057));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n18058));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n18059));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n18060));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n18061));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n18062));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n18063));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n18064));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n18065));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n18066));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n18054));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n18055));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n18052));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n18053));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n18050));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n18051));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_646_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2994), 
            .I3(n28596), .O(n2998[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_646_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2994), 
            .I3(n28595), .O(n2998[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_24 (.CI(n28595), .I0(encoder0_position[22]), .I1(n2994), 
            .CO(n28596));
    SB_LUT4 add_646_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2994), 
            .I3(n28594), .O(n2998[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_23 (.CI(n28594), .I0(encoder0_position[21]), .I1(n2994), 
            .CO(n28595));
    SB_LUT4 add_646_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2994), 
            .I3(n28593), .O(n2998[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_22 (.CI(n28593), .I0(encoder0_position[20]), .I1(n2994), 
            .CO(n28594));
    SB_LUT4 add_646_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2994), 
            .I3(n28592), .O(n2998[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_21 (.CI(n28592), .I0(encoder0_position[19]), .I1(n2994), 
            .CO(n28593));
    SB_LUT4 add_646_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2994), 
            .I3(n28591), .O(n2998[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_20 (.CI(n28591), .I0(encoder0_position[18]), .I1(n2994), 
            .CO(n28592));
    SB_LUT4 add_646_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2994), 
            .I3(n28590), .O(n2998[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_19 (.CI(n28590), .I0(encoder0_position[17]), .I1(n2994), 
            .CO(n28591));
    SB_LUT4 add_646_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2994), 
            .I3(n28589), .O(n2998[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_18 (.CI(n28589), .I0(encoder0_position[16]), .I1(n2994), 
            .CO(n28590));
    SB_LUT4 add_646_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2994), 
            .I3(n28588), .O(n2998[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_17 (.CI(n28588), .I0(encoder0_position[15]), .I1(n2994), 
            .CO(n28589));
    SB_LUT4 add_646_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2994), 
            .I3(n28587), .O(n2998[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_16 (.CI(n28587), .I0(encoder0_position[14]), .I1(n2994), 
            .CO(n28588));
    SB_LUT4 add_646_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2994), 
            .I3(n28586), .O(n2998[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_15 (.CI(n28586), .I0(encoder0_position[13]), .I1(n2994), 
            .CO(n28587));
    SB_LUT4 add_646_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2994), 
            .I3(n28585), .O(n2998[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_14 (.CI(n28585), .I0(encoder0_position[12]), .I1(n2994), 
            .CO(n28586));
    SB_LUT4 add_646_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2994), 
            .I3(n28584), .O(n2998[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_13 (.CI(n28584), .I0(encoder0_position[11]), .I1(n2994), 
            .CO(n28585));
    SB_LUT4 add_646_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2994), 
            .I3(n28583), .O(n2998[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_12 (.CI(n28583), .I0(encoder0_position[10]), .I1(n2994), 
            .CO(n28584));
    SB_LUT4 add_646_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2994), 
            .I3(n28582), .O(n2998[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_11 (.CI(n28582), .I0(encoder0_position[9]), .I1(n2994), 
            .CO(n28583));
    SB_LUT4 add_646_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2994), 
            .I3(n28581), .O(n2998[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_10 (.CI(n28581), .I0(encoder0_position[8]), .I1(n2994), 
            .CO(n28582));
    SB_LUT4 add_646_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2994), 
            .I3(n28580), .O(n2998[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_9 (.CI(n28580), .I0(encoder0_position[7]), .I1(n2994), 
            .CO(n28581));
    SB_LUT4 add_646_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2994), 
            .I3(n28579), .O(n2998[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_8 (.CI(n28579), .I0(encoder0_position[6]), .I1(n2994), 
            .CO(n28580));
    SB_LUT4 add_646_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2994), 
            .I3(n28578), .O(n2998[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_7 (.CI(n28578), .I0(encoder0_position[5]), .I1(n2994), 
            .CO(n28579));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17523));   // quad.v(35[10] 41[6])
    SB_LUT4 add_646_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2994), 
            .I3(n28577), .O(n2998[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_6 (.CI(n28577), .I0(encoder0_position[4]), .I1(n2994), 
            .CO(n28578));
    SB_LUT4 add_646_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2994), 
            .I3(n28576), .O(n2998[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_5 (.CI(n28576), .I0(encoder0_position[3]), .I1(n2994), 
            .CO(n28577));
    SB_LUT4 add_646_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2994), 
            .I3(n28575), .O(n2998[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_4 (.CI(n28575), .I0(encoder0_position[2]), .I1(n2994), 
            .CO(n28576));
    SB_LUT4 add_646_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2994), 
            .I3(n28574), .O(n2998[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_3 (.CI(n28574), .I0(encoder0_position[1]), .I1(n2994), 
            .CO(n28575));
    SB_LUT4 add_646_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n28573), .O(n2998[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_646_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_646_2 (.CI(n28573), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n28574));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_646_1 (.CI(GND_net), .I0(n2994), .I1(n2994), .CO(n28573));
    SB_LUT4 i923_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2994));   // quad.v(37[5] 40[8])
    defparam i923_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    \grp_debouncer(2,5)_U0  debounce (.n18101(n18101), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .GND_net(GND_net), .n37457(n37457), 
            .PIN_2_c_0(PIN_2_c_0), .n17526(n17526), .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18101, data_o, clk32MHz, reg_B, GND_net, 
            n37457, PIN_2_c_0, n17526, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18101;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n37457;
    input PIN_2_c_0;
    input n17526;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3559;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18101));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n37457), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i23421_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23421_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1203__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n37457));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1203__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1203__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17526));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i23430_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23430_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i23423_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23423_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n18075, encoder1_position, clk32MHz, 
            n18076, n18077, n18078, n18079, n18080, n18081, n18095, 
            n18096, n18097, n18093, n18094, n18091, n18092, n18089, 
            n18090, n18087, n18088, n18085, n18086, n18082, n18083, 
            n18084, n2948, GND_net, data_o, n17525, count_enable, 
            n18161, PIN_6_c_0, reg_B, PIN_7_c_1, n37455, n17539) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18075;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n18076;
    input n18077;
    input n18078;
    input n18079;
    input n18080;
    input n18081;
    input n18095;
    input n18096;
    input n18097;
    input n18093;
    input n18094;
    input n18091;
    input n18092;
    input n18089;
    input n18090;
    input n18087;
    input n18088;
    input n18085;
    input n18086;
    input n18082;
    input n18083;
    input n18084;
    output [23:0]n2948;
    input GND_net;
    output [1:0]data_o;
    input n17525;
    output count_enable;
    input n18161;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    output n37455;
    input n17539;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n2935, n28630, B_delayed, n28629, A_delayed, count_direction, 
        n28628, n28627, n28626, n28625, n28624, n28623, n28622, 
        n28621, n28620, n28619, n28618, n28617, n28616, n28615, 
        n28614, n28613, n28612, n28611, n28610, n28609, n28608, 
        n28607;
    
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n18075));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n18076));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n18077));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n18078));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n18079));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n18080));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n18081));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18095));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18096));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18097));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18093));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18094));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18091));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18092));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18089));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18090));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18087));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18088));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18085));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18086));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n18082));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n18083));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n18084));   // quad.v(35[10] 41[6])
    SB_LUT4 add_620_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2935), 
            .I3(n28630), .O(n2948[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_LUT4 add_620_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2935), 
            .I3(n28629), .O(n2948[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_620_24 (.CI(n28629), .I0(encoder1_position[22]), .I1(n2935), 
            .CO(n28630));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_620_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2935), 
            .I3(n28628), .O(n2948[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_23 (.CI(n28628), .I0(encoder1_position[21]), .I1(n2935), 
            .CO(n28629));
    SB_LUT4 add_620_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2935), 
            .I3(n28627), .O(n2948[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_22 (.CI(n28627), .I0(encoder1_position[20]), .I1(n2935), 
            .CO(n28628));
    SB_LUT4 add_620_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2935), 
            .I3(n28626), .O(n2948[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_21 (.CI(n28626), .I0(encoder1_position[19]), .I1(n2935), 
            .CO(n28627));
    SB_LUT4 add_620_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2935), 
            .I3(n28625), .O(n2948[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_20 (.CI(n28625), .I0(encoder1_position[18]), .I1(n2935), 
            .CO(n28626));
    SB_LUT4 add_620_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2935), 
            .I3(n28624), .O(n2948[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_19 (.CI(n28624), .I0(encoder1_position[17]), .I1(n2935), 
            .CO(n28625));
    SB_LUT4 add_620_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2935), 
            .I3(n28623), .O(n2948[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_18 (.CI(n28623), .I0(encoder1_position[16]), .I1(n2935), 
            .CO(n28624));
    SB_LUT4 add_620_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2935), 
            .I3(n28622), .O(n2948[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_17 (.CI(n28622), .I0(encoder1_position[15]), .I1(n2935), 
            .CO(n28623));
    SB_LUT4 add_620_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2935), 
            .I3(n28621), .O(n2948[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_16 (.CI(n28621), .I0(encoder1_position[14]), .I1(n2935), 
            .CO(n28622));
    SB_LUT4 add_620_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2935), 
            .I3(n28620), .O(n2948[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_15 (.CI(n28620), .I0(encoder1_position[13]), .I1(n2935), 
            .CO(n28621));
    SB_LUT4 add_620_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2935), 
            .I3(n28619), .O(n2948[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_14 (.CI(n28619), .I0(encoder1_position[12]), .I1(n2935), 
            .CO(n28620));
    SB_LUT4 add_620_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2935), 
            .I3(n28618), .O(n2948[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_13 (.CI(n28618), .I0(encoder1_position[11]), .I1(n2935), 
            .CO(n28619));
    SB_LUT4 add_620_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2935), 
            .I3(n28617), .O(n2948[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_12 (.CI(n28617), .I0(encoder1_position[10]), .I1(n2935), 
            .CO(n28618));
    SB_LUT4 add_620_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2935), 
            .I3(n28616), .O(n2948[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_11 (.CI(n28616), .I0(encoder1_position[9]), .I1(n2935), 
            .CO(n28617));
    SB_LUT4 add_620_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2935), 
            .I3(n28615), .O(n2948[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_10 (.CI(n28615), .I0(encoder1_position[8]), .I1(n2935), 
            .CO(n28616));
    SB_LUT4 add_620_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2935), 
            .I3(n28614), .O(n2948[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_9 (.CI(n28614), .I0(encoder1_position[7]), .I1(n2935), 
            .CO(n28615));
    SB_LUT4 add_620_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2935), 
            .I3(n28613), .O(n2948[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_8 (.CI(n28613), .I0(encoder1_position[6]), .I1(n2935), 
            .CO(n28614));
    SB_LUT4 add_620_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2935), 
            .I3(n28612), .O(n2948[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_7 (.CI(n28612), .I0(encoder1_position[5]), .I1(n2935), 
            .CO(n28613));
    SB_LUT4 add_620_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2935), 
            .I3(n28611), .O(n2948[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_6 (.CI(n28611), .I0(encoder1_position[4]), .I1(n2935), 
            .CO(n28612));
    SB_LUT4 add_620_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2935), 
            .I3(n28610), .O(n2948[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_5 (.CI(n28610), .I0(encoder1_position[3]), .I1(n2935), 
            .CO(n28611));
    SB_LUT4 add_620_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2935), 
            .I3(n28609), .O(n2948[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_4 (.CI(n28609), .I0(encoder1_position[2]), .I1(n2935), 
            .CO(n28610));
    SB_LUT4 add_620_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2935), 
            .I3(n28608), .O(n2948[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_3 (.CI(n28608), .I0(encoder1_position[1]), .I1(n2935), 
            .CO(n28609));
    SB_LUT4 add_620_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n28607), .O(n2948[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_620_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_620_2 (.CI(n28607), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n28608));
    SB_CARRY add_620_1 (.CI(GND_net), .I0(n2935), .I1(n2935), .CO(n28607));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17525));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i933_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2935));   // quad.v(37[5] 40[8])
    defparam i933_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n18161(n18161), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B}), .PIN_7_c_1(PIN_7_c_1), 
            .GND_net(GND_net), .n37455(n37455), .n17539(n17539)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n18161, data_o, clk32MHz, PIN_6_c_0, reg_B, 
            PIN_7_c_1, GND_net, n37455, n17539) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18161;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    input GND_net;
    output n37455;
    input n17539;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3559;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18161));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_6_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_7_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n37455), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i23443_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23443_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1204__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1204__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1204__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17539));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i23452_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23452_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i23445_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23445_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n37455));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (GND_net, VCC_net, PIN_19_c_0, 
            CLK_c, \half_duty_new[0] , n18136, \half_duty[0][6] , n18137, 
            \half_duty[0][7] , n18134, \half_duty[0][4] , n18135, \half_duty[0][5] , 
            n18132, \half_duty[0][2] , n18133, \half_duty[0][3] , n18131, 
            \half_duty[0][1] , n1144, \half_duty[0][0] , \half_duty_new[1] , 
            \half_duty_new[2] , \half_duty_new[3] , \half_duty_new[4] , 
            \half_duty_new[5] , \half_duty_new[6] , \half_duty_new[7] , 
            pwm_setpoint, n17531) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input GND_net;
    input VCC_net;
    output PIN_19_c_0;
    input CLK_c;
    output \half_duty_new[0] ;
    input n18136;
    output \half_duty[0][6] ;
    input n18137;
    output \half_duty[0][7] ;
    input n18134;
    output \half_duty[0][4] ;
    input n18135;
    output \half_duty[0][5] ;
    input n18132;
    output \half_duty[0][2] ;
    input n18133;
    output \half_duty[0][3] ;
    input n18131;
    output \half_duty[0][1] ;
    output n1144;
    output \half_duty[0][0] ;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[5] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input [22:0]pwm_setpoint;
    input n17531;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n29243;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n29244;
    wire [10:0]n49;
    
    wire pwm_out_0__N_582, n17118;
    wire [9:0]half_duty_new_9__N_664;
    
    wire pause_counter_0, n36266, pause_counter_0__N_612;
    wire [10:0]pwm_out_0__N_587;
    
    wire n8, n9, n39091, n2, n5, n4, n7, n39103, n6, n22, 
        n10, n3, n1, pwm_out_0__N_586, n21, n13, n12, n18, n16, 
        n17, n15, n28468, n28467, n28466, n28465, n28464, n28463, 
        n28462, n28461, n28460, n28459, n28458;
    wire [22:0]n5612;
    
    wire n28856, n28855, n28854, n28853, n28852, n28851, n28850, 
        n28849, n28848, n28847, n28846, n28845, n20, n28844, n28843, 
        n28842, n28841, n28840, n28839, n28838, n28837, n28836, 
        n28835, n19, n6_adj_3889, n28834, n28833, n28832, n28831, 
        n28830, n28829, n28828, n28827, n28826, n28825, n28824, 
        n28823, n28822, n28821, n28820, n28819, n28818, n28817, 
        n28816, n28815, n28814, n29252, n29251, n29250, n29249, 
        n29248, n29247, n29246, n29245;
    
    SB_CARRY count_0__1201_add_4_3 (.CI(n29243), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n29244));
    SB_LUT4 count_0__1201_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n29243));
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n17118), .D(pwm_out_0__N_582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_664[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n18136));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n18137));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n18134));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0][5] ), .C(CLK_c), .D(n18135));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n18132));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n18133));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n18131));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i37360_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_582), .I2(GND_net), 
            .I3(GND_net), .O(n36266));
    defparam i37360_2_lut.LUT_INIT = 16'h1111;
    SB_DFFESR count_0__1201__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[10]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[9]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[8]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[7]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[6]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[5]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[4]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1201__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[3]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n36266));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0][5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i7_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[6]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR count_0__1201__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[2]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32310_2_lut (.I0(n8), .I1(n9), .I2(GND_net), .I3(GND_net), 
            .O(n39091));
    defparam i32310_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32322_4_lut (.I0(n2), .I1(n5), .I2(n4), .I3(n7), .O(n39103));
    defparam i32322_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(\count[0] [10]), .I1(n39103), .I2(n39091), 
            .I3(n6), .O(n22));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i9_4_lut (.I0(n10), .I1(n3), .I2(n1), .I3(pwm_out_0__N_586), 
            .O(n21));
    defparam i9_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut (.I0(n21), .I1(pause_counter_0), .I2(pwm_out_0__N_582), 
            .I3(n22), .O(n17118));
    defparam i1_4_lut.LUT_INIT = 16'h2303;
    SB_LUT4 i2_4_lut (.I0(\half_duty[0][1] ), .I1(\half_duty[0][6] ), .I2(\count[0] [1]), 
            .I3(\count[0] [6]), .O(n13));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_855 (.I0(\half_duty[0][5] ), .I1(\half_duty[0][4] ), 
            .I2(\count[0] [5]), .I3(\count[0] [4]), .O(n12));   // vhdl/pwm.vhd(80[8:31])
    defparam i1_4_lut_adj_855.LUT_INIT = 16'h7bde;
    SB_DFFESR count_0__1201__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[1]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i7_3_lut (.I0(n13), .I1(\count[0] [8]), .I2(\count[0] [9]), 
            .I3(GND_net), .O(n18));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(\count[0] [10]), .I1(\half_duty[0][0] ), .I2(\count[0] [0]), 
            .I3(GND_net), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i6_3_lut (.I0(\half_duty[0][2] ), .I1(n12), .I2(\count[0] [2]), 
            .I3(GND_net), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i4_4_lut (.I0(\half_duty[0][3] ), .I1(\half_duty[0][7] ), .I2(\count[0] [3]), 
            .I3(\count[0] [7]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10_4_lut_adj_856 (.I0(n15), .I1(n17), .I2(n16), .I3(n18), 
            .O(pwm_out_0__N_582));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_856.LUT_INIT = 16'hfffe;
    SB_DFFESR count_0__1201__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[0]), .R(n1144));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_612));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY pwm_out_0__I_20_13 (.CI(n28468), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_586));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n28467), .I0(VCC_net), .I1(VCC_net), 
            .CO(n28468));
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_664[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_664[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_664[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_664[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(\half_duty_new[5] ), .C(CLK_c), .D(half_duty_new_9__N_664[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_664[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_664[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n28466), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n28466), .I0(VCC_net), .I1(VCC_net), 
            .CO(n28467));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n28465), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_10 (.CI(n28465), .I0(GND_net), .I1(VCC_net), 
            .CO(n28466));
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_587[7]), 
            .I3(n28464), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n28464), .I0(GND_net), .I1(pwm_out_0__N_587[7]), 
            .CO(n28465));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_587[6]), 
            .I3(n28463), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n28463), .I0(VCC_net), .I1(pwm_out_0__N_587[6]), 
            .CO(n28464));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_587[5]), 
            .I3(n28462), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n28462), .I0(GND_net), .I1(pwm_out_0__N_587[5]), 
            .CO(n28463));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_587[4]), 
            .I3(n28461), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n28461), .I0(GND_net), .I1(pwm_out_0__N_587[4]), 
            .CO(n28462));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_587[3]), 
            .I3(n28460), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n28460), .I0(GND_net), .I1(pwm_out_0__N_587[3]), 
            .CO(n28461));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_587[2]), 
            .I3(n28459), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n28459), .I0(GND_net), .I1(pwm_out_0__N_587[2]), 
            .CO(n28460));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_587[1]), 
            .I3(n28458), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_3 (.CI(n28458), .I0(GND_net), .I1(pwm_out_0__N_587[1]), 
            .CO(n28459));
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_587[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_587[0]), 
            .CO(n28458));
    SB_LUT4 add_2052_24_lut (.I0(GND_net), .I1(n5612[22]), .I2(pwm_setpoint[22]), 
            .I3(n28856), .O(half_duty_new_9__N_664[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2052_23_lut (.I0(GND_net), .I1(n5612[21]), .I2(pwm_setpoint[21]), 
            .I3(n28855), .O(half_duty_new_9__N_664[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_23 (.CI(n28855), .I0(n5612[21]), .I1(pwm_setpoint[21]), 
            .CO(n28856));
    SB_LUT4 add_2052_22_lut (.I0(GND_net), .I1(n5612[20]), .I2(pwm_setpoint[20]), 
            .I3(n28854), .O(half_duty_new_9__N_664[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_22 (.CI(n28854), .I0(n5612[20]), .I1(pwm_setpoint[20]), 
            .CO(n28855));
    SB_LUT4 add_2052_21_lut (.I0(GND_net), .I1(n5612[19]), .I2(pwm_setpoint[19]), 
            .I3(n28853), .O(half_duty_new_9__N_664[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_21 (.CI(n28853), .I0(n5612[19]), .I1(pwm_setpoint[19]), 
            .CO(n28854));
    SB_LUT4 add_2052_20_lut (.I0(GND_net), .I1(n5612[18]), .I2(pwm_setpoint[18]), 
            .I3(n28852), .O(half_duty_new_9__N_664[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_20 (.CI(n28852), .I0(n5612[18]), .I1(pwm_setpoint[18]), 
            .CO(n28853));
    SB_LUT4 add_2052_19_lut (.I0(GND_net), .I1(n5612[17]), .I2(pwm_setpoint[17]), 
            .I3(n28851), .O(half_duty_new_9__N_664[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_19 (.CI(n28851), .I0(n5612[17]), .I1(pwm_setpoint[17]), 
            .CO(n28852));
    SB_LUT4 add_2052_18_lut (.I0(GND_net), .I1(n5612[16]), .I2(pwm_setpoint[16]), 
            .I3(n28850), .O(half_duty_new_9__N_664[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_18 (.CI(n28850), .I0(n5612[16]), .I1(pwm_setpoint[16]), 
            .CO(n28851));
    SB_LUT4 add_2052_17_lut (.I0(GND_net), .I1(n5612[15]), .I2(pwm_setpoint[15]), 
            .I3(n28849), .O(half_duty_new_9__N_664[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2052_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2052_17 (.CI(n28849), .I0(n5612[15]), .I1(pwm_setpoint[15]), 
            .CO(n28850));
    SB_CARRY add_2052_16 (.CI(n28848), .I0(n5612[14]), .I1(pwm_setpoint[14]), 
            .CO(n28849));
    SB_CARRY add_2052_15 (.CI(n28847), .I0(n5612[13]), .I1(pwm_setpoint[13]), 
            .CO(n28848));
    SB_CARRY add_2052_14 (.CI(n28846), .I0(n5612[12]), .I1(pwm_setpoint[12]), 
            .CO(n28847));
    SB_CARRY add_2052_13 (.CI(n28845), .I0(n5612[11]), .I1(pwm_setpoint[11]), 
            .CO(n28846));
    SB_LUT4 i8_4_lut (.I0(\count[0] [6]), .I1(\count[0] [0]), .I2(\count[0] [10]), 
            .I3(\count[0] [1]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hbfff;
    SB_CARRY add_2052_12 (.CI(n28844), .I0(n5612[10]), .I1(pwm_setpoint[10]), 
            .CO(n28845));
    SB_CARRY add_2052_11 (.CI(n28843), .I0(n5612[9]), .I1(pwm_setpoint[9]), 
            .CO(n28844));
    SB_CARRY add_2052_10 (.CI(n28842), .I0(n5612[8]), .I1(pwm_setpoint[8]), 
            .CO(n28843));
    SB_CARRY add_2052_9 (.CI(n28841), .I0(n5612[7]), .I1(pwm_setpoint[7]), 
            .CO(n28842));
    SB_CARRY add_2052_8 (.CI(n28840), .I0(n5612[6]), .I1(pwm_setpoint[6]), 
            .CO(n28841));
    SB_CARRY add_2052_7 (.CI(n28839), .I0(n5612[5]), .I1(pwm_setpoint[5]), 
            .CO(n28840));
    SB_CARRY add_2052_6 (.CI(n28838), .I0(n5612[4]), .I1(pwm_setpoint[4]), 
            .CO(n28839));
    SB_CARRY add_2052_5 (.CI(n28837), .I0(n5612[3]), .I1(pwm_setpoint[3]), 
            .CO(n28838));
    SB_CARRY add_2052_4 (.CI(n28836), .I0(n5612[2]), .I1(pwm_setpoint[2]), 
            .CO(n28837));
    SB_CARRY add_2052_3 (.CI(n28835), .I0(n5612[1]), .I1(pwm_setpoint[1]), 
            .CO(n28836));
    SB_LUT4 i7_4_lut (.I0(pause_counter_0), .I1(\count[0] [9]), .I2(\count[0] [8]), 
            .I3(\count[0] [7]), .O(n19));
    defparam i7_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut (.I0(\count[0] [4]), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n6_adj_3889));
    defparam i1_3_lut.LUT_INIT = 16'h0202;
    SB_CARRY add_2052_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n28835));
    SB_LUT4 add_2060_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n28834), .O(n5612[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2060_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n28833), .O(n5612[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_22 (.CI(n28833), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n28834));
    SB_LUT4 add_2060_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n28832), .O(n5612[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_21 (.CI(n28832), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n28833));
    SB_LUT4 add_2060_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n28831), .O(n5612[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_20 (.CI(n28831), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n28832));
    SB_LUT4 add_2060_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n28830), .O(n5612[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_19 (.CI(n28830), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n28831));
    SB_LUT4 add_2060_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n28829), .O(n5612[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_18 (.CI(n28829), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n28830));
    SB_LUT4 add_2060_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n28828), .O(n5612[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_17 (.CI(n28828), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n28829));
    SB_LUT4 add_2060_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n28827), .O(n5612[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_16 (.CI(n28827), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n28828));
    SB_LUT4 add_2060_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n28826), .O(n5612[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_15 (.CI(n28826), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n28827));
    SB_LUT4 add_2060_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n28825), .O(n5612[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_14 (.CI(n28825), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n28826));
    SB_LUT4 add_2060_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n28824), .O(n5612[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_13 (.CI(n28824), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n28825));
    SB_LUT4 add_2060_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n28823), .O(n5612[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_12 (.CI(n28823), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n28824));
    SB_LUT4 add_2060_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n28822), .O(n5612[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_11 (.CI(n28822), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n28823));
    SB_LUT4 add_2060_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n28821), .O(n5612[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_10 (.CI(n28821), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n28822));
    SB_LUT4 add_2060_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n28820), .O(n5612[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_9 (.CI(n28820), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n28821));
    SB_LUT4 add_2060_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n28819), .O(n5612[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_8 (.CI(n28819), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n28820));
    SB_LUT4 add_2060_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n28818), .O(n5612[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_7 (.CI(n28818), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n28819));
    SB_LUT4 add_2060_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n28817), .O(n5612[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_6 (.CI(n28817), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n28818));
    SB_LUT4 add_2060_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n28816), .O(n5612[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_5 (.CI(n28816), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n28817));
    SB_LUT4 add_2060_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n28815), .O(n5612[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_4 (.CI(n28815), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n28816));
    SB_LUT4 i4_4_lut_adj_857 (.I0(\count[0] [5]), .I1(\count[0] [2]), .I2(\count[0] [3]), 
            .I3(n6_adj_3889), .O(n1144));
    defparam i4_4_lut_adj_857.LUT_INIT = 16'h8000;
    SB_LUT4 add_2060_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n28814), .O(n5612[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_3 (.CI(n28814), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n28815));
    SB_LUT4 add_2060_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5612[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2060_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2060_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n28814));
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n17531));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 count_0__1201_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n29252), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1201_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n29251), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_11 (.CI(n29251), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n29252));
    SB_LUT4 count_0__1201_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n29250), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_10 (.CI(n29250), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n29251));
    SB_LUT4 count_0__1201_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n29249), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_9 (.CI(n29249), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n29250));
    SB_LUT4 count_0__1201_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n29248), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_8 (.CI(n29248), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n29249));
    SB_LUT4 count_0__1201_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n29247), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_7 (.CI(n29247), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n29248));
    SB_LUT4 count_0__1201_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n29246), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_6 (.CI(n29246), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n29247));
    SB_LUT4 count_0__1201_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n29245), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_5 (.CI(n29245), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n29246));
    SB_LUT4 count_0__1201_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n29244), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1201_add_4_4 (.CI(n29244), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n29245));
    SB_LUT4 count_0__1201_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n29243), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1201_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, IntegralLimit, \Ki[1] , \Ki[0] , \Ki[2] , 
            \Ki[3] , \Kp[1] , \Kp[0] , \Ki[4] , \Ki[5] , \Kp[2] , 
            \Kp[3] , \Ki[6] , \Kp[4] , \Ki[7] , \Kp[5] , \Kp[6] , 
            \Kp[7] , duty, PWMLimit, clk32MHz, VCC_net, n44224, 
            motor_state, n25, setpoint) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input [23:0]IntegralLimit;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Ki[6] ;
    input \Kp[4] ;
    input \Ki[7] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    output [23:0]duty;
    input [23:0]PWMLimit;
    input clk32MHz;
    input VCC_net;
    output n44224;
    input [23:0]motor_state;
    input n25;
    input [23:0]setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n30423;
    wire [10:0]n8304;
    
    wire n30424;
    wire [11:0]n8290;
    
    wire n30422;
    wire [23:0]n257;
    
    wire n13, n10;
    wire [23:0]n1;
    
    wire n12, n35, n30, n30421, n545, n30420;
    wire [8:0]n8032;
    wire [7:0]n8043;
    
    wire n554, n30207;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    
    wire n98, n30208, n29, n481, n30206, n472, n30419, n11, 
        n9, n41613, n42341, n408, n30205;
    wire [23:0]duty_23__N_3478;
    wire [23:0]n3054;
    wire [23:0]n3079;
    
    wire n28571, n28572, n19, n17, n15, n42299, n25_c, n23_adj_3561, 
        n21, n43203, n31, n29_adj_3562, n27, n42708, n399, n30418, 
        n335, n30204, n28570, n39, n28702, n326, n30417, n262, 
        n30203, n28703, n37, n28701, n28569, n171, n189, n30202, 
        n253, n30416, n47, n116, n180, n30415;
    wire [9:0]n8020;
    
    wire n30201, n38, n107, n30200;
    wire [12:0]n8275;
    
    wire n30414, n30199, n30413, n244;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n107_adj_3564, n38_adj_3565, n317, n35_adj_3566, n28700, 
        n33, n28699, n30412, n31_adj_3568, n28698, n390, n180_adj_3570, 
        n253_adj_3571, n37_adj_3572, n33_adj_3573, n43347, n463, n326_adj_3574, 
        n536, n399_adj_3576, n472_adj_3577, n545_adj_3578, n43, n16;
    wire [47:0]n155;
    
    wire n256, n6_adj_3580, n42758, n42759, n101, n32, n110, n41, 
        n174, n183, n317_adj_3582, n390_adj_3583, n463_adj_3584, n247, 
        n30411, n30410, n308, n256_adj_3585, n320, n393, n329, 
        n402, n466, n539, n551, n30198, n165, n475, n548, n30409, 
        n113, n536_adj_3588, n28568, n44, n186_adj_3589, n381, n454, 
        n104, n527, n35_adj_3590, n177, n8_adj_3591, n29_adj_3592, 
        n28697, n45, n24, n542, n30408, n478, n30197, n41563, 
        n41463, n469, n30407, n27_adj_3594, n28696;
    wire [23:0]duty_23__N_3355;
    wire [23:0]\PID_CONTROLLER.err_23__N_3379 ;
    
    wire n28567, n259_adj_3596, n405, n30196, n396, n30406, n250, 
        n332, n30195, n323, n30405, n30404, n30194, n30403, n92, 
        n23_adj_3597, n30193;
    wire [13:0]n8259;
    
    wire n30402, n30401;
    wire [10:0]n8007;
    
    wire n30192, n165_adj_3598, n238, n25_adj_3599, n28695, n30191, 
        n311, n101_adj_3600, n41_adj_3601, n39_adj_3602, n30400, n32_adj_3603, 
        n30399, n30190, n30398, n45_adj_3604, n43_adj_3605, n30189, 
        n23_adj_3606, n28694, n37_adj_3607, n30397, n30188, n21_adj_3608, 
        n28693, n29_adj_3609, n30396, n30187, n28566, n30395, n31_adj_3610, 
        n384, n30394, n30186, n30185, n30393, n23_adj_3611, n25_adj_3612, 
        n41453, n42936, n30392, n174_adj_3613, n30184, n30391, n28565, 
        n30183, n42202, n41179, n4, n42754, n35_adj_3614, n33_adj_3615, 
        n11_adj_3616, n13_adj_3617, n15_adj_3618, n457, n530, n27_adj_3619, 
        n9_adj_3620, n30390, n42755, n41534, n41522, n41519, n43373, 
        n42204, n43456, n43457, n39_adj_3622, n43433, n41_adj_3623, 
        n41468, n17_adj_3624, n19_adj_3625, n21_adj_3626, n41741, 
        n41720;
    wire [11:0]n7993;
    
    wire n30182, n43183, n40, n19_adj_3627, n28692, n28564;
    wire [14:0]n8242;
    
    wire n30389, n30388, n30387, n30181, n17_adj_3628, n28691, n30180, 
        n30386, n30179, n30385, n30178, n30177, n43185, n47_adj_3629, 
        n12_adj_3630, n30_adj_3631, n30384, n30383, n41789, n42437, 
        n42427, n43248, n15_adj_3632, n28690, n42784, n43360, n30176, 
        n30382, n30175, n13_adj_3633, n28689, n30381, n30174, n30380, 
        n30173, n6_adj_3634, n43047, n43048, n30172, n11_adj_3635, 
        n28688, n30379, n16_adj_3636, n24_adj_3637, n41623, n8_adj_3638, 
        n41619, n42932, n42192, n30378, n4_adj_3639, n43045, n43046, 
        n30377, n238_adj_3640, n448, n9_adj_3641, n28687, n311_adj_3642, 
        n521, n41696, n384_adj_3643, n30376, n10_adj_3644, n41692, 
        n43288, n247_adj_3645;
    wire [12:0]n7978;
    
    wire n30171, n30170, n42194, n43426, n43427, n43415, n7_adj_3646, 
        n28686, n41625, n30169, n43343, n42200, n43345, n5, n28685;
    wire [15:0]n8224;
    
    wire n30375, n30374, duty_23__N_3502, n3, n28684, n28563, n457_adj_3648, 
        n30373, n28562, n530_adj_3649, n30168, n30167, n30372, n30166, 
        n30371;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3454 ;
    
    wire n320_adj_3651, n30370, n542_adj_3652, n30165, n469_adj_3653, 
        n30164, n396_adj_3654, n30163, n30369, n323_adj_3655, n30162, 
        n30368, n28561, n30367, n533, n30366, n250_adj_3656, n30161, 
        n177_adj_3657, n30160, n35_adj_3658, n104_adj_3659, n460, 
        n30365, n28560, n387, n30364, n95, n26;
    wire [13:0]n7962;
    
    wire n30159, n168, n314, n30363, n241, n241_adj_3660, n30362, 
        n314_adj_3661, n30158, n86, n17_adj_3662, n387_adj_3663, n168_adj_3664, 
        n30361, n30157, n28559, n26_adj_3665, n95_adj_3666, n30156;
    wire [16:0]n8205;
    
    wire n30360, n30155, n30359, n30358, n30154, n28558, n30357;
    wire [21:0]n7798;
    wire [20:0]n7822;
    
    wire n29693, n30153, n29692, n539_adj_3667, n30152, n30356, 
        n466_adj_3668, n30151, n29691, n29690, n393_adj_3669, n29689, 
        n30355, n30150, n30354, n30353, n29688, n460_adj_3670, n30149, 
        n159, n29687, n29686, n30352, n533_adj_3671, n28557, n30148, 
        n30351, n29685, n30350, n30349, n30147, n29684, n30348, 
        n30347;
    wire [14:0]n7945;
    
    wire n30146, n30346, n30145, n30144, n232, n29683, n30345;
    wire [17:0]n8185;
    
    wire n30344, n30343, n30342, n30341, n30143, n30340, n30339, 
        n30338, n30142, n30337, n29682, n30141, n30336, n30335, 
        n28556, n30334, n30140, n30139, n29681, n30333, n30332, 
        n30331, n30138, n30330, n28555, n29680, n30137, n29679, 
        n30136, n30135, n305, n515, n29678, n235, n30329, n442, 
        n29677, n369, n29676, n244_adj_3672, n30134, n296, n29675, 
        n162, n30328, n20_adj_3673, n89;
    wire [18:0]n8164;
    
    wire n30327, n30326, n30325, n171_adj_3674, n30133, n223, n29674, 
        n30324, n29_adj_3675, n98_adj_3676, n150, n29673, n28554, 
        n378, n8_adj_3677, n77, n30323;
    wire [15:0]n7927;
    
    wire n30132, n30131, n30130, n30322, n28553, n30321, n30129, 
        n451, n524, n30320, n30128, n30319, n30318, n17_adj_3678, 
        n9_adj_3679, n28552, n30317, n11_adj_3680, n41395, n41385, 
        n45150, n42651, n42635, n45132, n42633, n42625, n30316, 
        n45126, n30127, n30126, n41854, n41868, n43_adj_3681, n16_adj_3682;
    wire [23:0]n28;
    
    wire \PID_CONTROLLER.integral_23__N_3451 , n41800, n8_adj_3683, n45_adj_3684, 
        n24_adj_3685, n41889, n30315, n42529, n42521, n43264, n42832, 
        n43368, n42055, n45119, n30314, n42603, n45114, n12_adj_3686, 
        n41948, n45137, n30125, n10_adj_3687, n30_adj_3688, n43113, 
        n30124, n41982, n45117, n42880, n45143, n43276, n45108, 
        n43446, n45105, n16_adj_3689, n30313, n41895, n24_adj_3690, 
        n6_adj_3691, n43065, n43066, n41899, n8_adj_3692, n45103, 
        n42928, n42172, n4_adj_3693, n43053, n43054, n12_adj_3694, 
        n41830, n10_adj_3695, n30_adj_3696, n41834, n43286, n42184, 
        n43424, n43425, n43417, n6_adj_3697, n43055, n43056, n41808, 
        n42930, n42182, n28551, n30312, n41_adj_3698, n41812, n43339, 
        n42190, n43341, n4_adj_3699, n43061, n43062, n41964, n43284, 
        n42174, n30311, n43422, n43423, n43419, n41901, n43335, 
        n42180, \PID_CONTROLLER.integral_23__N_3453 , n30123, n43337, 
        n30310, n30122, n30121, n30120;
    wire [19:0]n8142;
    
    wire n30309, n30308, n30119, n30118, n30307, n30306, n28550;
    wire [16:0]n7908;
    
    wire n30117, n30116, n30305, n30304, n30115, n30303, n30114, 
        n30113, n30302, n30112, n30111, n30301, n30110, n30300, 
        n30109, n30108, n30299, n30107, n30298, n30106, n30297, 
        n30105, n30296, n30104, n30295, n30103, n30102, n23_adj_3701, 
        n92_adj_3702, n375, n30294;
    wire [17:0]n7888;
    
    wire n30101, n302, n30293, n30100, n229, n30292, n30099, n156, 
        n30291, n30098, n14_adj_3703, n83, n30097;
    wire [20:0]n8119;
    
    wire n30290, n30096, n30289, n30095, n30094, n30093, n30288, 
        n30092, n30287, n30091, n30286, n527_adj_3704, n30090, n30285, 
        n454_adj_3705, n30089, n381_adj_3706, n30088, n30284, n308_adj_3707, 
        n30087, n30283, n235_adj_3708, n30086, n30282, n162_adj_3709, 
        n30085;
    wire [5:0]n8359;
    
    wire n31074, n490, n30470, n30281, n20_adj_3710, n89_adj_3711;
    wire [4:0]n8367;
    
    wire n417, n30469, n30280;
    wire [18:0]n7867;
    
    wire n30084, n30083, n30279, n30082, n344, n30468, n30278, 
        n30081, n30277, n30080, n271_adj_3712, n30467, n30079, n198, 
        n30466, n56, n125_adj_3713, n518, n30276, n30078;
    wire [6:0]n8350;
    
    wire n560, n30465, n445, n30275, n30077, n30076, n372, n30274, 
        n487, n30464, n30075, n299, n30273, n30074, n226, n30272, 
        n414, n30463, n30073, n153, n30271, n524_adj_3714, n30072, 
        n451_adj_3715, n30071, n341, n30462, n11_adj_3716, n80, 
        n378_adj_3717, n30070, n305_adj_3718, n30069, n41237;
    wire [21:0]n8095;
    
    wire n30270, n30269, n232_adj_3719, n30068, n268_adj_3720, n30461, 
        n159_adj_3721, n30067, n17_adj_3722, n86_adj_3723, n30268;
    wire [19:0]n7845;
    
    wire n30066, n195_adj_3724, n30460, n30267, n53, n122, n30065, 
        n30064, n30063;
    wire [7:0]n8340;
    
    wire n30459, n557, n30458, n30062, n30266, n30061, n30265, 
        n30060, n30059, n484, n30457, n30264, n411, n30456, n30263, 
        n30058, n30057, n30262, n338, n30455, n30056, n30261, 
        n30055, n30260, n30054, n265_adj_3726, n30454, n30259, n521_adj_3727, 
        n30053, n30258, n448_adj_3728, n30052, n192_adj_3729, n30453, 
        n30257, n375_adj_3730, n30051, n30256, n302_adj_3731, n30050, 
        n50, n119, n229_adj_3732, n30049, n30255, n156_adj_3733, 
        n30048, n512, n30254, n14_adj_3734, n83_adj_3735;
    wire [8:0]n8329;
    
    wire n30452, n30047, n439, n30253, n30046, n30045, n30451, 
        n366, n30252, n30044, n293, n30251, n554_adj_3744, n30450, 
        n30043, n481_adj_3745, n30449, n220, n30250, n30042, n30041, 
        n147, n30249, n30040, n5_adj_3746, n74, n408_adj_3747, n30448, 
        n335_adj_3748, n30447, n30039, n30248, n30038, n30247, n30037, 
        n262_adj_3749, n30446, n30246, n189_adj_3750, n30445, n29303, 
        n30036, n30245, n29302, n30035, n47_adj_3751, n116_adj_3752, 
        n30244, n29301, n30034, n29300, n30243, n30242, n518_adj_3753, 
        n30033;
    wire [9:0]n8317;
    
    wire n30444, n29299, n30241, n445_adj_3754, n30032, n29298, 
        n30443, n372_adj_3755, n30031, n29297, n30240, n29296, n30442, 
        n30239, n299_adj_3756, n30030, n226_adj_3757, n30029, n29295, 
        n29294, n30238, n29293, n30237, n153_adj_3758, n30028, n551_adj_3759, 
        n30441, n29292, n30236, n11_adj_3760, n80_adj_3761, n29291;
    wire [0:0]n6244;
    
    wire n30027, n30235, n30026, n25020, n478_adj_3762, n30440, 
        n29290, n30025, n29289, n30234, n30024, n29288, n515_adj_3763, 
        n30233, n30023, n405_adj_3764, n30439, n30022, n29287, n442_adj_3765, 
        n30232, n30021, n29286, n29285, n369_adj_3766, n30231, n30020, 
        n29284, n332_adj_3767, n30438, n296_adj_3768, n30230, n30019, 
        n29283, n29282, n223_adj_3769, n30229, n30018, n259_adj_3770, 
        n30437, n150_adj_3771, n30228, n30017, n30016, n29281, n186_adj_3772, 
        n30436, n8_adj_3773, n77_adj_3774, n30015, n44_adj_3775, n113_adj_3776;
    wire [5:0]n8062;
    
    wire n37137, n490_adj_3777, n30227, n30014;
    wire [4:0]n8070;
    
    wire n417_adj_3778, n30226, n30435, n30434, n344_adj_3779, n30225, 
        n30013, n30433, n30012, n271_adj_3780, n30224, n512_adj_3781, 
        n30011, n198_adj_3782, n30223, n30432, n56_adj_3783, n125_adj_3784, 
        n439_adj_3785, n30010;
    wire [23:0]n1_adj_3887;
    
    wire n28752, n28751, n366_adj_3787, n30009, n28750, n28749, 
        n293_adj_3790, n30008, n28748, n28747, n28746, n28745;
    wire [6:0]n8053;
    
    wire n560_adj_3795, n30222, n28744, n487_adj_3797, n30221, n28743, 
        n220_adj_3799, n30007, n28742, n28741, n28740, n28739, n548_adj_3804, 
        n30431, n147_adj_3805, n30006, n28738, n28737, n414_adj_3808, 
        n30220, n5_adj_3809, n74_adj_3810, n28736, n341_adj_3812, 
        n30219, n28735, n28734, n28733, n28732, n28731, n28730, 
        n475_adj_3820, n30430;
    wire [23:0]n1_adj_3888;
    
    wire n28729, n28728, n268_adj_3823, n30218, n28727, n402_adj_3825, 
        n30429, n28726, n28725, n28724, n28723, n28722, n28721, 
        n28720, n28719, n195_adj_3834, n30217, n28718, n53_adj_3836, 
        n122_adj_3837, n28717, n28716, n329_adj_3840, n30428, n30216, 
        n28715, n28714, n557_adj_3843, n30215, n28713, n28712, n28711, 
        n28710, n256_adj_3848, n30427, n28709, n28708, n484_adj_3851, 
        n30214, n28707, n28706, n28705, n28704, n411_adj_3858, n30213, 
        n183_adj_3859, n30426, n338_adj_3860, n30212, n41_adj_3861, 
        n110_adj_3862, n265_adj_3863, n30211, n30425, n192_adj_3865, 
        n30210, n50_adj_3866, n119_adj_3867, n30209, n28399, n28340;
    wire [2:0]n8380;
    
    wire n4_adj_3868;
    wire [3:0]n8374;
    
    wire n28374, n4_adj_3869, n6_adj_3870, n28297, n6_adj_3871;
    wire [3:0]n8077;
    wire [1:0]n8088;
    
    wire n4_adj_3872;
    wire [2:0]n8083;
    
    wire n12_adj_3873, n8_adj_3874, n11_adj_3875, n6_adj_3876, n28267, 
        n18_adj_3877, n13_adj_3878, n4_adj_3879, n28242, n28208, n4_adj_3880, 
        n28165, n137, n207, n68, n8_adj_3881, n6_adj_3882, n7_adj_3883, 
        n8_adj_3884, n4_adj_3885, n37855, n5_adj_3886;
    
    SB_CARRY add_3748_11 (.CI(n30423), .I0(n8304[8]), .I1(GND_net), .CO(n30424));
    SB_LUT4 add_3748_10_lut (.I0(GND_net), .I1(n8304[7]), .I2(GND_net), 
            .I3(n30422), .O(n8290[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12), .I1(n257[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3748_10 (.CI(n30422), .I0(n8304[7]), .I1(GND_net), .CO(n30423));
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3748_9_lut (.I0(GND_net), .I1(n8304[6]), .I2(GND_net), 
            .I3(n30421), .O(n8290[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3748_9 (.CI(n30421), .I0(n8304[6]), .I1(GND_net), .CO(n30422));
    SB_LUT4 add_3748_8_lut (.I0(GND_net), .I1(n8304[5]), .I2(n545), .I3(n30420), 
            .O(n8290[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_8_lut (.I0(GND_net), .I1(n8043[5]), .I2(n554), .I3(n30207), 
            .O(n8032[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3729_8 (.CI(n30207), .I0(n8043[5]), .I1(n554), .CO(n30208));
    SB_CARRY add_3748_8 (.CI(n30420), .I0(n8304[5]), .I1(n545), .CO(n30421));
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3729_7_lut (.I0(GND_net), .I1(n8043[4]), .I2(n481), .I3(n30206), 
            .O(n8032[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3748_7_lut (.I0(GND_net), .I1(n8304[4]), .I2(n472), .I3(n30419), 
            .O(n8290[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35487_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n41613), 
            .O(n42341));
    defparam i35487_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3729_7 (.CI(n30206), .I0(n8043[4]), .I1(n481), .CO(n30207));
    SB_LUT4 add_3729_6_lut (.I0(GND_net), .I1(n8043[3]), .I2(n408), .I3(n30205), 
            .O(n8032[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_24_lut (.I0(GND_net), .I1(n3054[22]), .I2(n3079[22]), 
            .I3(n28571), .O(duty_23__N_3478[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_24 (.CI(n28571), .I0(n3054[22]), .I1(n3079[22]), 
            .CO(n28572));
    SB_CARRY add_3748_7 (.CI(n30419), .I0(n8304[4]), .I1(n472), .CO(n30420));
    SB_CARRY add_3729_6 (.CI(n30205), .I0(n8043[3]), .I1(n408), .CO(n30206));
    SB_LUT4 i35445_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n42341), 
            .O(n42299));
    defparam i35445_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36349_4_lut (.I0(n25_c), .I1(n23_adj_3561), .I2(n21), .I3(n42299), 
            .O(n43203));
    defparam i36349_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35854_4_lut (.I0(n31), .I1(n29_adj_3562), .I2(n27), .I3(n43203), 
            .O(n42708));
    defparam i35854_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_3748_6_lut (.I0(GND_net), .I1(n8304[3]), .I2(n399), .I3(n30418), 
            .O(n8290[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_5_lut (.I0(GND_net), .I1(n8043[2]), .I2(n335), .I3(n30204), 
            .O(n8032[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3748_6 (.CI(n30418), .I0(n8304[3]), .I1(n399), .CO(n30419));
    SB_CARRY add_3729_5 (.CI(n30204), .I0(n8043[2]), .I1(n335), .CO(n30205));
    SB_LUT4 add_654_23_lut (.I0(GND_net), .I1(n3054[21]), .I2(n3079[21]), 
            .I3(n28570), .O(duty_23__N_3478[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n28702), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3748_5_lut (.I0(GND_net), .I1(n8304[2]), .I2(n326), .I3(n30417), 
            .O(n8290[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_4_lut (.I0(GND_net), .I1(n8043[1]), .I2(n262), .I3(n30203), 
            .O(n8032[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n28702), .I0(GND_net), .I1(n1[19]), 
            .CO(n28703));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n28701), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_654_23 (.CI(n28570), .I0(n3054[21]), .I1(n3079[21]), 
            .CO(n28571));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n28701), .I0(GND_net), .I1(n1[18]), 
            .CO(n28702));
    SB_LUT4 add_654_22_lut (.I0(GND_net), .I1(n3054[20]), .I2(n3079[20]), 
            .I3(n28569), .O(duty_23__N_3478[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3748_5 (.CI(n30417), .I0(n8304[2]), .I1(n326), .CO(n30418));
    SB_CARRY add_3729_4 (.CI(n30203), .I0(n8043[1]), .I1(n262), .CO(n30204));
    SB_LUT4 add_3729_3_lut (.I0(GND_net), .I1(n8043[0]), .I2(n189), .I3(n30202), 
            .O(n8032[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3748_4_lut (.I0(GND_net), .I1(n8304[1]), .I2(n253), .I3(n30416), 
            .O(n8290[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_3 (.CI(n30202), .I0(n8043[0]), .I1(n189), .CO(n30203));
    SB_CARRY add_3748_4 (.CI(n30416), .I0(n8304[1]), .I1(n253), .CO(n30417));
    SB_LUT4 add_3729_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n8032[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3748_3_lut (.I0(GND_net), .I1(n8304[0]), .I2(n180), .I3(n30415), 
            .O(n8290[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n30202));
    SB_CARRY add_3748_3 (.CI(n30415), .I0(n8304[0]), .I1(n180), .CO(n30416));
    SB_LUT4 add_3728_11_lut (.I0(GND_net), .I1(n8032[8]), .I2(GND_net), 
            .I3(n30201), .O(n8020[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3748_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8290[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_10_lut (.I0(GND_net), .I1(n8032[7]), .I2(GND_net), 
            .I3(n30200), .O(n8020[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3748_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n30415));
    SB_CARRY add_3728_10 (.CI(n30200), .I0(n8032[7]), .I1(GND_net), .CO(n30201));
    SB_LUT4 add_3747_14_lut (.I0(GND_net), .I1(n8290[11]), .I2(GND_net), 
            .I3(n30414), .O(n8275[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_9_lut (.I0(GND_net), .I1(n8032[6]), .I2(GND_net), 
            .I3(n30199), .O(n8020[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3747_13_lut (.I0(GND_net), .I1(n8290[10]), .I2(GND_net), 
            .I3(n30413), .O(n8275[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_9 (.CI(n30199), .I0(n8032[6]), .I1(GND_net), .CO(n30200));
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3564));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_13 (.CI(n30413), .I0(n8290[10]), .I1(GND_net), .CO(n30414));
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3565));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n28700), .O(n35_adj_3566)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n28700), .I0(GND_net), .I1(n1[17]), 
            .CO(n28701));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n28699), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n28699), .I0(GND_net), .I1(n1[16]), 
            .CO(n28700));
    SB_LUT4 add_3747_12_lut (.I0(GND_net), .I1(n8290[9]), .I2(GND_net), 
            .I3(n30412), .O(n8275[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n28698), .O(n31_adj_3568)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3570));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_3571));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36493_4_lut (.I0(n37_adj_3572), .I1(n35), .I2(n33_adj_3573), 
            .I3(n42708), .O(n43347));
    defparam i36493_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_3574));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_3576));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_3577));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_3578));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_652_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256), 
            .I3(GND_net), .O(n3079[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35904_3_lut (.I0(n6_adj_3580), .I1(n257[10]), .I2(n21), .I3(GND_net), 
            .O(n42758));   // verilog/motorControl.v(46[19:35])
    defparam i35904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35905_3_lut (.I0(n42758), .I1(n257[11]), .I2(n23_adj_3561), 
            .I3(GND_net), .O(n42759));   // verilog/motorControl.v(46[19:35])
    defparam i35905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_3582));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_3583));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_3584));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256), 
            .I3(GND_net), .O(n3079[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_652_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256), 
            .I3(GND_net), .O(n3079[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_12 (.CI(n30412), .I0(n8290[9]), .I1(GND_net), .CO(n30413));
    SB_LUT4 add_3747_11_lut (.I0(GND_net), .I1(n8290[8]), .I2(GND_net), 
            .I3(n30411), .O(n8275[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3747_11 (.CI(n30411), .I0(n8290[8]), .I1(GND_net), .CO(n30412));
    SB_LUT4 add_3747_10_lut (.I0(GND_net), .I1(n8290[7]), .I2(GND_net), 
            .I3(n30410), .O(n8275[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_10 (.CI(n30410), .I0(n8290[7]), .I1(GND_net), .CO(n30411));
    SB_CARRY add_654_22 (.CI(n28569), .I0(n3054[20]), .I1(n3079[20]), 
            .CO(n28570));
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3585));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256), 
            .I3(GND_net), .O(n3079[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3728_8_lut (.I0(GND_net), .I1(n8032[5]), .I2(n551), .I3(n30198), 
            .O(n8020[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3747_9_lut (.I0(GND_net), .I1(n8290[6]), .I2(GND_net), 
            .I3(n30409), .O(n8275[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_3588));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_654_21_lut (.I0(GND_net), .I1(n3054[19]), .I2(n3079[19]), 
            .I3(n28568), .O(duty_23__N_3478[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3589));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3590));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n28698), .I0(GND_net), .I1(n1[15]), 
            .CO(n28699));
    SB_LUT4 mux_652_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256), 
            .I3(GND_net), .O(n3079[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17), 
            .I3(GND_net), .O(n8_adj_3591));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n28697), .O(n29_adj_3592)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16), .I1(n257[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n28697), .I0(GND_net), .I1(n1[14]), 
            .CO(n28698));
    SB_CARRY add_3747_9 (.CI(n30409), .I0(n8290[6]), .I1(GND_net), .CO(n30410));
    SB_CARRY add_3728_8 (.CI(n30198), .I0(n8032[5]), .I1(n551), .CO(n30199));
    SB_LUT4 add_3747_8_lut (.I0(GND_net), .I1(n8290[5]), .I2(n542), .I3(n30408), 
            .O(n8275[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_7_lut (.I0(GND_net), .I1(n8032[4]), .I2(n478), .I3(n30197), 
            .O(n8020[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3747_8 (.CI(n30408), .I0(n8290[5]), .I1(n542), .CO(n30409));
    SB_CARRY add_3728_7 (.CI(n30197), .I0(n8032[4]), .I1(n478), .CO(n30198));
    SB_LUT4 i34610_4_lut (.I0(n43), .I1(n25_c), .I2(n23_adj_3561), .I3(n41563), 
            .O(n41463));
    defparam i34610_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3747_7_lut (.I0(GND_net), .I1(n8290[4]), .I2(n469), .I3(n30407), 
            .O(n8275[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n28696), .O(n27_adj_3594)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_654_21 (.CI(n28568), .I0(n3054[19]), .I1(n3079[19]), 
            .CO(n28569));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3355[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_654_20_lut (.I0(GND_net), .I1(n3054[18]), .I2(n3079[18]), 
            .I3(n28567), .O(duty_23__N_3478[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3596));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_7 (.CI(n30407), .I0(n8290[4]), .I1(n469), .CO(n30408));
    SB_LUT4 add_3728_6_lut (.I0(GND_net), .I1(n8032[3]), .I2(n405), .I3(n30196), 
            .O(n8020[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3747_6_lut (.I0(GND_net), .I1(n8290[3]), .I2(n396), .I3(n30406), 
            .O(n8275[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_6 (.CI(n30196), .I0(n8032[3]), .I1(n405), .CO(n30197));
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_6 (.CI(n30406), .I0(n8290[3]), .I1(n396), .CO(n30407));
    SB_LUT4 add_3728_5_lut (.I0(GND_net), .I1(n8032[2]), .I2(n332), .I3(n30195), 
            .O(n8020[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n28696), .I0(GND_net), .I1(n1[13]), 
            .CO(n28697));
    SB_LUT4 add_3747_5_lut (.I0(GND_net), .I1(n8290[2]), .I2(n323), .I3(n30405), 
            .O(n8275[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_5 (.CI(n30195), .I0(n8032[2]), .I1(n332), .CO(n30196));
    SB_CARRY add_3747_5 (.CI(n30405), .I0(n8290[2]), .I1(n323), .CO(n30406));
    SB_LUT4 add_3747_4_lut (.I0(GND_net), .I1(n8290[1]), .I2(n250), .I3(n30404), 
            .O(n8275[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_4_lut (.I0(GND_net), .I1(n8032[1]), .I2(n259_adj_3596), 
            .I3(n30194), .O(n8020[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3747_4 (.CI(n30404), .I0(n8290[1]), .I1(n250), .CO(n30405));
    SB_LUT4 add_3747_3_lut (.I0(GND_net), .I1(n8290[0]), .I2(n177), .I3(n30403), 
            .O(n8275[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_4 (.CI(n30194), .I0(n8032[1]), .I1(n259_adj_3596), 
            .CO(n30195));
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_3 (.CI(n30403), .I0(n8290[0]), .I1(n177), .CO(n30404));
    SB_LUT4 add_3747_2_lut (.I0(GND_net), .I1(n35_adj_3590), .I2(n104), 
            .I3(GND_net), .O(n8275[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3747_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3597));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3728_3_lut (.I0(GND_net), .I1(n8032[0]), .I2(n186_adj_3589), 
            .I3(n30193), .O(n8020[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_3 (.CI(n30193), .I0(n8032[0]), .I1(n186_adj_3589), 
            .CO(n30194));
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3747_2 (.CI(GND_net), .I0(n35_adj_3590), .I1(n104), .CO(n30403));
    SB_LUT4 add_3728_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n8020[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3746_15_lut (.I0(GND_net), .I1(n8275[12]), .I2(GND_net), 
            .I3(n30402), .O(n8259[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n30193));
    SB_LUT4 add_3746_14_lut (.I0(GND_net), .I1(n8275[11]), .I2(GND_net), 
            .I3(n30401), .O(n8259[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3727_12_lut (.I0(GND_net), .I1(n8020[9]), .I2(GND_net), 
            .I3(n30192), .O(n8007[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_14 (.CI(n30401), .I0(n8275[11]), .I1(GND_net), .CO(n30402));
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3598));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256), 
            .I3(GND_net), .O(n3079[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n28695), .O(n25_adj_3599)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3727_11_lut (.I0(GND_net), .I1(n8020[8]), .I2(GND_net), 
            .I3(n30191), .O(n8007[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3727_11 (.CI(n30191), .I0(n8020[8]), .I1(GND_net), .CO(n30192));
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3600));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3601));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3602));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3746_13_lut (.I0(GND_net), .I1(n8275[10]), .I2(GND_net), 
            .I3(n30400), .O(n8259[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3603));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3746_13 (.CI(n30400), .I0(n8275[10]), .I1(GND_net), .CO(n30401));
    SB_LUT4 add_3746_12_lut (.I0(GND_net), .I1(n8275[9]), .I2(GND_net), 
            .I3(n30399), .O(n8259[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3727_10_lut (.I0(GND_net), .I1(n8020[7]), .I2(GND_net), 
            .I3(n30190), .O(n8007[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_12 (.CI(n30399), .I0(n8275[9]), .I1(GND_net), .CO(n30400));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n28695), .I0(GND_net), .I1(n1[12]), 
            .CO(n28696));
    SB_LUT4 add_3746_11_lut (.I0(GND_net), .I1(n8275[8]), .I2(GND_net), 
            .I3(n30398), .O(n8259[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3604));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3727_10 (.CI(n30190), .I0(n8020[7]), .I1(GND_net), .CO(n30191));
    SB_CARRY add_3746_11 (.CI(n30398), .I0(n8275[8]), .I1(GND_net), .CO(n30399));
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3605));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3727_9_lut (.I0(GND_net), .I1(n8020[6]), .I2(GND_net), 
            .I3(n30189), .O(n8007[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n28694), .O(n23_adj_3606)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3607));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n28694), .I0(GND_net), .I1(n1[11]), 
            .CO(n28695));
    SB_LUT4 add_3746_10_lut (.I0(GND_net), .I1(n8275[7]), .I2(GND_net), 
            .I3(n30397), .O(n8259[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_9 (.CI(n30189), .I0(n8020[6]), .I1(GND_net), .CO(n30190));
    SB_CARRY add_3746_10 (.CI(n30397), .I0(n8275[7]), .I1(GND_net), .CO(n30398));
    SB_LUT4 add_3727_8_lut (.I0(GND_net), .I1(n8020[5]), .I2(n548), .I3(n30188), 
            .O(n8007[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n28693), .O(n21_adj_3608)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3609));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3746_9_lut (.I0(GND_net), .I1(n8275[6]), .I2(GND_net), 
            .I3(n30396), .O(n8259[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_20 (.CI(n28567), .I0(n3054[18]), .I1(n3079[18]), 
            .CO(n28568));
    SB_CARRY add_3727_8 (.CI(n30188), .I0(n8020[5]), .I1(n548), .CO(n30189));
    SB_LUT4 add_3727_7_lut (.I0(GND_net), .I1(n8020[4]), .I2(n475), .I3(n30187), 
            .O(n8007[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_19_lut (.I0(GND_net), .I1(n3054[17]), .I2(n3079[17]), 
            .I3(n28566), .O(duty_23__N_3478[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_9 (.CI(n30396), .I0(n8275[6]), .I1(GND_net), .CO(n30397));
    SB_LUT4 add_3746_8_lut (.I0(GND_net), .I1(n8275[5]), .I2(n539), .I3(n30395), 
            .O(n8259[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3610));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3746_8 (.CI(n30395), .I0(n8275[5]), .I1(n539), .CO(n30396));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n28693), .I0(GND_net), .I1(n1[10]), 
            .CO(n28694));
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3746_7_lut (.I0(GND_net), .I1(n8275[4]), .I2(n466), .I3(n30394), 
            .O(n8259[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_7 (.CI(n30187), .I0(n8020[4]), .I1(n475), .CO(n30188));
    SB_LUT4 add_3727_6_lut (.I0(GND_net), .I1(n8020[3]), .I2(n402), .I3(n30186), 
            .O(n8007[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_6 (.CI(n30186), .I0(n8020[3]), .I1(n402), .CO(n30187));
    SB_LUT4 add_3727_5_lut (.I0(GND_net), .I1(n8020[2]), .I2(n329), .I3(n30185), 
            .O(n8007[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_19 (.CI(n28566), .I0(n3054[17]), .I1(n3079[17]), 
            .CO(n28567));
    SB_CARRY add_3746_7 (.CI(n30394), .I0(n8275[4]), .I1(n466), .CO(n30395));
    SB_LUT4 add_3746_6_lut (.I0(GND_net), .I1(n8275[3]), .I2(n393), .I3(n30393), 
            .O(n8259[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3611));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3746_6 (.CI(n30393), .I0(n8275[3]), .I1(n393), .CO(n30394));
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3612));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36082_4_lut (.I0(n24), .I1(n8_adj_3591), .I2(n45), .I3(n41453), 
            .O(n42936));   // verilog/motorControl.v(46[19:35])
    defparam i36082_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3746_5_lut (.I0(GND_net), .I1(n8275[2]), .I2(n320), .I3(n30392), 
            .O(n8259[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_5 (.CI(n30392), .I0(n8275[2]), .I1(n320), .CO(n30393));
    SB_CARRY add_3727_5 (.CI(n30185), .I0(n8020[2]), .I1(n329), .CO(n30186));
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_3613));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3727_4_lut (.I0(GND_net), .I1(n8020[1]), .I2(n256_adj_3585), 
            .I3(n30184), .O(n8007[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3746_4_lut (.I0(GND_net), .I1(n8275[1]), .I2(n247), .I3(n30391), 
            .O(n8259[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_18_lut (.I0(GND_net), .I1(n3054[16]), .I2(n3079[16]), 
            .I3(n28565), .O(duty_23__N_3478[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_4 (.CI(n30184), .I0(n8020[1]), .I1(n256_adj_3585), 
            .CO(n30185));
    SB_CARRY add_3746_4 (.CI(n30391), .I0(n8275[1]), .I1(n247), .CO(n30392));
    SB_LUT4 add_3727_3_lut (.I0(GND_net), .I1(n8020[0]), .I2(n183), .I3(n30183), 
            .O(n8007[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35348_3_lut (.I0(n42759), .I1(n257[12]), .I2(n25_c), .I3(GND_net), 
            .O(n42202));   // verilog/motorControl.v(46[19:35])
    defparam i35348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n41179), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35900_3_lut (.I0(n4), .I1(n257[13]), .I2(n27), .I3(GND_net), 
            .O(n42754));   // verilog/motorControl.v(46[19:35])
    defparam i35900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3614));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3615));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3616));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3617));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3618));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3619));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3620));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3746_3_lut (.I0(GND_net), .I1(n8275[0]), .I2(n174), .I3(n30390), 
            .O(n8259[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_3 (.CI(n30183), .I0(n8020[0]), .I1(n183), .CO(n30184));
    SB_LUT4 add_3727_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n8007[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_3 (.CI(n30390), .I0(n8275[0]), .I1(n174), .CO(n30391));
    SB_CARRY add_3727_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n30183));
    SB_LUT4 i35901_3_lut (.I0(n42754), .I1(n257[14]), .I2(n29_adj_3562), 
            .I3(GND_net), .O(n42755));   // verilog/motorControl.v(46[19:35])
    defparam i35901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34669_4_lut (.I0(n33_adj_3573), .I1(n31), .I2(n29_adj_3562), 
            .I3(n41534), .O(n41522));
    defparam i34669_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36519_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n41519), 
            .O(n43373));   // verilog/motorControl.v(46[19:35])
    defparam i36519_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35350_3_lut (.I0(n42755), .I1(n257[15]), .I2(n31), .I3(GND_net), 
            .O(n42204));   // verilog/motorControl.v(46[19:35])
    defparam i35350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36602_4_lut (.I0(n42204), .I1(n43373), .I2(n35), .I3(n41522), 
            .O(n43456));   // verilog/motorControl.v(46[19:35])
    defparam i36602_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36603_3_lut (.I0(n43456), .I1(n257[18]), .I2(n37_adj_3572), 
            .I3(GND_net), .O(n43457));   // verilog/motorControl.v(46[19:35])
    defparam i36603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36579_3_lut (.I0(n43457), .I1(n257[19]), .I2(n39_adj_3622), 
            .I3(GND_net), .O(n43433));   // verilog/motorControl.v(46[19:35])
    defparam i36579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34615_4_lut (.I0(n43), .I1(n41_adj_3623), .I2(n39_adj_3622), 
            .I3(n43347), .O(n41468));
    defparam i34615_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3624));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3625));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3626));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34887_4_lut (.I0(n21_adj_3626), .I1(n19_adj_3625), .I2(n17_adj_3624), 
            .I3(n9_adj_3620), .O(n41741));
    defparam i34887_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34866_4_lut (.I0(n27_adj_3619), .I1(n15_adj_3618), .I2(n13_adj_3617), 
            .I3(n11_adj_3616), .O(n41720));
    defparam i34866_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3726_13_lut (.I0(GND_net), .I1(n8007[10]), .I2(GND_net), 
            .I3(n30182), .O(n7993[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_18 (.CI(n28565), .I0(n3054[16]), .I1(n3079[16]), 
            .CO(n28566));
    SB_LUT4 i36329_4_lut (.I0(n42202), .I1(n42936), .I2(n45), .I3(n41463), 
            .O(n43183));   // verilog/motorControl.v(46[19:35])
    defparam i36329_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36548_3_lut (.I0(n43433), .I1(n257[20]), .I2(n41_adj_3623), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(46[19:35])
    defparam i36548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n28692), .O(n19_adj_3627)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3746_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8259[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3746_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_17_lut (.I0(GND_net), .I1(n3054[15]), .I2(n3079[15]), 
            .I3(n28564), .O(duty_23__N_3478[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3746_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n30390));
    SB_LUT4 add_3745_16_lut (.I0(GND_net), .I1(n8259[13]), .I2(GND_net), 
            .I3(n30389), .O(n8242[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3745_15_lut (.I0(GND_net), .I1(n8259[12]), .I2(GND_net), 
            .I3(n30388), .O(n8242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_15 (.CI(n30388), .I0(n8259[12]), .I1(GND_net), .CO(n30389));
    SB_LUT4 add_3745_14_lut (.I0(GND_net), .I1(n8259[11]), .I2(GND_net), 
            .I3(n30387), .O(n8242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3726_12_lut (.I0(GND_net), .I1(n8007[9]), .I2(GND_net), 
            .I3(n30181), .O(n7993[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n28692), .I0(GND_net), .I1(n1[9]), 
            .CO(n28693));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n28691), .O(n17_adj_3628)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3726_12 (.CI(n30181), .I0(n8007[9]), .I1(GND_net), .CO(n30182));
    SB_LUT4 add_3726_11_lut (.I0(GND_net), .I1(n8007[8]), .I2(GND_net), 
            .I3(n30180), .O(n7993[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_14 (.CI(n30387), .I0(n8259[11]), .I1(GND_net), .CO(n30388));
    SB_CARRY add_3726_11 (.CI(n30180), .I0(n8007[8]), .I1(GND_net), .CO(n30181));
    SB_LUT4 add_3745_13_lut (.I0(GND_net), .I1(n8259[10]), .I2(GND_net), 
            .I3(n30386), .O(n8242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3726_10_lut (.I0(GND_net), .I1(n8007[7]), .I2(GND_net), 
            .I3(n30179), .O(n7993[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_13 (.CI(n30386), .I0(n8259[10]), .I1(GND_net), .CO(n30387));
    SB_LUT4 add_3745_12_lut (.I0(GND_net), .I1(n8259[9]), .I2(GND_net), 
            .I3(n30385), .O(n8242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_10 (.CI(n30179), .I0(n8007[7]), .I1(GND_net), .CO(n30180));
    SB_LUT4 add_3726_9_lut (.I0(GND_net), .I1(n8007[6]), .I2(GND_net), 
            .I3(n30178), .O(n7993[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_9 (.CI(n30178), .I0(n8007[6]), .I1(GND_net), .CO(n30179));
    SB_CARRY add_3745_12 (.CI(n30385), .I0(n8259[9]), .I1(GND_net), .CO(n30386));
    SB_LUT4 add_3726_8_lut (.I0(GND_net), .I1(n8007[5]), .I2(n545_adj_3578), 
            .I3(n30177), .O(n7993[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36331_4_lut (.I0(n40), .I1(n43183), .I2(n45), .I3(n41468), 
            .O(n43185));   // verilog/motorControl.v(46[19:35])
    defparam i36331_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36332_3_lut (.I0(n43185), .I1(duty[23]), .I2(n47_adj_3629), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(46[19:35])
    defparam i36332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256), 
            .I3(GND_net), .O(n3079[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n28691), .I0(GND_net), .I1(n1[8]), 
            .CO(n28692));
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_3630), .I1(duty[17]), .I2(n35_adj_3614), 
            .I3(GND_net), .O(n30_adj_3631));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3745_11_lut (.I0(GND_net), .I1(n8259[8]), .I2(GND_net), 
            .I3(n30384), .O(n8242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_11 (.CI(n30384), .I0(n8259[8]), .I1(GND_net), .CO(n30385));
    SB_CARRY add_3726_8 (.CI(n30177), .I0(n8007[5]), .I1(n545_adj_3578), 
            .CO(n30178));
    SB_LUT4 add_3745_10_lut (.I0(GND_net), .I1(n8259[7]), .I2(GND_net), 
            .I3(n30383), .O(n8242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35583_4_lut (.I0(n13_adj_3617), .I1(n11_adj_3616), .I2(n9_adj_3620), 
            .I3(n41789), .O(n42437));
    defparam i35583_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35573_4_lut (.I0(n19_adj_3625), .I1(n17_adj_3624), .I2(n15_adj_3618), 
            .I3(n42437), .O(n42427));
    defparam i35573_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36394_4_lut (.I0(n25_adj_3612), .I1(n23_adj_3611), .I2(n21_adj_3626), 
            .I3(n42427), .O(n43248));
    defparam i36394_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3745_10 (.CI(n30383), .I0(n8259[7]), .I1(GND_net), .CO(n30384));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n28690), .O(n15_adj_3632)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35930_4_lut (.I0(n31_adj_3610), .I1(n29_adj_3609), .I2(n27_adj_3619), 
            .I3(n43248), .O(n42784));
    defparam i35930_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36506_4_lut (.I0(n37_adj_3607), .I1(n35_adj_3614), .I2(n33_adj_3615), 
            .I3(n42784), .O(n43360));
    defparam i36506_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3726_7_lut (.I0(GND_net), .I1(n8007[4]), .I2(n472_adj_3577), 
            .I3(n30176), .O(n7993[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3745_9_lut (.I0(GND_net), .I1(n8259[6]), .I2(GND_net), 
            .I3(n30382), .O(n8242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_7 (.CI(n30176), .I0(n8007[4]), .I1(n472_adj_3577), 
            .CO(n30177));
    SB_LUT4 add_3726_6_lut (.I0(GND_net), .I1(n8007[3]), .I2(n399_adj_3576), 
            .I3(n30175), .O(n7993[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_9 (.CI(n30382), .I0(n8259[6]), .I1(GND_net), .CO(n30383));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n28690), .I0(GND_net), .I1(n1[7]), 
            .CO(n28691));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n28689), .O(n13_adj_3633)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3745_8_lut (.I0(GND_net), .I1(n8259[5]), .I2(n536), .I3(n30381), 
            .O(n8242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_6 (.CI(n30175), .I0(n8007[3]), .I1(n399_adj_3576), 
            .CO(n30176));
    SB_LUT4 add_3726_5_lut (.I0(GND_net), .I1(n8007[2]), .I2(n326_adj_3574), 
            .I3(n30174), .O(n7993[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_5 (.CI(n30174), .I0(n8007[2]), .I1(n326_adj_3574), 
            .CO(n30175));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n28689), .I0(GND_net), .I1(n1[6]), 
            .CO(n28690));
    SB_CARRY add_3745_8 (.CI(n30381), .I0(n8259[5]), .I1(n536), .CO(n30382));
    SB_LUT4 add_3745_7_lut (.I0(GND_net), .I1(n8259[4]), .I2(n463), .I3(n30380), 
            .O(n8242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3726_4_lut (.I0(GND_net), .I1(n8007[1]), .I2(n253_adj_3571), 
            .I3(n30173), .O(n7993[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_4 (.CI(n30173), .I0(n8007[1]), .I1(n253_adj_3571), 
            .CO(n30174));
    SB_LUT4 i36193_3_lut (.I0(n6_adj_3634), .I1(duty[10]), .I2(n21_adj_3626), 
            .I3(GND_net), .O(n43047));   // verilog/motorControl.v(44[10:25])
    defparam i36193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36194_3_lut (.I0(n43047), .I1(duty[11]), .I2(n23_adj_3611), 
            .I3(GND_net), .O(n43048));   // verilog/motorControl.v(44[10:25])
    defparam i36194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3745_7 (.CI(n30380), .I0(n8259[4]), .I1(n463), .CO(n30381));
    SB_LUT4 add_3726_3_lut (.I0(GND_net), .I1(n8007[0]), .I2(n180_adj_3570), 
            .I3(n30172), .O(n7993[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n28688), .O(n11_adj_3635)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3745_6_lut (.I0(GND_net), .I1(n8259[3]), .I2(n390), .I3(n30379), 
            .O(n8242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_3636), .I1(duty[22]), .I2(n45_adj_3604), 
            .I3(GND_net), .O(n24_adj_3637));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34770_4_lut (.I0(n43_adj_3605), .I1(n25_adj_3612), .I2(n23_adj_3611), 
            .I3(n41741), .O(n41623));
    defparam i34770_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36078_4_lut (.I0(n24_adj_3637), .I1(n8_adj_3638), .I2(n45_adj_3604), 
            .I3(n41619), .O(n42932));   // verilog/motorControl.v(44[10:25])
    defparam i36078_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3745_6 (.CI(n30379), .I0(n8259[3]), .I1(n390), .CO(n30380));
    SB_CARRY add_3726_3 (.CI(n30172), .I0(n8007[0]), .I1(n180_adj_3570), 
            .CO(n30173));
    SB_LUT4 i35338_3_lut (.I0(n43048), .I1(duty[12]), .I2(n25_adj_3612), 
            .I3(GND_net), .O(n42192));   // verilog/motorControl.v(44[10:25])
    defparam i35338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3745_5_lut (.I0(GND_net), .I1(n8259[2]), .I2(n317), .I3(n30378), 
            .O(n8242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_3639));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i36191_3_lut (.I0(n4_adj_3639), .I1(duty[13]), .I2(n27_adj_3619), 
            .I3(GND_net), .O(n43045));   // verilog/motorControl.v(44[10:25])
    defparam i36191_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3745_5 (.CI(n30378), .I0(n8259[2]), .I1(n317), .CO(n30379));
    SB_LUT4 i36192_3_lut (.I0(n43045), .I1(duty[14]), .I2(n29_adj_3609), 
            .I3(GND_net), .O(n43046));   // verilog/motorControl.v(44[10:25])
    defparam i36192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3726_2_lut (.I0(GND_net), .I1(n38_adj_3565), .I2(n107_adj_3564), 
            .I3(GND_net), .O(n7993[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3745_4_lut (.I0(GND_net), .I1(n8259[1]), .I2(n244), .I3(n30377), 
            .O(n8242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3640));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n28688), .I0(GND_net), .I1(n1[5]), 
            .CO(n28689));
    SB_CARRY add_654_17 (.CI(n28564), .I0(n3054[15]), .I1(n3079[15]), 
            .CO(n28565));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n28687), .O(n9_adj_3641)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3642));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34842_4_lut (.I0(n33_adj_3615), .I1(n31_adj_3610), .I2(n29_adj_3609), 
            .I3(n41720), .O(n41696));
    defparam i34842_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n28687), .I0(GND_net), .I1(n1[4]), 
            .CO(n28688));
    SB_CARRY add_3726_2 (.CI(GND_net), .I0(n38_adj_3565), .I1(n107_adj_3564), 
            .CO(n30172));
    SB_CARRY add_3745_4 (.CI(n30377), .I0(n8259[1]), .I1(n244), .CO(n30378));
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_3643));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3745_3_lut (.I0(GND_net), .I1(n8259[0]), .I2(n171), .I3(n30376), 
            .O(n8242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3745_3 (.CI(n30376), .I0(n8259[0]), .I1(n171), .CO(n30377));
    SB_LUT4 i36434_4_lut (.I0(n30_adj_3631), .I1(n10_adj_3644), .I2(n35_adj_3614), 
            .I3(n41692), .O(n43288));   // verilog/motorControl.v(44[10:25])
    defparam i36434_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_3645));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3725_14_lut (.I0(GND_net), .I1(n7993[11]), .I2(GND_net), 
            .I3(n30171), .O(n7978[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3725_13_lut (.I0(GND_net), .I1(n7993[10]), .I2(GND_net), 
            .I3(n30170), .O(n7978[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35340_3_lut (.I0(n43046), .I1(duty[15]), .I2(n31_adj_3610), 
            .I3(GND_net), .O(n42194));   // verilog/motorControl.v(44[10:25])
    defparam i35340_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3725_13 (.CI(n30170), .I0(n7993[10]), .I1(GND_net), .CO(n30171));
    SB_LUT4 add_3745_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n8242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3745_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36572_4_lut (.I0(n42194), .I1(n43288), .I2(n35_adj_3614), 
            .I3(n41696), .O(n43426));   // verilog/motorControl.v(44[10:25])
    defparam i36572_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3745_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n30376));
    SB_LUT4 i36573_3_lut (.I0(n43426), .I1(duty[18]), .I2(n37_adj_3607), 
            .I3(GND_net), .O(n43427));   // verilog/motorControl.v(44[10:25])
    defparam i36573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36561_3_lut (.I0(n43427), .I1(duty[19]), .I2(n39_adj_3602), 
            .I3(GND_net), .O(n43415));   // verilog/motorControl.v(44[10:25])
    defparam i36561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n28686), .O(n7_adj_3646)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n28686), .I0(GND_net), .I1(n1[3]), 
            .CO(n28687));
    SB_LUT4 i34772_4_lut (.I0(n43_adj_3605), .I1(n41_adj_3601), .I2(n39_adj_3602), 
            .I3(n43360), .O(n41625));
    defparam i34772_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3725_12_lut (.I0(GND_net), .I1(n7993[9]), .I2(GND_net), 
            .I3(n30169), .O(n7978[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36489_4_lut (.I0(n42192), .I1(n42932), .I2(n45_adj_3604), 
            .I3(n41623), .O(n43343));   // verilog/motorControl.v(44[10:25])
    defparam i36489_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35346_3_lut (.I0(n43415), .I1(duty[20]), .I2(n41_adj_3601), 
            .I3(GND_net), .O(n42200));   // verilog/motorControl.v(44[10:25])
    defparam i35346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36491_4_lut (.I0(n42200), .I1(n43343), .I2(n45_adj_3604), 
            .I3(n41625), .O(n43345));   // verilog/motorControl.v(44[10:25])
    defparam i36491_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n28685), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3744_17_lut (.I0(GND_net), .I1(n8242[14]), .I2(GND_net), 
            .I3(n30375), .O(n8224[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3744_16_lut (.I0(GND_net), .I1(n8242[13]), .I2(GND_net), 
            .I3(n30374), .O(n8224[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n28685), .I0(GND_net), .I1(n1[2]), 
            .CO(n28686));
    SB_LUT4 mux_652_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256), 
            .I3(GND_net), .O(n3079[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36492_3_lut (.I0(n43345), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3502));   // verilog/motorControl.v(44[10:25])
    defparam i36492_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n28684), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_654_16_lut (.I0(GND_net), .I1(n3054[14]), .I2(n3079[14]), 
            .I3(n28563), .O(duty_23__N_3478[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_12 (.CI(n30169), .I0(n7993[9]), .I1(GND_net), .CO(n30170));
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_3648));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3478[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_654_16 (.CI(n28563), .I0(n3054[14]), .I1(n3079[14]), 
            .CO(n28564));
    SB_CARRY add_3744_16 (.CI(n30374), .I0(n8242[13]), .I1(GND_net), .CO(n30375));
    SB_LUT4 add_3744_15_lut (.I0(GND_net), .I1(n8242[12]), .I2(GND_net), 
            .I3(n30373), .O(n8224[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_15_lut (.I0(GND_net), .I1(n3054[13]), .I2(n3079[13]), 
            .I3(n28562), .O(duty_23__N_3478[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n28684), .I0(GND_net), .I1(n1[1]), 
            .CO(n28685));
    SB_CARRY add_3744_15 (.CI(n30373), .I0(n8242[12]), .I1(GND_net), .CO(n30374));
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_3649));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3725_11_lut (.I0(GND_net), .I1(n7993[8]), .I2(GND_net), 
            .I3(n30168), .O(n7978[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3725_11 (.CI(n30168), .I0(n7993[8]), .I1(GND_net), .CO(n30169));
    SB_LUT4 add_3725_10_lut (.I0(GND_net), .I1(n7993[7]), .I2(GND_net), 
            .I3(n30167), .O(n7978[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3744_14_lut (.I0(GND_net), .I1(n8242[11]), .I2(GND_net), 
            .I3(n30372), .O(n8224[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_14 (.CI(n30372), .I0(n8242[11]), .I1(GND_net), .CO(n30373));
    SB_CARRY add_3725_10 (.CI(n30167), .I0(n7993[7]), .I1(GND_net), .CO(n30168));
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3725_9_lut (.I0(GND_net), .I1(n7993[6]), .I2(GND_net), 
            .I3(n30166), .O(n7978[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_9 (.CI(n30166), .I0(n7993[6]), .I1(GND_net), .CO(n30167));
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3744_13_lut (.I0(GND_net), .I1(n8242[10]), .I2(GND_net), 
            .I3(n30371), .O(n8224[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_13 (.CI(n30371), .I0(n8242[10]), .I1(GND_net), .CO(n30372));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3454 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n28684));
    SB_LUT4 mux_652_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n3079[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i19973_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n3054[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i19973_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_3651));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3744_12_lut (.I0(GND_net), .I1(n8242[9]), .I2(GND_net), 
            .I3(n30370), .O(n8224[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3725_8_lut (.I0(GND_net), .I1(n7993[5]), .I2(n542_adj_3652), 
            .I3(n30165), .O(n7978[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_8 (.CI(n30165), .I0(n7993[5]), .I1(n542_adj_3652), 
            .CO(n30166));
    SB_LUT4 add_3725_7_lut (.I0(GND_net), .I1(n7993[4]), .I2(n469_adj_3653), 
            .I3(n30164), .O(n7978[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_7 (.CI(n30164), .I0(n7993[4]), .I1(n469_adj_3653), 
            .CO(n30165));
    SB_LUT4 add_3725_6_lut (.I0(GND_net), .I1(n7993[3]), .I2(n396_adj_3654), 
            .I3(n30163), .O(n7978[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_12 (.CI(n30370), .I0(n8242[9]), .I1(GND_net), .CO(n30371));
    SB_LUT4 add_3744_11_lut (.I0(GND_net), .I1(n8242[8]), .I2(GND_net), 
            .I3(n30369), .O(n8224[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_15 (.CI(n28562), .I0(n3054[13]), .I1(n3079[13]), 
            .CO(n28563));
    SB_CARRY add_3725_6 (.CI(n30163), .I0(n7993[3]), .I1(n396_adj_3654), 
            .CO(n30164));
    SB_LUT4 add_3725_5_lut (.I0(GND_net), .I1(n7993[2]), .I2(n323_adj_3655), 
            .I3(n30162), .O(n7978[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_11 (.CI(n30369), .I0(n8242[8]), .I1(GND_net), .CO(n30370));
    SB_LUT4 add_3744_10_lut (.I0(GND_net), .I1(n8242[7]), .I2(GND_net), 
            .I3(n30368), .O(n8224[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_14_lut (.I0(GND_net), .I1(n3054[12]), .I2(n3079[12]), 
            .I3(n28561), .O(duty_23__N_3478[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_10 (.CI(n30368), .I0(n8242[7]), .I1(GND_net), .CO(n30369));
    SB_LUT4 add_3744_9_lut (.I0(GND_net), .I1(n8242[6]), .I2(GND_net), 
            .I3(n30367), .O(n8224[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_9 (.CI(n30367), .I0(n8242[6]), .I1(GND_net), .CO(n30368));
    SB_LUT4 add_3744_8_lut (.I0(GND_net), .I1(n8242[5]), .I2(n533), .I3(n30366), 
            .O(n8224[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_5 (.CI(n30162), .I0(n7993[2]), .I1(n323_adj_3655), 
            .CO(n30163));
    SB_LUT4 add_3725_4_lut (.I0(GND_net), .I1(n7993[1]), .I2(n250_adj_3656), 
            .I3(n30161), .O(n7978[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_4 (.CI(n30161), .I0(n7993[1]), .I1(n250_adj_3656), 
            .CO(n30162));
    SB_LUT4 add_3725_3_lut (.I0(GND_net), .I1(n7993[0]), .I2(n177_adj_3657), 
            .I3(n30160), .O(n7978[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_14 (.CI(n28561), .I0(n3054[12]), .I1(n3079[12]), 
            .CO(n28562));
    SB_CARRY add_3725_3 (.CI(n30160), .I0(n7993[0]), .I1(n177_adj_3657), 
            .CO(n30161));
    SB_CARRY add_3744_8 (.CI(n30366), .I0(n8242[5]), .I1(n533), .CO(n30367));
    SB_LUT4 add_3725_2_lut (.I0(GND_net), .I1(n35_adj_3658), .I2(n104_adj_3659), 
            .I3(GND_net), .O(n7978[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3744_7_lut (.I0(GND_net), .I1(n8242[4]), .I2(n460), .I3(n30365), 
            .O(n8224[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_2 (.CI(GND_net), .I0(n35_adj_3658), .I1(n104_adj_3659), 
            .CO(n30160));
    SB_LUT4 add_654_13_lut (.I0(GND_net), .I1(n3054[11]), .I2(n3079[11]), 
            .I3(n28560), .O(duty_23__N_3478[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_652_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256), 
            .I3(GND_net), .O(n3079[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3744_7 (.CI(n30365), .I0(n8242[4]), .I1(n460), .CO(n30366));
    SB_LUT4 add_3744_6_lut (.I0(GND_net), .I1(n8242[3]), .I2(n387), .I3(n30364), 
            .O(n8224[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3744_6 (.CI(n30364), .I0(n8242[3]), .I1(n387), .CO(n30365));
    SB_LUT4 add_3724_15_lut (.I0(GND_net), .I1(n7978[12]), .I2(GND_net), 
            .I3(n30159), .O(n7962[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3744_5_lut (.I0(GND_net), .I1(n8242[2]), .I2(n314), .I3(n30363), 
            .O(n8224[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_5 (.CI(n30363), .I0(n8242[2]), .I1(n314), .CO(n30364));
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3744_4_lut (.I0(GND_net), .I1(n8242[1]), .I2(n241_adj_3660), 
            .I3(n30362), .O(n8224[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3661));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3744_4 (.CI(n30362), .I0(n8242[1]), .I1(n241_adj_3660), 
            .CO(n30363));
    SB_LUT4 add_3724_14_lut (.I0(GND_net), .I1(n7978[11]), .I2(GND_net), 
            .I3(n30158), .O(n7962[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_13 (.CI(n28560), .I0(n3054[11]), .I1(n3079[11]), 
            .CO(n28561));
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3662));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_3663));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3744_3_lut (.I0(GND_net), .I1(n8242[0]), .I2(n168_adj_3664), 
            .I3(n30361), .O(n8224[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_14 (.CI(n30158), .I0(n7978[11]), .I1(GND_net), .CO(n30159));
    SB_LUT4 add_3724_13_lut (.I0(GND_net), .I1(n7978[10]), .I2(GND_net), 
            .I3(n30157), .O(n7962[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_3 (.CI(n30361), .I0(n8242[0]), .I1(n168_adj_3664), 
            .CO(n30362));
    SB_CARRY add_3724_13 (.CI(n30157), .I0(n7978[10]), .I1(GND_net), .CO(n30158));
    SB_LUT4 add_654_12_lut (.I0(GND_net), .I1(n3054[10]), .I2(n3079[10]), 
            .I3(n28559), .O(duty_23__N_3478[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3744_2_lut (.I0(GND_net), .I1(n26_adj_3665), .I2(n95_adj_3666), 
            .I3(GND_net), .O(n8224[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_12_lut (.I0(GND_net), .I1(n7978[9]), .I2(GND_net), 
            .I3(n30156), .O(n7962[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_12 (.CI(n28559), .I0(n3054[10]), .I1(n3079[10]), 
            .CO(n28560));
    SB_CARRY add_3724_12 (.CI(n30156), .I0(n7978[9]), .I1(GND_net), .CO(n30157));
    SB_CARRY add_3744_2 (.CI(GND_net), .I0(n26_adj_3665), .I1(n95_adj_3666), 
            .CO(n30361));
    SB_LUT4 add_3743_18_lut (.I0(GND_net), .I1(n8224[15]), .I2(GND_net), 
            .I3(n30360), .O(n8205[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_11_lut (.I0(GND_net), .I1(n7978[8]), .I2(GND_net), 
            .I3(n30155), .O(n7962[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_11 (.CI(n30155), .I0(n7978[8]), .I1(GND_net), .CO(n30156));
    SB_LUT4 add_3743_17_lut (.I0(GND_net), .I1(n8224[14]), .I2(GND_net), 
            .I3(n30359), .O(n8205[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_17 (.CI(n30359), .I0(n8224[14]), .I1(GND_net), .CO(n30360));
    SB_LUT4 add_3743_16_lut (.I0(GND_net), .I1(n8224[13]), .I2(GND_net), 
            .I3(n30358), .O(n8205[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_10_lut (.I0(GND_net), .I1(n7978[7]), .I2(GND_net), 
            .I3(n30154), .O(n7962[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_11_lut (.I0(GND_net), .I1(n3054[9]), .I2(n3079[9]), 
            .I3(n28558), .O(duty_23__N_3478[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_16 (.CI(n30358), .I0(n8224[13]), .I1(GND_net), .CO(n30359));
    SB_CARRY add_3724_10 (.CI(n30154), .I0(n7978[7]), .I1(GND_net), .CO(n30155));
    SB_LUT4 add_3743_15_lut (.I0(GND_net), .I1(n8224[12]), .I2(GND_net), 
            .I3(n30357), .O(n8205[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_23_lut (.I0(GND_net), .I1(n7822[20]), .I2(GND_net), 
            .I3(n29693), .O(n7798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_9_lut (.I0(GND_net), .I1(n7978[6]), .I2(GND_net), 
            .I3(n30153), .O(n7962[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_11 (.CI(n28558), .I0(n3054[9]), .I1(n3079[9]), .CO(n28559));
    SB_LUT4 add_3716_22_lut (.I0(GND_net), .I1(n7822[19]), .I2(GND_net), 
            .I3(n29692), .O(n7798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_9 (.CI(n30153), .I0(n7978[6]), .I1(GND_net), .CO(n30154));
    SB_LUT4 add_3724_8_lut (.I0(GND_net), .I1(n7978[5]), .I2(n539_adj_3667), 
            .I3(n30152), .O(n7962[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_15 (.CI(n30357), .I0(n8224[12]), .I1(GND_net), .CO(n30358));
    SB_CARRY add_3716_22 (.CI(n29692), .I0(n7822[19]), .I1(GND_net), .CO(n29693));
    SB_LUT4 add_3743_14_lut (.I0(GND_net), .I1(n8224[11]), .I2(GND_net), 
            .I3(n30356), .O(n8205[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_8 (.CI(n30152), .I0(n7978[5]), .I1(n539_adj_3667), 
            .CO(n30153));
    SB_LUT4 add_3724_7_lut (.I0(GND_net), .I1(n7978[4]), .I2(n466_adj_3668), 
            .I3(n30151), .O(n7962[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_21_lut (.I0(GND_net), .I1(n7822[18]), .I2(GND_net), 
            .I3(n29691), .O(n7798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_14 (.CI(n30356), .I0(n8224[11]), .I1(GND_net), .CO(n30357));
    SB_CARRY add_3724_7 (.CI(n30151), .I0(n7978[4]), .I1(n466_adj_3668), 
            .CO(n30152));
    SB_CARRY add_3716_21 (.CI(n29691), .I0(n7822[18]), .I1(GND_net), .CO(n29692));
    SB_LUT4 add_3716_20_lut (.I0(GND_net), .I1(n7822[17]), .I2(GND_net), 
            .I3(n29690), .O(n7798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_20 (.CI(n29690), .I0(n7822[17]), .I1(GND_net), .CO(n29691));
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_3669));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3716_19_lut (.I0(GND_net), .I1(n7822[16]), .I2(GND_net), 
            .I3(n29689), .O(n7798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_19 (.CI(n29689), .I0(n7822[16]), .I1(GND_net), .CO(n29690));
    SB_LUT4 add_3743_13_lut (.I0(GND_net), .I1(n8224[10]), .I2(GND_net), 
            .I3(n30355), .O(n8205[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_13 (.CI(n30355), .I0(n8224[10]), .I1(GND_net), .CO(n30356));
    SB_LUT4 add_3724_6_lut (.I0(GND_net), .I1(n7978[3]), .I2(n393_adj_3669), 
            .I3(n30150), .O(n7962[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3743_12_lut (.I0(GND_net), .I1(n8224[9]), .I2(GND_net), 
            .I3(n30354), .O(n8205[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_3668));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_3667));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3743_12 (.CI(n30354), .I0(n8224[9]), .I1(GND_net), .CO(n30355));
    SB_LUT4 add_3743_11_lut (.I0(GND_net), .I1(n8224[8]), .I2(GND_net), 
            .I3(n30353), .O(n8205[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_11 (.CI(n30353), .I0(n8224[8]), .I1(GND_net), .CO(n30354));
    SB_LUT4 add_3716_18_lut (.I0(GND_net), .I1(n7822[15]), .I2(GND_net), 
            .I3(n29688), .O(n7798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_18 (.CI(n29688), .I0(n7822[15]), .I1(GND_net), .CO(n29689));
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3670));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3724_6 (.CI(n30150), .I0(n7978[3]), .I1(n393_adj_3669), 
            .CO(n30151));
    SB_LUT4 add_3724_5_lut (.I0(GND_net), .I1(n7978[2]), .I2(n320_adj_3651), 
            .I3(n30149), .O(n7962[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3716_17_lut (.I0(GND_net), .I1(n7822[14]), .I2(GND_net), 
            .I3(n29687), .O(n7798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_17 (.CI(n29687), .I0(n7822[14]), .I1(GND_net), .CO(n29688));
    SB_LUT4 add_3716_16_lut (.I0(GND_net), .I1(n7822[13]), .I2(GND_net), 
            .I3(n29686), .O(n7798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3743_10_lut (.I0(GND_net), .I1(n8224[7]), .I2(GND_net), 
            .I3(n30352), .O(n8205[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_10 (.CI(n30352), .I0(n8224[7]), .I1(GND_net), .CO(n30353));
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_3671));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3724_5 (.CI(n30149), .I0(n7978[2]), .I1(n320_adj_3651), 
            .CO(n30150));
    SB_LUT4 add_654_10_lut (.I0(GND_net), .I1(n3054[8]), .I2(n3079[8]), 
            .I3(n28557), .O(duty_23__N_3478[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_16 (.CI(n29686), .I0(n7822[13]), .I1(GND_net), .CO(n29687));
    SB_LUT4 add_3724_4_lut (.I0(GND_net), .I1(n7978[1]), .I2(n247_adj_3645), 
            .I3(n30148), .O(n7962[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3743_9_lut (.I0(GND_net), .I1(n8224[6]), .I2(GND_net), 
            .I3(n30351), .O(n8205[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_15_lut (.I0(GND_net), .I1(n7822[12]), .I2(GND_net), 
            .I3(n29685), .O(n7798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_9 (.CI(n30351), .I0(n8224[6]), .I1(GND_net), .CO(n30352));
    SB_LUT4 add_3743_8_lut (.I0(GND_net), .I1(n8224[5]), .I2(n530), .I3(n30350), 
            .O(n8205[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_4 (.CI(n30148), .I0(n7978[1]), .I1(n247_adj_3645), 
            .CO(n30149));
    SB_CARRY add_3743_8 (.CI(n30350), .I0(n8224[5]), .I1(n530), .CO(n30351));
    SB_LUT4 add_3743_7_lut (.I0(GND_net), .I1(n8224[4]), .I2(n457), .I3(n30349), 
            .O(n8205[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_3_lut (.I0(GND_net), .I1(n7978[0]), .I2(n174_adj_3613), 
            .I3(n30147), .O(n7962[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_7 (.CI(n30349), .I0(n8224[4]), .I1(n457), .CO(n30350));
    SB_CARRY add_3724_3 (.CI(n30147), .I0(n7978[0]), .I1(n174_adj_3613), 
            .CO(n30148));
    SB_CARRY add_3716_15 (.CI(n29685), .I0(n7822[12]), .I1(GND_net), .CO(n29686));
    SB_LUT4 add_3716_14_lut (.I0(GND_net), .I1(n7822[11]), .I2(GND_net), 
            .I3(n29684), .O(n7798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3743_6_lut (.I0(GND_net), .I1(n8224[3]), .I2(n384), .I3(n30348), 
            .O(n8205[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_2_lut (.I0(GND_net), .I1(n32_adj_3603), .I2(n101_adj_3600), 
            .I3(GND_net), .O(n7962[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_6 (.CI(n30348), .I0(n8224[3]), .I1(n384), .CO(n30349));
    SB_LUT4 add_3743_5_lut (.I0(GND_net), .I1(n8224[2]), .I2(n311), .I3(n30347), 
            .O(n8205[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_2 (.CI(GND_net), .I0(n32_adj_3603), .I1(n101_adj_3600), 
            .CO(n30147));
    SB_CARRY add_3743_5 (.CI(n30347), .I0(n8224[2]), .I1(n311), .CO(n30348));
    SB_LUT4 add_3723_16_lut (.I0(GND_net), .I1(n7962[13]), .I2(GND_net), 
            .I3(n30146), .O(n7945[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_14 (.CI(n29684), .I0(n7822[11]), .I1(GND_net), .CO(n29685));
    SB_LUT4 add_3743_4_lut (.I0(GND_net), .I1(n8224[1]), .I2(n238), .I3(n30346), 
            .O(n8205[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_15_lut (.I0(GND_net), .I1(n7962[12]), .I2(GND_net), 
            .I3(n30145), .O(n7945[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_15 (.CI(n30145), .I0(n7962[12]), .I1(GND_net), .CO(n30146));
    SB_CARRY add_3743_4 (.CI(n30346), .I0(n8224[1]), .I1(n238), .CO(n30347));
    SB_LUT4 add_3723_14_lut (.I0(GND_net), .I1(n7962[11]), .I2(GND_net), 
            .I3(n30144), .O(n7945[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3716_13_lut (.I0(GND_net), .I1(n7822[10]), .I2(GND_net), 
            .I3(n29683), .O(n7798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_10 (.CI(n28557), .I0(n3054[8]), .I1(n3079[8]), .CO(n28558));
    SB_LUT4 add_3743_3_lut (.I0(GND_net), .I1(n8224[0]), .I2(n165_adj_3598), 
            .I3(n30345), .O(n8205[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_14 (.CI(n30144), .I0(n7962[11]), .I1(GND_net), .CO(n30145));
    SB_CARRY add_3743_3 (.CI(n30345), .I0(n8224[0]), .I1(n165_adj_3598), 
            .CO(n30346));
    SB_LUT4 add_3743_2_lut (.I0(GND_net), .I1(n23_adj_3597), .I2(n92), 
            .I3(GND_net), .O(n8205[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_2 (.CI(GND_net), .I0(n23_adj_3597), .I1(n92), .CO(n30345));
    SB_LUT4 add_3742_19_lut (.I0(GND_net), .I1(n8205[16]), .I2(GND_net), 
            .I3(n30344), .O(n8185[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3742_18_lut (.I0(GND_net), .I1(n8205[15]), .I2(GND_net), 
            .I3(n30343), .O(n8185[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_18 (.CI(n30343), .I0(n8205[15]), .I1(GND_net), .CO(n30344));
    SB_LUT4 add_3742_17_lut (.I0(GND_net), .I1(n8205[14]), .I2(GND_net), 
            .I3(n30342), .O(n8185[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_17 (.CI(n30342), .I0(n8205[14]), .I1(GND_net), .CO(n30343));
    SB_LUT4 add_3742_16_lut (.I0(GND_net), .I1(n8205[13]), .I2(GND_net), 
            .I3(n30341), .O(n8185[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_13_lut (.I0(GND_net), .I1(n7962[10]), .I2(GND_net), 
            .I3(n30143), .O(n7945[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_16 (.CI(n30341), .I0(n8205[13]), .I1(GND_net), .CO(n30342));
    SB_LUT4 add_3742_15_lut (.I0(GND_net), .I1(n8205[12]), .I2(GND_net), 
            .I3(n30340), .O(n8185[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_15 (.CI(n30340), .I0(n8205[12]), .I1(GND_net), .CO(n30341));
    SB_CARRY add_3723_13 (.CI(n30143), .I0(n7962[10]), .I1(GND_net), .CO(n30144));
    SB_LUT4 add_3742_14_lut (.I0(GND_net), .I1(n8205[11]), .I2(GND_net), 
            .I3(n30339), .O(n8185[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_14 (.CI(n30339), .I0(n8205[11]), .I1(GND_net), .CO(n30340));
    SB_LUT4 add_3742_13_lut (.I0(GND_net), .I1(n8205[10]), .I2(GND_net), 
            .I3(n30338), .O(n8185[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_12_lut (.I0(GND_net), .I1(n7962[9]), .I2(GND_net), 
            .I3(n30142), .O(n7945[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_13 (.CI(n30338), .I0(n8205[10]), .I1(GND_net), .CO(n30339));
    SB_CARRY add_3723_12 (.CI(n30142), .I0(n7962[9]), .I1(GND_net), .CO(n30143));
    SB_LUT4 add_3742_12_lut (.I0(GND_net), .I1(n8205[9]), .I2(GND_net), 
            .I3(n30337), .O(n8185[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_13 (.CI(n29683), .I0(n7822[10]), .I1(GND_net), .CO(n29684));
    SB_CARRY add_3742_12 (.CI(n30337), .I0(n8205[9]), .I1(GND_net), .CO(n30338));
    SB_LUT4 add_3716_12_lut (.I0(GND_net), .I1(n7822[9]), .I2(GND_net), 
            .I3(n29682), .O(n7798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_11_lut (.I0(GND_net), .I1(n7962[8]), .I2(GND_net), 
            .I3(n30141), .O(n7945[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3742_11_lut (.I0(GND_net), .I1(n8205[8]), .I2(GND_net), 
            .I3(n30336), .O(n8185[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_11 (.CI(n30336), .I0(n8205[8]), .I1(GND_net), .CO(n30337));
    SB_LUT4 add_3742_10_lut (.I0(GND_net), .I1(n8205[7]), .I2(GND_net), 
            .I3(n30335), .O(n8185[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_9_lut (.I0(GND_net), .I1(n3054[7]), .I2(n3079[7]), 
            .I3(n28556), .O(duty_23__N_3478[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_9 (.CI(n28556), .I0(n3054[7]), .I1(n3079[7]), .CO(n28557));
    SB_CARRY add_3742_10 (.CI(n30335), .I0(n8205[7]), .I1(GND_net), .CO(n30336));
    SB_CARRY add_3723_11 (.CI(n30141), .I0(n7962[8]), .I1(GND_net), .CO(n30142));
    SB_LUT4 add_3742_9_lut (.I0(GND_net), .I1(n8205[6]), .I2(GND_net), 
            .I3(n30334), .O(n8185[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_10_lut (.I0(GND_net), .I1(n7962[7]), .I2(GND_net), 
            .I3(n30140), .O(n7945[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_9 (.CI(n30334), .I0(n8205[6]), .I1(GND_net), .CO(n30335));
    SB_CARRY add_3723_10 (.CI(n30140), .I0(n7962[7]), .I1(GND_net), .CO(n30141));
    SB_LUT4 add_3723_9_lut (.I0(GND_net), .I1(n7962[6]), .I2(GND_net), 
            .I3(n30139), .O(n7945[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_12 (.CI(n29682), .I0(n7822[9]), .I1(GND_net), .CO(n29683));
    SB_LUT4 add_3716_11_lut (.I0(GND_net), .I1(n7822[8]), .I2(GND_net), 
            .I3(n29681), .O(n7798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_9 (.CI(n30139), .I0(n7962[6]), .I1(GND_net), .CO(n30140));
    SB_LUT4 add_3742_8_lut (.I0(GND_net), .I1(n8205[5]), .I2(n527), .I3(n30333), 
            .O(n8185[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_8 (.CI(n30333), .I0(n8205[5]), .I1(n527), .CO(n30334));
    SB_LUT4 add_3742_7_lut (.I0(GND_net), .I1(n8205[4]), .I2(n454), .I3(n30332), 
            .O(n8185[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_7 (.CI(n30332), .I0(n8205[4]), .I1(n454), .CO(n30333));
    SB_CARRY add_3716_11 (.CI(n29681), .I0(n7822[8]), .I1(GND_net), .CO(n29682));
    SB_LUT4 add_3742_6_lut (.I0(GND_net), .I1(n8205[3]), .I2(n381), .I3(n30331), 
            .O(n8185[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_8_lut (.I0(GND_net), .I1(n7962[5]), .I2(n536_adj_3588), 
            .I3(n30138), .O(n7945[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_6 (.CI(n30331), .I0(n8205[3]), .I1(n381), .CO(n30332));
    SB_LUT4 add_3742_5_lut (.I0(GND_net), .I1(n8205[2]), .I2(n308), .I3(n30330), 
            .O(n8185[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_8_lut (.I0(GND_net), .I1(n3054[6]), .I2(n3079[6]), 
            .I3(n28555), .O(duty_23__N_3478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34710_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n41563));
    defparam i34710_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3723_8 (.CI(n30138), .I0(n7962[5]), .I1(n536_adj_3588), 
            .CO(n30139));
    SB_LUT4 add_3716_10_lut (.I0(GND_net), .I1(n7822[7]), .I2(GND_net), 
            .I3(n29680), .O(n7798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_7_lut (.I0(GND_net), .I1(n7962[4]), .I2(n463_adj_3584), 
            .I3(n30137), .O(n7945[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_10 (.CI(n29680), .I0(n7822[7]), .I1(GND_net), .CO(n29681));
    SB_CARRY add_3723_7 (.CI(n30137), .I0(n7962[4]), .I1(n463_adj_3584), 
            .CO(n30138));
    SB_LUT4 add_3716_9_lut (.I0(GND_net), .I1(n7822[6]), .I2(GND_net), 
            .I3(n29679), .O(n7798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_6_lut (.I0(GND_net), .I1(n7962[3]), .I2(n390_adj_3583), 
            .I3(n30136), .O(n7945[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_5 (.CI(n30330), .I0(n8205[2]), .I1(n308), .CO(n30331));
    SB_CARRY add_3723_6 (.CI(n30136), .I0(n7962[3]), .I1(n390_adj_3583), 
            .CO(n30137));
    SB_LUT4 add_3723_5_lut (.I0(GND_net), .I1(n7962[2]), .I2(n317_adj_3582), 
            .I3(n30135), .O(n7945[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_9 (.CI(n29679), .I0(n7822[6]), .I1(GND_net), .CO(n29680));
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256), 
            .I3(GND_net), .O(n3079[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3716_8_lut (.I0(GND_net), .I1(n7822[5]), .I2(n515), .I3(n29678), 
            .O(n7798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_8 (.CI(n29678), .I0(n7822[5]), .I1(n515), .CO(n29679));
    SB_LUT4 add_3742_4_lut (.I0(GND_net), .I1(n8205[1]), .I2(n235), .I3(n30329), 
            .O(n8185[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_5 (.CI(n30135), .I0(n7962[2]), .I1(n317_adj_3582), 
            .CO(n30136));
    SB_LUT4 add_3716_7_lut (.I0(GND_net), .I1(n7822[4]), .I2(n442), .I3(n29677), 
            .O(n7798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_7 (.CI(n29677), .I0(n7822[4]), .I1(n442), .CO(n29678));
    SB_LUT4 add_3716_6_lut (.I0(GND_net), .I1(n7822[3]), .I2(n369), .I3(n29676), 
            .O(n7798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_4_lut (.I0(GND_net), .I1(n7962[1]), .I2(n244_adj_3672), 
            .I3(n30134), .O(n7945[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_6 (.CI(n29676), .I0(n7822[3]), .I1(n369), .CO(n29677));
    SB_LUT4 add_3716_5_lut (.I0(GND_net), .I1(n7822[2]), .I2(n296), .I3(n29675), 
            .O(n7798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_4 (.CI(n30329), .I0(n8205[1]), .I1(n235), .CO(n30330));
    SB_CARRY add_3723_4 (.CI(n30134), .I0(n7962[1]), .I1(n244_adj_3672), 
            .CO(n30135));
    SB_LUT4 add_3742_3_lut (.I0(GND_net), .I1(n8205[0]), .I2(n162), .I3(n30328), 
            .O(n8185[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_3 (.CI(n30328), .I0(n8205[0]), .I1(n162), .CO(n30329));
    SB_LUT4 add_3742_2_lut (.I0(GND_net), .I1(n20_adj_3673), .I2(n89), 
            .I3(GND_net), .O(n8185[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_2 (.CI(GND_net), .I0(n20_adj_3673), .I1(n89), .CO(n30328));
    SB_LUT4 add_3741_20_lut (.I0(GND_net), .I1(n8185[17]), .I2(GND_net), 
            .I3(n30327), .O(n8164[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_19_lut (.I0(GND_net), .I1(n8185[16]), .I2(GND_net), 
            .I3(n30326), .O(n8164[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_19 (.CI(n30326), .I0(n8185[16]), .I1(GND_net), .CO(n30327));
    SB_LUT4 add_3741_18_lut (.I0(GND_net), .I1(n8185[15]), .I2(GND_net), 
            .I3(n30325), .O(n8164[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_5 (.CI(n29675), .I0(n7822[2]), .I1(n296), .CO(n29676));
    SB_LUT4 add_3723_3_lut (.I0(GND_net), .I1(n7962[0]), .I2(n171_adj_3674), 
            .I3(n30133), .O(n7945[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_4_lut (.I0(GND_net), .I1(n7822[1]), .I2(n223), .I3(n29674), 
            .O(n7798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_4 (.CI(n29674), .I0(n7822[1]), .I1(n223), .CO(n29675));
    SB_CARRY add_3723_3 (.CI(n30133), .I0(n7962[0]), .I1(n171_adj_3674), 
            .CO(n30134));
    SB_LUT4 mux_652_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256), 
            .I3(GND_net), .O(n3079[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3573));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_654_8 (.CI(n28555), .I0(n3054[6]), .I1(n3079[6]), .CO(n28556));
    SB_CARRY add_3741_18 (.CI(n30325), .I0(n8185[15]), .I1(GND_net), .CO(n30326));
    SB_LUT4 add_3741_17_lut (.I0(GND_net), .I1(n8185[14]), .I2(GND_net), 
            .I3(n30324), .O(n8164[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_2_lut (.I0(GND_net), .I1(n29_adj_3675), .I2(n98_adj_3676), 
            .I3(GND_net), .O(n7945[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_3_lut (.I0(GND_net), .I1(n7822[0]), .I2(n150), .I3(n29673), 
            .O(n7798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_7_lut (.I0(GND_net), .I1(n3054[5]), .I2(n3079[5]), 
            .I3(n28554), .O(duty_23__N_3478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3716_3 (.CI(n29673), .I0(n7822[0]), .I1(n150), .CO(n29674));
    SB_CARRY add_3741_17 (.CI(n30324), .I0(n8185[14]), .I1(GND_net), .CO(n30325));
    SB_LUT4 add_3716_2_lut (.I0(GND_net), .I1(n8_adj_3677), .I2(n77), 
            .I3(GND_net), .O(n7798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_2 (.CI(GND_net), .I0(n8_adj_3677), .I1(n77), .CO(n29673));
    SB_CARRY add_3723_2 (.CI(GND_net), .I0(n29_adj_3675), .I1(n98_adj_3676), 
            .CO(n30133));
    SB_LUT4 add_3741_16_lut (.I0(GND_net), .I1(n8185[13]), .I2(GND_net), 
            .I3(n30323), .O(n8164[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_17_lut (.I0(GND_net), .I1(n7945[14]), .I2(GND_net), 
            .I3(n30132), .O(n7927[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_16_lut (.I0(GND_net), .I1(n7945[13]), .I2(GND_net), 
            .I3(n30131), .O(n7927[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_16 (.CI(n30131), .I0(n7945[13]), .I1(GND_net), .CO(n30132));
    SB_LUT4 add_3722_15_lut (.I0(GND_net), .I1(n7945[12]), .I2(GND_net), 
            .I3(n30130), .O(n7927[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_7 (.CI(n28554), .I0(n3054[5]), .I1(n3079[5]), .CO(n28555));
    SB_CARRY add_3741_16 (.CI(n30323), .I0(n8185[13]), .I1(GND_net), .CO(n30324));
    SB_LUT4 add_3741_15_lut (.I0(GND_net), .I1(n8185[12]), .I2(GND_net), 
            .I3(n30322), .O(n8164[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_15 (.CI(n30322), .I0(n8185[12]), .I1(GND_net), .CO(n30323));
    SB_CARRY add_3722_15 (.CI(n30130), .I0(n7945[12]), .I1(GND_net), .CO(n30131));
    SB_LUT4 add_654_6_lut (.I0(GND_net), .I1(n3054[4]), .I2(n3079[4]), 
            .I3(n28553), .O(duty_23__N_3478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_14_lut (.I0(GND_net), .I1(n8185[11]), .I2(GND_net), 
            .I3(n30321), .O(n8164[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_14_lut (.I0(GND_net), .I1(n7945[11]), .I2(GND_net), 
            .I3(n30129), .O(n7927[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_14 (.CI(n30321), .I0(n8185[11]), .I1(GND_net), .CO(n30322));
    SB_CARRY add_654_6 (.CI(n28553), .I0(n3054[4]), .I1(n3079[4]), .CO(n28554));
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3741_13_lut (.I0(GND_net), .I1(n8185[10]), .I2(GND_net), 
            .I3(n30320), .O(n8164[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_13 (.CI(n30320), .I0(n8185[10]), .I1(GND_net), .CO(n30321));
    SB_CARRY add_3722_14 (.CI(n30129), .I0(n7945[11]), .I1(GND_net), .CO(n30130));
    SB_LUT4 add_3722_13_lut (.I0(GND_net), .I1(n7945[10]), .I2(GND_net), 
            .I3(n30128), .O(n7927[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_12_lut (.I0(GND_net), .I1(n8185[9]), .I2(GND_net), 
            .I3(n30319), .O(n8164[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_12 (.CI(n30319), .I0(n8185[9]), .I1(GND_net), .CO(n30320));
    SB_LUT4 add_3741_11_lut (.I0(GND_net), .I1(n8185[8]), .I2(GND_net), 
            .I3(n30318), .O(n8164[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_11 (.CI(n30318), .I0(n8185[8]), .I1(GND_net), .CO(n30319));
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_3678));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_3679));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_654_5_lut (.I0(GND_net), .I1(n3054[3]), .I2(n3079[3]), 
            .I3(n28552), .O(duty_23__N_3478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_10_lut (.I0(GND_net), .I1(n8185[7]), .I2(GND_net), 
            .I3(n30317), .O(n8164[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_3680));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34542_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n41395));
    defparam i34542_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i34532_3_lut (.I0(n11_adj_3680), .I1(n9_adj_3679), .I2(n41395), 
            .I3(GND_net), .O(n41385));
    defparam i34532_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mux_652_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256), 
            .I3(GND_net), .O(n3079[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_654_5 (.CI(n28552), .I0(n3054[3]), .I1(n3079[3]), .CO(n28553));
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_420_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n45150));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_420_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35797_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n45150), 
            .I2(IntegralLimit[7]), .I3(n41385), .O(n42651));
    defparam i35797_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_3741_10 (.CI(n30317), .I0(n8185[7]), .I1(GND_net), .CO(n30318));
    SB_CARRY add_3722_13 (.CI(n30128), .I0(n7945[10]), .I1(GND_net), .CO(n30129));
    SB_LUT4 i35781_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3678), 
            .I2(IntegralLimit[9]), .I3(n42651), .O(n42635));
    defparam i35781_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_402_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n45132));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_402_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35779_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3678), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3679), .O(n42633));
    defparam i35779_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_3666));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35771_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n45132), 
            .I2(IntegralLimit[11]), .I3(n42633), .O(n42625));
    defparam i35771_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_3741_9_lut (.I0(GND_net), .I1(n8185[6]), .I2(GND_net), 
            .I3(n30316), .O(n8164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_396_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n45126));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_396_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3722_12_lut (.I0(GND_net), .I1(n7945[9]), .I2(GND_net), 
            .I3(n30127), .O(n7927[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_9 (.CI(n30316), .I0(n8185[6]), .I1(GND_net), .CO(n30317));
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3573), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3561));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3722_12 (.CI(n30127), .I0(n7945[9]), .I1(GND_net), .CO(n30128));
    SB_LUT4 add_3722_11_lut (.I0(GND_net), .I1(n7945[8]), .I2(GND_net), 
            .I3(n30126), .O(n7927[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35000_4_lut (.I0(n27_adj_3594), .I1(n15_adj_3632), .I2(n13_adj_3633), 
            .I3(n11_adj_3635), .O(n41854));
    defparam i35000_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3665));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35014_4_lut (.I0(n21_adj_3608), .I1(n19_adj_3627), .I2(n17_adj_3628), 
            .I3(n9_adj_3641), .O(n41868));
    defparam i35014_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_3681), .I3(GND_net), 
            .O(n16_adj_3682));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_DFFE \PID_CONTROLLER.integral_1202__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[0]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 i34946_2_lut (.I0(n43_adj_3681), .I1(n19_adj_3627), .I2(GND_net), 
            .I3(GND_net), .O(n41800));
    defparam i34946_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3628), .I3(GND_net), 
            .O(n8_adj_3683));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mux_652_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256), 
            .I3(GND_net), .O(n3079[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_3682), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_3684), .I3(GND_net), 
            .O(n24_adj_3685));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35035_2_lut (.I0(n7_adj_3646), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n41889));
    defparam i35035_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_3741_8_lut (.I0(GND_net), .I1(n8185[5]), .I2(n524), .I3(n30315), 
            .O(n8164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3664));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35675_4_lut (.I0(n13_adj_3633), .I1(n11_adj_3635), .I2(n9_adj_3641), 
            .I3(n41889), .O(n42529));
    defparam i35675_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35667_4_lut (.I0(n19_adj_3627), .I1(n17_adj_3628), .I2(n15_adj_3632), 
            .I3(n42529), .O(n42521));
    defparam i35667_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36410_4_lut (.I0(n25_adj_3599), .I1(n23_adj_3606), .I2(n21_adj_3608), 
            .I3(n42521), .O(n43264));
    defparam i36410_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3741_8 (.CI(n30315), .I0(n8185[5]), .I1(n524), .CO(n30316));
    SB_LUT4 i35978_4_lut (.I0(n31_adj_3568), .I1(n29_adj_3592), .I2(n27_adj_3594), 
            .I3(n43264), .O(n42832));
    defparam i35978_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36514_4_lut (.I0(n37), .I1(n35_adj_3566), .I2(n33), .I3(n42832), 
            .O(n43368));
    defparam i36514_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35201_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n45150), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3680), .O(n42055));
    defparam i35201_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_389_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n45119));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_389_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3741_7_lut (.I0(GND_net), .I1(n8185[4]), .I2(n451), .I3(n30314), 
            .O(n8164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35749_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n45119), 
            .I2(IntegralLimit[14]), .I3(n42055), .O(n42603));
    defparam i35749_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_384_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n45114));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_384_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3722_11 (.CI(n30126), .I0(n7945[8]), .I1(GND_net), .CO(n30127));
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_3686));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35094_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n41948));
    defparam i35094_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_407_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n45137));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_407_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3722_10_lut (.I0(GND_net), .I1(n7945[7]), .I2(GND_net), 
            .I3(n30125), .O(n7927[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3687));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_3686), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_3688));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3722_10 (.CI(n30125), .I0(n7945[7]), .I1(GND_net), .CO(n30126));
    SB_CARRY add_3741_7 (.CI(n30314), .I0(n8185[4]), .I1(n451), .CO(n30315));
    SB_LUT4 i36259_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n45132), 
            .I2(IntegralLimit[11]), .I3(n42635), .O(n43113));
    defparam i36259_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_3722_9_lut (.I0(GND_net), .I1(n7945[6]), .I2(GND_net), 
            .I3(n30124), .O(n7927[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3660));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35128_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n45126), 
            .I2(IntegralLimit[13]), .I3(n43113), .O(n41982));
    defparam i35128_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_387_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n45117));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_387_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36026_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n45117), 
            .I2(IntegralLimit[15]), .I3(n41982), .O(n42880));
    defparam i36026_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_413_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n45143));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_413_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36422_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n45143), 
            .I2(IntegralLimit[17]), .I3(n42880), .O(n43276));
    defparam i36422_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_378_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n45108));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_378_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36592_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n45108), 
            .I2(IntegralLimit[19]), .I3(n43276), .O(n43446));
    defparam i36592_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_375_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n45105));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3689));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3741_6_lut (.I0(GND_net), .I1(n8185[3]), .I2(n378), .I3(n30313), 
            .O(n8164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35041_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n41895));
    defparam i35041_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3689), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3690));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3691));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36211_3_lut (.I0(n6_adj_3691), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n43065));   // verilog/motorControl.v(39[10:34])
    defparam i36211_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36212_3_lut (.I0(n43065), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n43066));   // verilog/motorControl.v(39[10:34])
    defparam i36212_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3741_6 (.CI(n30313), .I0(n8185[3]), .I1(n378), .CO(n30314));
    SB_LUT4 i35045_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n45126), 
            .I2(IntegralLimit[21]), .I3(n42625), .O(n41899));
    defparam i35045_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i36074_4_lut (.I0(n24_adj_3690), .I1(n8_adj_3692), .I2(n45103), 
            .I3(n41895), .O(n42928));   // verilog/motorControl.v(39[10:34])
    defparam i36074_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35318_3_lut (.I0(n43066), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n42172));   // verilog/motorControl.v(39[10:34])
    defparam i35318_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256), 
            .I3(GND_net), .O(n3079[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3454 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_3693));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i36199_3_lut (.I0(n4_adj_3693), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_3594), .I3(GND_net), .O(n43053));   // verilog/motorControl.v(39[38:63])
    defparam i36199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36200_3_lut (.I0(n43053), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_3592), .I3(GND_net), .O(n43054));   // verilog/motorControl.v(39[38:63])
    defparam i36200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_3694));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34976_2_lut (.I0(n33), .I1(n15_adj_3632), .I2(GND_net), .I3(GND_net), 
            .O(n41830));
    defparam i34976_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3633), .I3(GND_net), 
            .O(n10_adj_3695));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3694), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_3566), .I3(GND_net), 
            .O(n30_adj_3696));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34980_4_lut (.I0(n33), .I1(n31_adj_3568), .I2(n29_adj_3592), 
            .I3(n41854), .O(n41834));
    defparam i34980_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36432_4_lut (.I0(n30_adj_3696), .I1(n10_adj_3695), .I2(n35_adj_3566), 
            .I3(n41830), .O(n43286));   // verilog/motorControl.v(39[38:63])
    defparam i36432_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35330_3_lut (.I0(n43054), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_3568), .I3(GND_net), .O(n42184));   // verilog/motorControl.v(39[38:63])
    defparam i35330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36570_4_lut (.I0(n42184), .I1(n43286), .I2(n35_adj_3566), 
            .I3(n41834), .O(n43424));   // verilog/motorControl.v(39[38:63])
    defparam i36570_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36571_3_lut (.I0(n43424), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n43425));   // verilog/motorControl.v(39[38:63])
    defparam i36571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36563_3_lut (.I0(n43425), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n43417));   // verilog/motorControl.v(39[38:63])
    defparam i36563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_3646), .I3(GND_net), 
            .O(n6_adj_3697));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36201_3_lut (.I0(n6_adj_3697), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_3608), .I3(GND_net), .O(n43055));   // verilog/motorControl.v(39[38:63])
    defparam i36201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3659));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36202_3_lut (.I0(n43055), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_3606), .I3(GND_net), .O(n43056));   // verilog/motorControl.v(39[38:63])
    defparam i36202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3658));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34954_4_lut (.I0(n43_adj_3681), .I1(n25_adj_3599), .I2(n23_adj_3606), 
            .I3(n41868), .O(n41808));
    defparam i34954_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36076_4_lut (.I0(n24_adj_3685), .I1(n8_adj_3683), .I2(n45_adj_3684), 
            .I3(n41800), .O(n42930));   // verilog/motorControl.v(39[38:63])
    defparam i36076_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35328_3_lut (.I0(n43056), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_3599), .I3(GND_net), .O(n42182));   // verilog/motorControl.v(39[38:63])
    defparam i35328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_3657));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_654_4_lut (.I0(GND_net), .I1(n3054[2]), .I2(n3079[2]), 
            .I3(n28551), .O(duty_23__N_3478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_4 (.CI(n28551), .I0(n3054[2]), .I1(n3079[2]), .CO(n28552));
    SB_CARRY add_3722_9 (.CI(n30124), .I0(n7945[6]), .I1(GND_net), .CO(n30125));
    SB_LUT4 add_3741_5_lut (.I0(GND_net), .I1(n8185[2]), .I2(n305), .I3(n30312), 
            .O(n8164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34958_4_lut (.I0(n43_adj_3681), .I1(n41_adj_3698), .I2(n39), 
            .I3(n43368), .O(n41812));
    defparam i34958_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36485_4_lut (.I0(n42182), .I1(n42930), .I2(n45_adj_3684), 
            .I3(n41808), .O(n43339));   // verilog/motorControl.v(39[38:63])
    defparam i36485_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35336_3_lut (.I0(n43417), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_3698), .I3(GND_net), .O(n42190));   // verilog/motorControl.v(39[38:63])
    defparam i35336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_3656));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3741_5 (.CI(n30312), .I0(n8185[2]), .I1(n305), .CO(n30313));
    SB_LUT4 i36487_4_lut (.I0(n42190), .I1(n43339), .I2(n45_adj_3684), 
            .I3(n41812), .O(n43341));   // verilog/motorControl.v(39[38:63])
    defparam i36487_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3699));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36207_3_lut (.I0(n4_adj_3699), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n43061));   // verilog/motorControl.v(39[10:34])
    defparam i36207_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36208_3_lut (.I0(n43061), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n43062));   // verilog/motorControl.v(39[10:34])
    defparam i36208_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35110_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n45114), 
            .I2(IntegralLimit[16]), .I3(n42603), .O(n41964));
    defparam i35110_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i36430_4_lut (.I0(n30_adj_3688), .I1(n10_adj_3687), .I2(n45137), 
            .I3(n41948), .O(n43284));   // verilog/motorControl.v(39[10:34])
    defparam i36430_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35320_3_lut (.I0(n43062), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n42174));   // verilog/motorControl.v(39[10:34])
    defparam i35320_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3741_4_lut (.I0(GND_net), .I1(n8185[1]), .I2(n232), .I3(n30311), 
            .O(n8164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36568_4_lut (.I0(n42174), .I1(n43284), .I2(n45137), .I3(n41964), 
            .O(n43422));   // verilog/motorControl.v(39[10:34])
    defparam i36568_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36569_3_lut (.I0(n43422), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n43423));   // verilog/motorControl.v(39[10:34])
    defparam i36569_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36565_3_lut (.I0(n43423), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n43419));   // verilog/motorControl.v(39[10:34])
    defparam i36565_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35047_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n45105), 
            .I2(IntegralLimit[21]), .I3(n43446), .O(n41901));
    defparam i35047_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_373_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n45103));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_373_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36481_4_lut (.I0(n42172), .I1(n42928), .I2(n45103), .I3(n41899), 
            .O(n43335));   // verilog/motorControl.v(39[10:34])
    defparam i36481_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35326_3_lut (.I0(n43419), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n42180));   // verilog/motorControl.v(39[10:34])
    defparam i35326_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36488_3_lut (.I0(n43341), .I1(\PID_CONTROLLER.integral_23__N_3454 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3453 ));   // verilog/motorControl.v(39[38:63])
    defparam i36488_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3722_8_lut (.I0(GND_net), .I1(n7945[5]), .I2(n533_adj_3671), 
            .I3(n30123), .O(n7927[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36483_4_lut (.I0(n42180), .I1(n43335), .I2(n45103), .I3(n41901), 
            .O(n43337));   // verilog/motorControl.v(39[10:34])
    defparam i36483_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3722_8 (.CI(n30123), .I0(n7945[5]), .I1(n533_adj_3671), 
            .CO(n30124));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_838_4_lut  (.I0(n43337), .I1(\PID_CONTROLLER.integral_23__N_3453 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3451 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_838_4_lut .LUT_INIT = 16'h80c8;
    SB_CARRY add_3741_4 (.CI(n30311), .I0(n8185[1]), .I1(n232), .CO(n30312));
    SB_LUT4 add_3741_3_lut (.I0(GND_net), .I1(n8185[0]), .I2(n159), .I3(n30310), 
            .O(n8164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_7_lut (.I0(GND_net), .I1(n7945[4]), .I2(n460_adj_3670), 
            .I3(n30122), .O(n7927[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_7 (.CI(n30122), .I0(n7945[4]), .I1(n460_adj_3670), 
            .CO(n30123));
    SB_LUT4 mux_652_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256), 
            .I3(GND_net), .O(n3079[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3741_3 (.CI(n30310), .I0(n8185[0]), .I1(n159), .CO(n30311));
    SB_LUT4 add_3722_6_lut (.I0(GND_net), .I1(n7945[3]), .I2(n387_adj_3663), 
            .I3(n30121), .O(n7927[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_2_lut (.I0(GND_net), .I1(n17_adj_3662), .I2(n86), 
            .I3(GND_net), .O(n8164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_6 (.CI(n30121), .I0(n7945[3]), .I1(n387_adj_3663), 
            .CO(n30122));
    SB_CARRY add_3741_2 (.CI(GND_net), .I0(n17_adj_3662), .I1(n86), .CO(n30310));
    SB_LUT4 add_3722_5_lut (.I0(GND_net), .I1(n7945[2]), .I2(n314_adj_3661), 
            .I3(n30120), .O(n7927[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_21_lut (.I0(GND_net), .I1(n8164[18]), .I2(GND_net), 
            .I3(n30309), .O(n8142[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_5 (.CI(n30120), .I0(n7945[2]), .I1(n314_adj_3661), 
            .CO(n30121));
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_3655));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37372_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n44224));   // verilog/motorControl.v(37[14] 56[8])
    defparam i37372_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_3654));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_3653));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_3652));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_652_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256), 
            .I3(GND_net), .O(n3079[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_652_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256), 
            .I3(GND_net), .O(n3079[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3740_20_lut (.I0(GND_net), .I1(n8164[17]), .I2(GND_net), 
            .I3(n30308), .O(n8142[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_4_lut (.I0(GND_net), .I1(n7945[1]), .I2(n241), .I3(n30119), 
            .O(n7927[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_20 (.CI(n30308), .I0(n8164[17]), .I1(GND_net), .CO(n30309));
    SB_CARRY add_3722_4 (.CI(n30119), .I0(n7945[1]), .I1(n241), .CO(n30120));
    SB_LUT4 add_3722_3_lut (.I0(GND_net), .I1(n7945[0]), .I2(n168), .I3(n30118), 
            .O(n7927[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_19_lut (.I0(GND_net), .I1(n8164[16]), .I2(GND_net), 
            .I3(n30307), .O(n8142[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_3 (.CI(n30118), .I0(n7945[0]), .I1(n168), .CO(n30119));
    SB_CARRY add_3740_19 (.CI(n30307), .I0(n8164[16]), .I1(GND_net), .CO(n30308));
    SB_LUT4 add_3722_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7927[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_18_lut (.I0(GND_net), .I1(n8164[15]), .I2(GND_net), 
            .I3(n30306), .O(n8142[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n30118));
    SB_LUT4 add_654_3_lut (.I0(GND_net), .I1(n3054[1]), .I2(n3079[1]), 
            .I3(n28550), .O(duty_23__N_3478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_654_3 (.CI(n28550), .I0(n3054[1]), .I1(n3079[1]), .CO(n28551));
    SB_CARRY add_3740_18 (.CI(n30306), .I0(n8164[15]), .I1(GND_net), .CO(n30307));
    SB_LUT4 add_3721_18_lut (.I0(GND_net), .I1(n7927[15]), .I2(GND_net), 
            .I3(n30117), .O(n7908[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_17_lut (.I0(GND_net), .I1(n7927[14]), .I2(GND_net), 
            .I3(n30116), .O(n7908[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_17_lut (.I0(GND_net), .I1(n8164[14]), .I2(GND_net), 
            .I3(n30305), .O(n8142[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_17 (.CI(n30305), .I0(n8164[14]), .I1(GND_net), .CO(n30306));
    SB_CARRY add_3721_17 (.CI(n30116), .I0(n7927[14]), .I1(GND_net), .CO(n30117));
    SB_LUT4 add_3740_16_lut (.I0(GND_net), .I1(n8164[13]), .I2(GND_net), 
            .I3(n30304), .O(n8142[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_16_lut (.I0(GND_net), .I1(n7927[13]), .I2(GND_net), 
            .I3(n30115), .O(n7908[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_16 (.CI(n30304), .I0(n8164[13]), .I1(GND_net), .CO(n30305));
    SB_CARRY add_3721_16 (.CI(n30115), .I0(n7927[13]), .I1(GND_net), .CO(n30116));
    SB_LUT4 add_3740_15_lut (.I0(GND_net), .I1(n8164[12]), .I2(GND_net), 
            .I3(n30303), .O(n8142[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_15_lut (.I0(GND_net), .I1(n7927[12]), .I2(GND_net), 
            .I3(n30114), .O(n7908[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_15 (.CI(n30114), .I0(n7927[12]), .I1(GND_net), .CO(n30115));
    SB_CARRY add_3740_15 (.CI(n30303), .I0(n8164[12]), .I1(GND_net), .CO(n30304));
    SB_LUT4 add_3721_14_lut (.I0(GND_net), .I1(n7927[11]), .I2(GND_net), 
            .I3(n30113), .O(n7908[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_14 (.CI(n30113), .I0(n7927[11]), .I1(GND_net), .CO(n30114));
    SB_LUT4 add_3740_14_lut (.I0(GND_net), .I1(n8164[11]), .I2(GND_net), 
            .I3(n30302), .O(n8142[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_13_lut (.I0(GND_net), .I1(n7927[10]), .I2(GND_net), 
            .I3(n30112), .O(n7908[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_13 (.CI(n30112), .I0(n7927[10]), .I1(GND_net), .CO(n30113));
    SB_CARRY add_3740_14 (.CI(n30302), .I0(n8164[11]), .I1(GND_net), .CO(n30303));
    SB_LUT4 add_3721_12_lut (.I0(GND_net), .I1(n7927[9]), .I2(GND_net), 
            .I3(n30111), .O(n7908[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_13_lut (.I0(GND_net), .I1(n8164[10]), .I2(GND_net), 
            .I3(n30301), .O(n8142[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_654_2_lut (.I0(GND_net), .I1(n3054[0]), .I2(n3079[0]), 
            .I3(GND_net), .O(duty_23__N_3478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_12 (.CI(n30111), .I0(n7927[9]), .I1(GND_net), .CO(n30112));
    SB_CARRY add_654_2 (.CI(GND_net), .I0(n3054[0]), .I1(n3079[0]), .CO(n28550));
    SB_CARRY add_3740_13 (.CI(n30301), .I0(n8164[10]), .I1(GND_net), .CO(n30302));
    SB_LUT4 add_3721_11_lut (.I0(GND_net), .I1(n7927[8]), .I2(GND_net), 
            .I3(n30110), .O(n7908[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_12_lut (.I0(GND_net), .I1(n8164[9]), .I2(GND_net), 
            .I3(n30300), .O(n8142[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_11 (.CI(n30110), .I0(n7927[8]), .I1(GND_net), .CO(n30111));
    SB_LUT4 add_3721_10_lut (.I0(GND_net), .I1(n7927[7]), .I2(GND_net), 
            .I3(n30109), .O(n7908[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_12 (.CI(n30300), .I0(n8164[9]), .I1(GND_net), .CO(n30301));
    SB_CARRY add_3721_10 (.CI(n30109), .I0(n7927[7]), .I1(GND_net), .CO(n30110));
    SB_LUT4 add_3721_9_lut (.I0(GND_net), .I1(n7927[6]), .I2(GND_net), 
            .I3(n30108), .O(n7908[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_11_lut (.I0(GND_net), .I1(n8164[8]), .I2(GND_net), 
            .I3(n30299), .O(n8142[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_9 (.CI(n30108), .I0(n7927[6]), .I1(GND_net), .CO(n30109));
    SB_CARRY add_3740_11 (.CI(n30299), .I0(n8164[8]), .I1(GND_net), .CO(n30300));
    SB_LUT4 add_3721_8_lut (.I0(GND_net), .I1(n7927[5]), .I2(n530_adj_3649), 
            .I3(n30107), .O(n7908[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_10_lut (.I0(GND_net), .I1(n8164[7]), .I2(GND_net), 
            .I3(n30298), .O(n8142[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_8 (.CI(n30107), .I0(n7927[5]), .I1(n530_adj_3649), 
            .CO(n30108));
    SB_CARRY add_3740_10 (.CI(n30298), .I0(n8164[7]), .I1(GND_net), .CO(n30299));
    SB_LUT4 add_3721_7_lut (.I0(GND_net), .I1(n7927[4]), .I2(n457_adj_3648), 
            .I3(n30106), .O(n7908[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_9_lut (.I0(GND_net), .I1(n8164[6]), .I2(GND_net), 
            .I3(n30297), .O(n8142[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_7 (.CI(n30106), .I0(n7927[4]), .I1(n457_adj_3648), 
            .CO(n30107));
    SB_LUT4 add_3721_6_lut (.I0(GND_net), .I1(n7927[3]), .I2(n384_adj_3643), 
            .I3(n30105), .O(n7908[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_9 (.CI(n30297), .I0(n8164[6]), .I1(GND_net), .CO(n30298));
    SB_CARRY add_3721_6 (.CI(n30105), .I0(n7927[3]), .I1(n384_adj_3643), 
            .CO(n30106));
    SB_LUT4 add_3740_8_lut (.I0(GND_net), .I1(n8164[5]), .I2(n521), .I3(n30296), 
            .O(n8142[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_5_lut (.I0(GND_net), .I1(n7927[2]), .I2(n311_adj_3642), 
            .I3(n30104), .O(n7908[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_8 (.CI(n30296), .I0(n8164[5]), .I1(n521), .CO(n30297));
    SB_CARRY add_3721_5 (.CI(n30104), .I0(n7927[2]), .I1(n311_adj_3642), 
            .CO(n30105));
    SB_LUT4 add_3740_7_lut (.I0(GND_net), .I1(n8164[4]), .I2(n448), .I3(n30295), 
            .O(n8142[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_4_lut (.I0(GND_net), .I1(n7927[1]), .I2(n238_adj_3640), 
            .I3(n30103), .O(n7908[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_4 (.CI(n30103), .I0(n7927[1]), .I1(n238_adj_3640), 
            .CO(n30104));
    SB_CARRY add_3740_7 (.CI(n30295), .I0(n8164[4]), .I1(n448), .CO(n30296));
    SB_LUT4 add_3721_3_lut (.I0(GND_net), .I1(n7927[0]), .I2(n165), .I3(n30102), 
            .O(n7908[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_3 (.CI(n30102), .I0(n7927[0]), .I1(n165), .CO(n30103));
    SB_LUT4 add_3721_2_lut (.I0(GND_net), .I1(n23_adj_3701), .I2(n92_adj_3702), 
            .I3(GND_net), .O(n7908[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_6_lut (.I0(GND_net), .I1(n8164[3]), .I2(n375), .I3(n30294), 
            .O(n8142[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3355[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_3740_6 (.CI(n30294), .I0(n8164[3]), .I1(n375), .CO(n30295));
    SB_CARRY add_3721_2 (.CI(GND_net), .I0(n23_adj_3701), .I1(n92_adj_3702), 
            .CO(n30102));
    SB_LUT4 add_3720_19_lut (.I0(GND_net), .I1(n7908[16]), .I2(GND_net), 
            .I3(n30101), .O(n7888[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_5_lut (.I0(GND_net), .I1(n8164[2]), .I2(n302), .I3(n30293), 
            .O(n8142[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_5 (.CI(n30293), .I0(n8164[2]), .I1(n302), .CO(n30294));
    SB_LUT4 add_3720_18_lut (.I0(GND_net), .I1(n7908[15]), .I2(GND_net), 
            .I3(n30100), .O(n7888[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_18 (.CI(n30100), .I0(n7908[15]), .I1(GND_net), .CO(n30101));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3355[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_3740_4_lut (.I0(GND_net), .I1(n8164[1]), .I2(n229), .I3(n30292), 
            .O(n8142[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_17_lut (.I0(GND_net), .I1(n7908[14]), .I2(GND_net), 
            .I3(n30099), .O(n7888[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_4 (.CI(n30292), .I0(n8164[1]), .I1(n229), .CO(n30293));
    SB_CARRY add_3720_17 (.CI(n30099), .I0(n7908[14]), .I1(GND_net), .CO(n30100));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3355[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3355[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3355[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3355[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3355[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3355[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3355[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3355[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3355[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3355[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3355[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3355[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3355[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3355[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3355[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3355[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3355[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3355[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3355[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3355[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3355[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_3740_3_lut (.I0(GND_net), .I1(n8164[0]), .I2(n156), .I3(n30291), 
            .O(n8142[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_16_lut (.I0(GND_net), .I1(n7908[13]), .I2(GND_net), 
            .I3(n30098), .O(n7888[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_3 (.CI(n30291), .I0(n8164[0]), .I1(n156), .CO(n30292));
    SB_LUT4 add_3740_2_lut (.I0(GND_net), .I1(n14_adj_3703), .I2(n83), 
            .I3(GND_net), .O(n8142[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_16 (.CI(n30098), .I0(n7908[13]), .I1(GND_net), .CO(n30099));
    SB_CARRY add_3740_2 (.CI(GND_net), .I0(n14_adj_3703), .I1(n83), .CO(n30291));
    SB_LUT4 add_3720_15_lut (.I0(GND_net), .I1(n7908[12]), .I2(GND_net), 
            .I3(n30097), .O(n7888[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_15 (.CI(n30097), .I0(n7908[12]), .I1(GND_net), .CO(n30098));
    SB_LUT4 add_3739_22_lut (.I0(GND_net), .I1(n8142[19]), .I2(GND_net), 
            .I3(n30290), .O(n8119[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_14_lut (.I0(GND_net), .I1(n7908[11]), .I2(GND_net), 
            .I3(n30096), .O(n7888[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_21_lut (.I0(GND_net), .I1(n8142[18]), .I2(GND_net), 
            .I3(n30289), .O(n8119[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_14 (.CI(n30096), .I0(n7908[11]), .I1(GND_net), .CO(n30097));
    SB_LUT4 add_3720_13_lut (.I0(GND_net), .I1(n7908[10]), .I2(GND_net), 
            .I3(n30095), .O(n7888[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_13 (.CI(n30095), .I0(n7908[10]), .I1(GND_net), .CO(n30096));
    SB_LUT4 add_3720_12_lut (.I0(GND_net), .I1(n7908[9]), .I2(GND_net), 
            .I3(n30094), .O(n7888[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_21 (.CI(n30289), .I0(n8142[18]), .I1(GND_net), .CO(n30290));
    SB_CARRY add_3720_12 (.CI(n30094), .I0(n7908[9]), .I1(GND_net), .CO(n30095));
    SB_LUT4 add_3720_11_lut (.I0(GND_net), .I1(n7908[8]), .I2(GND_net), 
            .I3(n30093), .O(n7888[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_20_lut (.I0(GND_net), .I1(n8142[17]), .I2(GND_net), 
            .I3(n30288), .O(n8119[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_11 (.CI(n30093), .I0(n7908[8]), .I1(GND_net), .CO(n30094));
    SB_CARRY add_3739_20 (.CI(n30288), .I0(n8142[17]), .I1(GND_net), .CO(n30289));
    SB_LUT4 add_3720_10_lut (.I0(GND_net), .I1(n7908[7]), .I2(GND_net), 
            .I3(n30092), .O(n7888[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_19_lut (.I0(GND_net), .I1(n8142[16]), .I2(GND_net), 
            .I3(n30287), .O(n8119[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_10 (.CI(n30092), .I0(n7908[7]), .I1(GND_net), .CO(n30093));
    SB_LUT4 add_3720_9_lut (.I0(GND_net), .I1(n7908[6]), .I2(GND_net), 
            .I3(n30091), .O(n7888[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_19 (.CI(n30287), .I0(n8142[16]), .I1(GND_net), .CO(n30288));
    SB_CARRY add_3720_9 (.CI(n30091), .I0(n7908[6]), .I1(GND_net), .CO(n30092));
    SB_LUT4 add_3739_18_lut (.I0(GND_net), .I1(n8142[15]), .I2(GND_net), 
            .I3(n30286), .O(n8119[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_8_lut (.I0(GND_net), .I1(n7908[5]), .I2(n527_adj_3704), 
            .I3(n30090), .O(n7888[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_18 (.CI(n30286), .I0(n8142[15]), .I1(GND_net), .CO(n30287));
    SB_CARRY add_3720_8 (.CI(n30090), .I0(n7908[5]), .I1(n527_adj_3704), 
            .CO(n30091));
    SB_LUT4 add_3739_17_lut (.I0(GND_net), .I1(n8142[14]), .I2(GND_net), 
            .I3(n30285), .O(n8119[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_7_lut (.I0(GND_net), .I1(n7908[4]), .I2(n454_adj_3705), 
            .I3(n30089), .O(n7888[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_17 (.CI(n30285), .I0(n8142[14]), .I1(GND_net), .CO(n30286));
    SB_CARRY add_3720_7 (.CI(n30089), .I0(n7908[4]), .I1(n454_adj_3705), 
            .CO(n30090));
    SB_LUT4 add_3720_6_lut (.I0(GND_net), .I1(n7908[3]), .I2(n381_adj_3706), 
            .I3(n30088), .O(n7888[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_16_lut (.I0(GND_net), .I1(n8142[13]), .I2(GND_net), 
            .I3(n30284), .O(n8119[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_6 (.CI(n30088), .I0(n7908[3]), .I1(n381_adj_3706), 
            .CO(n30089));
    SB_LUT4 add_3720_5_lut (.I0(GND_net), .I1(n7908[2]), .I2(n308_adj_3707), 
            .I3(n30087), .O(n7888[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_16 (.CI(n30284), .I0(n8142[13]), .I1(GND_net), .CO(n30285));
    SB_CARRY add_3720_5 (.CI(n30087), .I0(n7908[2]), .I1(n308_adj_3707), 
            .CO(n30088));
    SB_LUT4 add_3739_15_lut (.I0(GND_net), .I1(n8142[12]), .I2(GND_net), 
            .I3(n30283), .O(n8119[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_4_lut (.I0(GND_net), .I1(n7908[1]), .I2(n235_adj_3708), 
            .I3(n30086), .O(n7888[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_15 (.CI(n30283), .I0(n8142[12]), .I1(GND_net), .CO(n30284));
    SB_CARRY add_3720_4 (.CI(n30086), .I0(n7908[1]), .I1(n235_adj_3708), 
            .CO(n30087));
    SB_LUT4 add_3739_14_lut (.I0(GND_net), .I1(n8142[11]), .I2(GND_net), 
            .I3(n30282), .O(n8119[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_14 (.CI(n30282), .I0(n8142[11]), .I1(GND_net), .CO(n30283));
    SB_LUT4 add_3720_3_lut (.I0(GND_net), .I1(n7908[0]), .I2(n162_adj_3709), 
            .I3(n30085), .O(n7888[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3754_7_lut (.I0(GND_net), .I1(n31074), .I2(n490), .I3(n30470), 
            .O(n8359[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_13_lut (.I0(GND_net), .I1(n8142[10]), .I2(GND_net), 
            .I3(n30281), .O(n8119[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_13 (.CI(n30281), .I0(n8142[10]), .I1(GND_net), .CO(n30282));
    SB_CARRY add_3720_3 (.CI(n30085), .I0(n7908[0]), .I1(n162_adj_3709), 
            .CO(n30086));
    SB_LUT4 add_3720_2_lut (.I0(GND_net), .I1(n20_adj_3710), .I2(n89_adj_3711), 
            .I3(GND_net), .O(n7888[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3754_6_lut (.I0(GND_net), .I1(n8367[3]), .I2(n417), .I3(n30469), 
            .O(n8359[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_12_lut (.I0(GND_net), .I1(n8142[9]), .I2(GND_net), 
            .I3(n30280), .O(n8119[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_2 (.CI(GND_net), .I0(n20_adj_3710), .I1(n89_adj_3711), 
            .CO(n30085));
    SB_LUT4 add_3719_20_lut (.I0(GND_net), .I1(n7888[17]), .I2(GND_net), 
            .I3(n30084), .O(n7867[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_12 (.CI(n30280), .I0(n8142[9]), .I1(GND_net), .CO(n30281));
    SB_LUT4 add_3719_19_lut (.I0(GND_net), .I1(n7888[16]), .I2(GND_net), 
            .I3(n30083), .O(n7867[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_19 (.CI(n30083), .I0(n7888[16]), .I1(GND_net), .CO(n30084));
    SB_CARRY add_3754_6 (.CI(n30469), .I0(n8367[3]), .I1(n417), .CO(n30470));
    SB_LUT4 add_3739_11_lut (.I0(GND_net), .I1(n8142[8]), .I2(GND_net), 
            .I3(n30279), .O(n8119[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_18_lut (.I0(GND_net), .I1(n7888[15]), .I2(GND_net), 
            .I3(n30082), .O(n7867[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3754_5_lut (.I0(GND_net), .I1(n8367[2]), .I2(n344), .I3(n30468), 
            .O(n8359[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_11 (.CI(n30279), .I0(n8142[8]), .I1(GND_net), .CO(n30280));
    SB_LUT4 add_3739_10_lut (.I0(GND_net), .I1(n8142[7]), .I2(GND_net), 
            .I3(n30278), .O(n8119[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_18 (.CI(n30082), .I0(n7888[15]), .I1(GND_net), .CO(n30083));
    SB_CARRY add_3754_5 (.CI(n30468), .I0(n8367[2]), .I1(n344), .CO(n30469));
    SB_CARRY add_3739_10 (.CI(n30278), .I0(n8142[7]), .I1(GND_net), .CO(n30279));
    SB_LUT4 add_3719_17_lut (.I0(GND_net), .I1(n7888[14]), .I2(GND_net), 
            .I3(n30081), .O(n7867[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_17 (.CI(n30081), .I0(n7888[14]), .I1(GND_net), .CO(n30082));
    SB_LUT4 add_3739_9_lut (.I0(GND_net), .I1(n8142[6]), .I2(GND_net), 
            .I3(n30277), .O(n8119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_16_lut (.I0(GND_net), .I1(n7888[13]), .I2(GND_net), 
            .I3(n30080), .O(n7867[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_16 (.CI(n30080), .I0(n7888[13]), .I1(GND_net), .CO(n30081));
    SB_LUT4 add_3754_4_lut (.I0(GND_net), .I1(n8367[1]), .I2(n271_adj_3712), 
            .I3(n30467), .O(n8359[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_15_lut (.I0(GND_net), .I1(n7888[12]), .I2(GND_net), 
            .I3(n30079), .O(n7867[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_4 (.CI(n30467), .I0(n8367[1]), .I1(n271_adj_3712), 
            .CO(n30468));
    SB_LUT4 add_3754_3_lut (.I0(GND_net), .I1(n8367[0]), .I2(n198), .I3(n30466), 
            .O(n8359[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_9 (.CI(n30277), .I0(n8142[6]), .I1(GND_net), .CO(n30278));
    SB_CARRY add_3719_15 (.CI(n30079), .I0(n7888[12]), .I1(GND_net), .CO(n30080));
    SB_CARRY add_3754_3 (.CI(n30466), .I0(n8367[0]), .I1(n198), .CO(n30467));
    SB_LUT4 add_3754_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_3713), 
            .I3(GND_net), .O(n8359[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_8_lut (.I0(GND_net), .I1(n8142[5]), .I2(n518), .I3(n30276), 
            .O(n8119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_14_lut (.I0(GND_net), .I1(n7888[11]), .I2(GND_net), 
            .I3(n30078), .O(n7867[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_14 (.CI(n30078), .I0(n7888[11]), .I1(GND_net), .CO(n30079));
    SB_CARRY add_3739_8 (.CI(n30276), .I0(n8142[5]), .I1(n518), .CO(n30277));
    SB_CARRY add_3754_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_3713), .CO(n30466));
    SB_LUT4 add_3753_8_lut (.I0(GND_net), .I1(n8359[5]), .I2(n560), .I3(n30465), 
            .O(n8350[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_7_lut (.I0(GND_net), .I1(n8142[4]), .I2(n445), .I3(n30275), 
            .O(n8119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_13_lut (.I0(GND_net), .I1(n7888[10]), .I2(GND_net), 
            .I3(n30077), .O(n7867[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_13 (.CI(n30077), .I0(n7888[10]), .I1(GND_net), .CO(n30078));
    SB_CARRY add_3739_7 (.CI(n30275), .I0(n8142[4]), .I1(n445), .CO(n30276));
    SB_LUT4 add_3719_12_lut (.I0(GND_net), .I1(n7888[9]), .I2(GND_net), 
            .I3(n30076), .O(n7867[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_12 (.CI(n30076), .I0(n7888[9]), .I1(GND_net), .CO(n30077));
    SB_LUT4 add_3739_6_lut (.I0(GND_net), .I1(n8142[3]), .I2(n372), .I3(n30274), 
            .O(n8119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_7_lut (.I0(GND_net), .I1(n8359[4]), .I2(n487), .I3(n30464), 
            .O(n8350[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_11_lut (.I0(GND_net), .I1(n7888[8]), .I2(GND_net), 
            .I3(n30075), .O(n7867[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_6 (.CI(n30274), .I0(n8142[3]), .I1(n372), .CO(n30275));
    SB_CARRY add_3719_11 (.CI(n30075), .I0(n7888[8]), .I1(GND_net), .CO(n30076));
    SB_LUT4 add_3739_5_lut (.I0(GND_net), .I1(n8142[2]), .I2(n299), .I3(n30273), 
            .O(n8119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_7 (.CI(n30464), .I0(n8359[4]), .I1(n487), .CO(n30465));
    SB_LUT4 add_3719_10_lut (.I0(GND_net), .I1(n7888[7]), .I2(GND_net), 
            .I3(n30074), .O(n7867[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_5 (.CI(n30273), .I0(n8142[2]), .I1(n299), .CO(n30274));
    SB_CARRY add_3719_10 (.CI(n30074), .I0(n7888[7]), .I1(GND_net), .CO(n30075));
    SB_LUT4 add_3739_4_lut (.I0(GND_net), .I1(n8142[1]), .I2(n226), .I3(n30272), 
            .O(n8119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_6_lut (.I0(GND_net), .I1(n8359[3]), .I2(n414), .I3(n30463), 
            .O(n8350[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_9_lut (.I0(GND_net), .I1(n7888[6]), .I2(GND_net), 
            .I3(n30073), .O(n7867[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_9 (.CI(n30073), .I0(n7888[6]), .I1(GND_net), .CO(n30074));
    SB_CARRY add_3739_4 (.CI(n30272), .I0(n8142[1]), .I1(n226), .CO(n30273));
    SB_CARRY add_3753_6 (.CI(n30463), .I0(n8359[3]), .I1(n414), .CO(n30464));
    SB_LUT4 add_3739_3_lut (.I0(GND_net), .I1(n8142[0]), .I2(n153), .I3(n30271), 
            .O(n8119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_8_lut (.I0(GND_net), .I1(n7888[5]), .I2(n524_adj_3714), 
            .I3(n30072), .O(n7867[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_3 (.CI(n30271), .I0(n8142[0]), .I1(n153), .CO(n30272));
    SB_CARRY add_3719_8 (.CI(n30072), .I0(n7888[5]), .I1(n524_adj_3714), 
            .CO(n30073));
    SB_LUT4 add_3719_7_lut (.I0(GND_net), .I1(n7888[4]), .I2(n451_adj_3715), 
            .I3(n30071), .O(n7867[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_5_lut (.I0(GND_net), .I1(n8359[2]), .I2(n341), .I3(n30462), 
            .O(n8350[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_2_lut (.I0(GND_net), .I1(n11_adj_3716), .I2(n80), 
            .I3(GND_net), .O(n8119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_7 (.CI(n30071), .I0(n7888[4]), .I1(n451_adj_3715), 
            .CO(n30072));
    SB_LUT4 add_3719_6_lut (.I0(GND_net), .I1(n7888[3]), .I2(n378_adj_3717), 
            .I3(n30070), .O(n7867[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_2 (.CI(GND_net), .I0(n11_adj_3716), .I1(n80), .CO(n30271));
    SB_CARRY add_3719_6 (.CI(n30070), .I0(n7888[3]), .I1(n378_adj_3717), 
            .CO(n30071));
    SB_LUT4 add_3719_5_lut (.I0(GND_net), .I1(n7888[2]), .I2(n305_adj_3718), 
            .I3(n30069), .O(n7867[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_5 (.CI(n30462), .I0(n8359[2]), .I1(n341), .CO(n30463));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n8095[21]), 
            .I2(GND_net), .I3(n30270), .O(n41237)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3719_5 (.CI(n30069), .I0(n7888[2]), .I1(n305_adj_3718), 
            .CO(n30070));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8095[20]), .I2(GND_net), 
            .I3(n30269), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_4_lut (.I0(GND_net), .I1(n7888[1]), .I2(n232_adj_3719), 
            .I3(n30068), .O(n7867[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_4_lut (.I0(GND_net), .I1(n8359[1]), .I2(n268_adj_3720), 
            .I3(n30461), .O(n8350[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n30269), .I0(n8095[20]), .I1(GND_net), 
            .CO(n30270));
    SB_CARRY add_3719_4 (.CI(n30068), .I0(n7888[1]), .I1(n232_adj_3719), 
            .CO(n30069));
    SB_LUT4 add_3719_3_lut (.I0(GND_net), .I1(n7888[0]), .I2(n159_adj_3721), 
            .I3(n30067), .O(n7867[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_3 (.CI(n30067), .I0(n7888[0]), .I1(n159_adj_3721), 
            .CO(n30068));
    SB_LUT4 add_3719_2_lut (.I0(GND_net), .I1(n17_adj_3722), .I2(n86_adj_3723), 
            .I3(GND_net), .O(n7867[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_2 (.CI(GND_net), .I0(n17_adj_3722), .I1(n86_adj_3723), 
            .CO(n30067));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8095[19]), .I2(GND_net), 
            .I3(n30268), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_4 (.CI(n30461), .I0(n8359[1]), .I1(n268_adj_3720), 
            .CO(n30462));
    SB_LUT4 add_3718_21_lut (.I0(GND_net), .I1(n7867[18]), .I2(GND_net), 
            .I3(n30066), .O(n7845[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_3_lut (.I0(GND_net), .I1(n8359[0]), .I2(n195_adj_3724), 
            .I3(n30460), .O(n8350[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n30268), .I0(n8095[19]), .I1(GND_net), 
            .CO(n30269));
    SB_CARRY add_3753_3 (.CI(n30460), .I0(n8359[0]), .I1(n195_adj_3724), 
            .CO(n30461));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8095[18]), .I2(GND_net), 
            .I3(n30267), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3753_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n8350[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_20_lut (.I0(GND_net), .I1(n7867[17]), .I2(GND_net), 
            .I3(n30065), .O(n7845[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_20 (.CI(n30065), .I0(n7867[17]), .I1(GND_net), .CO(n30066));
    SB_CARRY add_3753_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n30460));
    SB_LUT4 add_3718_19_lut (.I0(GND_net), .I1(n7867[16]), .I2(GND_net), 
            .I3(n30064), .O(n7845[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_19 (.CI(n30064), .I0(n7867[16]), .I1(GND_net), .CO(n30065));
    SB_LUT4 add_3718_18_lut (.I0(GND_net), .I1(n7867[15]), .I2(GND_net), 
            .I3(n30063), .O(n7845[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_9_lut (.I0(GND_net), .I1(n8350[6]), .I2(GND_net), 
            .I3(n30459), .O(n8340[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_18 (.CI(n30063), .I0(n7867[15]), .I1(GND_net), .CO(n30064));
    SB_LUT4 add_3752_8_lut (.I0(GND_net), .I1(n8350[5]), .I2(n557), .I3(n30458), 
            .O(n8340[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n30267), .I0(n8095[18]), .I1(GND_net), 
            .CO(n30268));
    SB_LUT4 add_3718_17_lut (.I0(GND_net), .I1(n7867[14]), .I2(GND_net), 
            .I3(n30062), .O(n7845[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_17 (.CI(n30062), .I0(n7867[14]), .I1(GND_net), .CO(n30063));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8095[17]), .I2(GND_net), 
            .I3(n30266), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_16_lut (.I0(GND_net), .I1(n7867[13]), .I2(GND_net), 
            .I3(n30061), .O(n7845[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n30266), .I0(n8095[17]), .I1(GND_net), 
            .CO(n30267));
    SB_CARRY add_3718_16 (.CI(n30061), .I0(n7867[13]), .I1(GND_net), .CO(n30062));
    SB_CARRY add_3752_8 (.CI(n30458), .I0(n8350[5]), .I1(n557), .CO(n30459));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8095[16]), .I2(GND_net), 
            .I3(n30265), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_15_lut (.I0(GND_net), .I1(n7867[12]), .I2(GND_net), 
            .I3(n30060), .O(n7845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_15 (.CI(n30060), .I0(n7867[12]), .I1(GND_net), .CO(n30061));
    SB_CARRY mult_11_add_1225_19 (.CI(n30265), .I0(n8095[16]), .I1(GND_net), 
            .CO(n30266));
    SB_LUT4 add_3718_14_lut (.I0(GND_net), .I1(n7867[11]), .I2(GND_net), 
            .I3(n30059), .O(n7845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_7_lut (.I0(GND_net), .I1(n8350[4]), .I2(n484), .I3(n30457), 
            .O(n8340[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_7 (.CI(n30457), .I0(n8350[4]), .I1(n484), .CO(n30458));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8095[15]), .I2(GND_net), 
            .I3(n30264), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_14 (.CI(n30059), .I0(n7867[11]), .I1(GND_net), .CO(n30060));
    SB_LUT4 add_3752_6_lut (.I0(GND_net), .I1(n8350[3]), .I2(n411), .I3(n30456), 
            .O(n8340[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n30264), .I0(n8095[15]), .I1(GND_net), 
            .CO(n30265));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8095[14]), .I2(GND_net), 
            .I3(n30263), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_13_lut (.I0(GND_net), .I1(n7867[10]), .I2(GND_net), 
            .I3(n30058), .O(n7845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_13 (.CI(n30058), .I0(n7867[10]), .I1(GND_net), .CO(n30059));
    SB_CARRY add_3752_6 (.CI(n30456), .I0(n8350[3]), .I1(n411), .CO(n30457));
    SB_CARRY mult_11_add_1225_17 (.CI(n30263), .I0(n8095[14]), .I1(GND_net), 
            .CO(n30264));
    SB_LUT4 add_3718_12_lut (.I0(GND_net), .I1(n7867[9]), .I2(GND_net), 
            .I3(n30057), .O(n7845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8095[13]), .I2(GND_net), 
            .I3(n30262), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_12 (.CI(n30057), .I0(n7867[9]), .I1(GND_net), .CO(n30058));
    SB_LUT4 add_3752_5_lut (.I0(GND_net), .I1(n8350[2]), .I2(n338), .I3(n30455), 
            .O(n8340[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n30262), .I0(n8095[13]), .I1(GND_net), 
            .CO(n30263));
    SB_LUT4 add_3718_11_lut (.I0(GND_net), .I1(n7867[8]), .I2(GND_net), 
            .I3(n30056), .O(n7845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8095[12]), .I2(GND_net), 
            .I3(n30261), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_11 (.CI(n30056), .I0(n7867[8]), .I1(GND_net), .CO(n30057));
    SB_CARRY add_3752_5 (.CI(n30455), .I0(n8350[2]), .I1(n338), .CO(n30456));
    SB_CARRY mult_11_add_1225_15 (.CI(n30261), .I0(n8095[12]), .I1(GND_net), 
            .CO(n30262));
    SB_LUT4 add_3718_10_lut (.I0(GND_net), .I1(n7867[7]), .I2(GND_net), 
            .I3(n30055), .O(n7845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8095[11]), .I2(GND_net), 
            .I3(n30260), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_10 (.CI(n30055), .I0(n7867[7]), .I1(GND_net), .CO(n30056));
    SB_LUT4 add_3718_9_lut (.I0(GND_net), .I1(n7867[6]), .I2(GND_net), 
            .I3(n30054), .O(n7845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_4_lut (.I0(GND_net), .I1(n8350[1]), .I2(n265_adj_3726), 
            .I3(n30454), .O(n8340[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n30260), .I0(n8095[11]), .I1(GND_net), 
            .CO(n30261));
    SB_CARRY add_3718_9 (.CI(n30054), .I0(n7867[6]), .I1(GND_net), .CO(n30055));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8095[10]), .I2(GND_net), 
            .I3(n30259), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_8_lut (.I0(GND_net), .I1(n7867[5]), .I2(n521_adj_3727), 
            .I3(n30053), .O(n7845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_4 (.CI(n30454), .I0(n8350[1]), .I1(n265_adj_3726), 
            .CO(n30455));
    SB_CARRY mult_11_add_1225_13 (.CI(n30259), .I0(n8095[10]), .I1(GND_net), 
            .CO(n30260));
    SB_CARRY add_3718_8 (.CI(n30053), .I0(n7867[5]), .I1(n521_adj_3727), 
            .CO(n30054));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8095[9]), .I2(GND_net), 
            .I3(n30258), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_7_lut (.I0(GND_net), .I1(n7867[4]), .I2(n448_adj_3728), 
            .I3(n30052), .O(n7845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_3_lut (.I0(GND_net), .I1(n8350[0]), .I2(n192_adj_3729), 
            .I3(n30453), .O(n8340[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n30258), .I0(n8095[9]), .I1(GND_net), 
            .CO(n30259));
    SB_CARRY add_3718_7 (.CI(n30052), .I0(n7867[4]), .I1(n448_adj_3728), 
            .CO(n30053));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8095[8]), .I2(GND_net), 
            .I3(n30257), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_6_lut (.I0(GND_net), .I1(n7867[3]), .I2(n375_adj_3730), 
            .I3(n30051), .O(n7845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_3 (.CI(n30453), .I0(n8350[0]), .I1(n192_adj_3729), 
            .CO(n30454));
    SB_CARRY mult_11_add_1225_11 (.CI(n30257), .I0(n8095[8]), .I1(GND_net), 
            .CO(n30258));
    SB_CARRY add_3718_6 (.CI(n30051), .I0(n7867[3]), .I1(n375_adj_3730), 
            .CO(n30052));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8095[7]), .I2(GND_net), 
            .I3(n30256), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_5_lut (.I0(GND_net), .I1(n7867[2]), .I2(n302_adj_3731), 
            .I3(n30050), .O(n7845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n8340[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n30256), .I0(n8095[7]), .I1(GND_net), 
            .CO(n30257));
    SB_CARRY add_3718_5 (.CI(n30050), .I0(n7867[2]), .I1(n302_adj_3731), 
            .CO(n30051));
    SB_LUT4 add_3718_4_lut (.I0(GND_net), .I1(n7867[1]), .I2(n229_adj_3732), 
            .I3(n30049), .O(n7845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8095[6]), .I2(GND_net), 
            .I3(n30255), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_4 (.CI(n30049), .I0(n7867[1]), .I1(n229_adj_3732), 
            .CO(n30050));
    SB_LUT4 add_3718_3_lut (.I0(GND_net), .I1(n7867[0]), .I2(n156_adj_3733), 
            .I3(n30048), .O(n7845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n30453));
    SB_CARRY mult_11_add_1225_9 (.CI(n30255), .I0(n8095[6]), .I1(GND_net), 
            .CO(n30256));
    SB_CARRY add_3718_3 (.CI(n30048), .I0(n7867[0]), .I1(n156_adj_3733), 
            .CO(n30049));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8095[5]), .I2(n512), 
            .I3(n30254), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_2_lut (.I0(GND_net), .I1(n14_adj_3734), .I2(n83_adj_3735), 
            .I3(GND_net), .O(n7845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_10_lut (.I0(GND_net), .I1(n8340[7]), .I2(GND_net), 
            .I3(n30452), .O(n8329[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n30254), .I0(n8095[5]), .I1(n512), 
            .CO(n30255));
    SB_CARRY add_3718_2 (.CI(GND_net), .I0(n14_adj_3734), .I1(n83_adj_3735), 
            .CO(n30048));
    SB_LUT4 add_3717_22_lut (.I0(GND_net), .I1(n7845[19]), .I2(GND_net), 
            .I3(n30047), .O(n7822[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8095[4]), .I2(n439), 
            .I3(n30253), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_21_lut (.I0(GND_net), .I1(n7845[18]), .I2(GND_net), 
            .I3(n30046), .O(n7822[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_21 (.CI(n30046), .I0(n7845[18]), .I1(GND_net), .CO(n30047));
    SB_CARRY mult_11_add_1225_7 (.CI(n30253), .I0(n8095[4]), .I1(n439), 
            .CO(n30254));
    SB_LUT4 add_3717_20_lut (.I0(GND_net), .I1(n7845[17]), .I2(GND_net), 
            .I3(n30045), .O(n7822[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_20 (.CI(n30045), .I0(n7845[17]), .I1(GND_net), .CO(n30046));
    SB_LUT4 add_3751_9_lut (.I0(GND_net), .I1(n8340[6]), .I2(GND_net), 
            .I3(n30451), .O(n8329[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8095[3]), .I2(n366), 
            .I3(n30252), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_19_lut (.I0(GND_net), .I1(n7845[16]), .I2(GND_net), 
            .I3(n30044), .O(n7822[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n30252), .I0(n8095[3]), .I1(n366), 
            .CO(n30253));
    SB_CARRY add_3717_19 (.CI(n30044), .I0(n7845[16]), .I1(GND_net), .CO(n30045));
    SB_DFFE \PID_CONTROLLER.integral_1202__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[1]));   // verilog/motorControl.v(40[21:33])
    SB_CARRY add_3751_9 (.CI(n30451), .I0(n8340[6]), .I1(GND_net), .CO(n30452));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8095[2]), .I2(n293), 
            .I3(n30251), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \PID_CONTROLLER.integral_1202__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1202__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[23]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 add_3751_8_lut (.I0(GND_net), .I1(n8340[5]), .I2(n554_adj_3744), 
            .I3(n30450), .O(n8329[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n30251), .I0(n8095[2]), .I1(n293), 
            .CO(n30252));
    SB_LUT4 add_3717_18_lut (.I0(GND_net), .I1(n7845[15]), .I2(GND_net), 
            .I3(n30043), .O(n7822[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_8 (.CI(n30450), .I0(n8340[5]), .I1(n554_adj_3744), 
            .CO(n30451));
    SB_LUT4 add_3751_7_lut (.I0(GND_net), .I1(n8340[4]), .I2(n481_adj_3745), 
            .I3(n30449), .O(n8329[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8095[1]), .I2(n220), 
            .I3(n30250), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_18 (.CI(n30043), .I0(n7845[15]), .I1(GND_net), .CO(n30044));
    SB_LUT4 add_3717_17_lut (.I0(GND_net), .I1(n7845[14]), .I2(GND_net), 
            .I3(n30042), .O(n7822[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_17 (.CI(n30042), .I0(n7845[14]), .I1(GND_net), .CO(n30043));
    SB_CARRY mult_11_add_1225_4 (.CI(n30250), .I0(n8095[1]), .I1(n220), 
            .CO(n30251));
    SB_LUT4 add_3717_16_lut (.I0(GND_net), .I1(n7845[13]), .I2(GND_net), 
            .I3(n30041), .O(n7822[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_7 (.CI(n30449), .I0(n8340[4]), .I1(n481_adj_3745), 
            .CO(n30450));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8095[0]), .I2(n147), 
            .I3(n30249), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n30249), .I0(n8095[0]), .I1(n147), 
            .CO(n30250));
    SB_CARRY add_3717_16 (.CI(n30041), .I0(n7845[13]), .I1(GND_net), .CO(n30042));
    SB_LUT4 add_3717_15_lut (.I0(GND_net), .I1(n7845[12]), .I2(GND_net), 
            .I3(n30040), .O(n7822[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_15 (.CI(n30040), .I0(n7845[12]), .I1(GND_net), .CO(n30041));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3746), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_6_lut (.I0(GND_net), .I1(n8340[3]), .I2(n408_adj_3747), 
            .I3(n30448), .O(n8329[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_6 (.CI(n30448), .I0(n8340[3]), .I1(n408_adj_3747), 
            .CO(n30449));
    SB_LUT4 add_3751_5_lut (.I0(GND_net), .I1(n8340[2]), .I2(n335_adj_3748), 
            .I3(n30447), .O(n8329[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_3746), .I1(n74), 
            .CO(n30249));
    SB_LUT4 add_3717_14_lut (.I0(GND_net), .I1(n7845[11]), .I2(GND_net), 
            .I3(n30039), .O(n7822[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_23_lut (.I0(GND_net), .I1(n8119[20]), .I2(GND_net), 
            .I3(n30248), .O(n8095[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_14 (.CI(n30039), .I0(n7845[11]), .I1(GND_net), .CO(n30040));
    SB_LUT4 add_3717_13_lut (.I0(GND_net), .I1(n7845[10]), .I2(GND_net), 
            .I3(n30038), .O(n7822[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_22_lut (.I0(GND_net), .I1(n8119[19]), .I2(GND_net), 
            .I3(n30247), .O(n8095[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_5 (.CI(n30447), .I0(n8340[2]), .I1(n335_adj_3748), 
            .CO(n30448));
    SB_CARRY add_3717_13 (.CI(n30038), .I0(n7845[10]), .I1(GND_net), .CO(n30039));
    SB_LUT4 add_3717_12_lut (.I0(GND_net), .I1(n7845[9]), .I2(GND_net), 
            .I3(n30037), .O(n7822[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_22 (.CI(n30247), .I0(n8119[19]), .I1(GND_net), .CO(n30248));
    SB_LUT4 add_3751_4_lut (.I0(GND_net), .I1(n8340[1]), .I2(n262_adj_3749), 
            .I3(n30446), .O(n8329[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_4 (.CI(n30446), .I0(n8340[1]), .I1(n262_adj_3749), 
            .CO(n30447));
    SB_LUT4 add_3738_21_lut (.I0(GND_net), .I1(n8119[18]), .I2(GND_net), 
            .I3(n30246), .O(n8095[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_3_lut (.I0(GND_net), .I1(n8340[0]), .I2(n189_adj_3750), 
            .I3(n30445), .O(n8329[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_21 (.CI(n30246), .I0(n8119[18]), .I1(GND_net), .CO(n30247));
    SB_CARRY add_3717_12 (.CI(n30037), .I0(n7845[9]), .I1(GND_net), .CO(n30038));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n29303), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_11_lut (.I0(GND_net), .I1(n7845[8]), .I2(GND_net), 
            .I3(n30036), .O(n7822[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_20_lut (.I0(GND_net), .I1(n8119[17]), .I2(GND_net), 
            .I3(n30245), .O(n8095[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_11 (.CI(n30036), .I0(n7845[8]), .I1(GND_net), .CO(n30037));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n29302), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_24  (.CI(n29302), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n29303));
    SB_CARRY add_3751_3 (.CI(n30445), .I0(n8340[0]), .I1(n189_adj_3750), 
            .CO(n30446));
    SB_CARRY add_3738_20 (.CI(n30245), .I0(n8119[17]), .I1(GND_net), .CO(n30246));
    SB_LUT4 add_3717_10_lut (.I0(GND_net), .I1(n7845[7]), .I2(GND_net), 
            .I3(n30035), .O(n7822[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_2_lut (.I0(GND_net), .I1(n47_adj_3751), .I2(n116_adj_3752), 
            .I3(GND_net), .O(n8329[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_19_lut (.I0(GND_net), .I1(n8119[16]), .I2(GND_net), 
            .I3(n30244), .O(n8095[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_10 (.CI(n30035), .I0(n7845[7]), .I1(GND_net), .CO(n30036));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n29301), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_19 (.CI(n30244), .I0(n8119[16]), .I1(GND_net), .CO(n30245));
    SB_LUT4 add_3717_9_lut (.I0(GND_net), .I1(n7845[6]), .I2(GND_net), 
            .I3(n30034), .O(n7822[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_23  (.CI(n29301), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n29302));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n29300), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_2 (.CI(GND_net), .I0(n47_adj_3751), .I1(n116_adj_3752), 
            .CO(n30445));
    SB_LUT4 add_3738_18_lut (.I0(GND_net), .I1(n8119[15]), .I2(GND_net), 
            .I3(n30243), .O(n8095[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_9 (.CI(n30034), .I0(n7845[6]), .I1(GND_net), .CO(n30035));
    SB_CARRY add_3738_18 (.CI(n30243), .I0(n8119[15]), .I1(GND_net), .CO(n30244));
    SB_LUT4 add_3738_17_lut (.I0(GND_net), .I1(n8119[14]), .I2(GND_net), 
            .I3(n30242), .O(n8095[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_8_lut (.I0(GND_net), .I1(n7845[5]), .I2(n518_adj_3753), 
            .I3(n30033), .O(n7822[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_22  (.CI(n29300), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n29301));
    SB_LUT4 add_3750_11_lut (.I0(GND_net), .I1(n8329[8]), .I2(GND_net), 
            .I3(n30444), .O(n8317[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_17 (.CI(n30242), .I0(n8119[14]), .I1(GND_net), .CO(n30243));
    SB_CARRY add_3717_8 (.CI(n30033), .I0(n7845[5]), .I1(n518_adj_3753), 
            .CO(n30034));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n29299), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_16_lut (.I0(GND_net), .I1(n8119[13]), .I2(GND_net), 
            .I3(n30241), .O(n8095[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_7_lut (.I0(GND_net), .I1(n7845[4]), .I2(n445_adj_3754), 
            .I3(n30032), .O(n7822[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_7 (.CI(n30032), .I0(n7845[4]), .I1(n445_adj_3754), 
            .CO(n30033));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_21  (.CI(n29299), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n29300));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n29298), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3750_10_lut (.I0(GND_net), .I1(n8329[7]), .I2(GND_net), 
            .I3(n30443), .O(n8317[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_16 (.CI(n30241), .I0(n8119[13]), .I1(GND_net), .CO(n30242));
    SB_LUT4 add_3717_6_lut (.I0(GND_net), .I1(n7845[3]), .I2(n372_adj_3755), 
            .I3(n30031), .O(n7822[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_20  (.CI(n29298), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n29299));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n29297), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_15_lut (.I0(GND_net), .I1(n8119[12]), .I2(GND_net), 
            .I3(n30240), .O(n8095[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_10 (.CI(n30443), .I0(n8329[7]), .I1(GND_net), .CO(n30444));
    SB_CARRY add_3717_6 (.CI(n30031), .I0(n7845[3]), .I1(n372_adj_3755), 
            .CO(n30032));
    SB_CARRY add_3738_15 (.CI(n30240), .I0(n8119[12]), .I1(GND_net), .CO(n30241));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_19  (.CI(n29297), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n29298));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n29296), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3750_9_lut (.I0(GND_net), .I1(n8329[6]), .I2(GND_net), 
            .I3(n30442), .O(n8317[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_14_lut (.I0(GND_net), .I1(n8119[11]), .I2(GND_net), 
            .I3(n30239), .O(n8095[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_5_lut (.I0(GND_net), .I1(n7845[2]), .I2(n299_adj_3756), 
            .I3(n30030), .O(n7822[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_18  (.CI(n29296), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n29297));
    SB_CARRY add_3738_14 (.CI(n30239), .I0(n8119[11]), .I1(GND_net), .CO(n30240));
    SB_CARRY add_3717_5 (.CI(n30030), .I0(n7845[2]), .I1(n299_adj_3756), 
            .CO(n30031));
    SB_LUT4 add_3717_4_lut (.I0(GND_net), .I1(n7845[1]), .I2(n226_adj_3757), 
            .I3(n30029), .O(n7822[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n29295), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_17  (.CI(n29295), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n29296));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n29294), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_16  (.CI(n29294), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n29295));
    SB_CARRY add_3750_9 (.CI(n30442), .I0(n8329[6]), .I1(GND_net), .CO(n30443));
    SB_LUT4 add_3738_13_lut (.I0(GND_net), .I1(n8119[10]), .I2(GND_net), 
            .I3(n30238), .O(n8095[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_4 (.CI(n30029), .I0(n7845[1]), .I1(n226_adj_3757), 
            .CO(n30030));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n29293), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_13 (.CI(n30238), .I0(n8119[10]), .I1(GND_net), .CO(n30239));
    SB_LUT4 add_3738_12_lut (.I0(GND_net), .I1(n8119[9]), .I2(GND_net), 
            .I3(n30237), .O(n8095[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_3_lut (.I0(GND_net), .I1(n7845[0]), .I2(n153_adj_3758), 
            .I3(n30028), .O(n7822[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_15  (.CI(n29293), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n29294));
    SB_LUT4 add_3750_8_lut (.I0(GND_net), .I1(n8329[5]), .I2(n551_adj_3759), 
            .I3(n30441), .O(n8317[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_12 (.CI(n30237), .I0(n8119[9]), .I1(GND_net), .CO(n30238));
    SB_CARRY add_3717_3 (.CI(n30028), .I0(n7845[0]), .I1(n153_adj_3758), 
            .CO(n30029));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n29292), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_11_lut (.I0(GND_net), .I1(n8119[8]), .I2(GND_net), 
            .I3(n30236), .O(n8095[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_2_lut (.I0(GND_net), .I1(n11_adj_3760), .I2(n80_adj_3761), 
            .I3(GND_net), .O(n7822[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_14  (.CI(n29292), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n29293));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n29291), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_2 (.CI(GND_net), .I0(n11_adj_3760), .I1(n80_adj_3761), 
            .CO(n30028));
    SB_CARRY add_3750_8 (.CI(n30441), .I0(n8329[5]), .I1(n551_adj_3759), 
            .CO(n30442));
    SB_CARRY add_3738_11 (.CI(n30236), .I0(n8119[8]), .I1(GND_net), .CO(n30237));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7798[21]), 
            .I2(GND_net), .I3(n30027), .O(n6244[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3738_10_lut (.I0(GND_net), .I1(n8119[7]), .I2(GND_net), 
            .I3(n30235), .O(n8095[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n25020), .I1(n7798[20]), .I2(GND_net), 
            .I3(n30026), .O(n3054[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_13  (.CI(n29291), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n29292));
    SB_LUT4 add_3750_7_lut (.I0(GND_net), .I1(n8329[4]), .I2(n478_adj_3762), 
            .I3(n30440), .O(n8317[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_10 (.CI(n30235), .I0(n8119[7]), .I1(GND_net), .CO(n30236));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n29290), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n30026), .I0(n7798[20]), .I1(GND_net), 
            .CO(n30027));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_12  (.CI(n29290), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n29291));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n25020), .I1(n7798[19]), .I2(GND_net), 
            .I3(n30025), .O(n3054[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n29289), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_9_lut (.I0(GND_net), .I1(n8119[6]), .I2(GND_net), 
            .I3(n30234), .O(n8095[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n30025), .I0(n7798[19]), .I1(GND_net), 
            .CO(n30026));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_11  (.CI(n29289), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n29290));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n25020), .I1(n7798[18]), .I2(GND_net), 
            .I3(n30024), .O(n3054[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n29288), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_7 (.CI(n30440), .I0(n8329[4]), .I1(n478_adj_3762), 
            .CO(n30441));
    SB_CARRY add_3738_9 (.CI(n30234), .I0(n8119[6]), .I1(GND_net), .CO(n30235));
    SB_CARRY mult_10_add_1225_21 (.CI(n30024), .I0(n7798[18]), .I1(GND_net), 
            .CO(n30025));
    SB_LUT4 add_3738_8_lut (.I0(GND_net), .I1(n8119[5]), .I2(n515_adj_3763), 
            .I3(n30233), .O(n8095[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n25020), .I1(n7798[17]), .I2(GND_net), 
            .I3(n30023), .O(n3054[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_10  (.CI(n29288), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n29289));
    SB_LUT4 add_3750_6_lut (.I0(GND_net), .I1(n8329[3]), .I2(n405_adj_3764), 
            .I3(n30439), .O(n8317[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_8 (.CI(n30233), .I0(n8119[5]), .I1(n515_adj_3763), 
            .CO(n30234));
    SB_CARRY mult_10_add_1225_20 (.CI(n30023), .I0(n7798[17]), .I1(GND_net), 
            .CO(n30024));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n25020), .I1(n7798[16]), .I2(GND_net), 
            .I3(n30022), .O(n3054[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n29287), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_9  (.CI(n29287), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n29288));
    SB_LUT4 add_3738_7_lut (.I0(GND_net), .I1(n8119[4]), .I2(n442_adj_3765), 
            .I3(n30232), .O(n8095[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n30022), .I0(n7798[16]), .I1(GND_net), 
            .CO(n30023));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n25020), .I1(n7798[15]), .I2(GND_net), 
            .I3(n30021), .O(n3054[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n29286), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_8  (.CI(n29286), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n29287));
    SB_CARRY add_3750_6 (.CI(n30439), .I0(n8329[3]), .I1(n405_adj_3764), 
            .CO(n30440));
    SB_CARRY add_3738_7 (.CI(n30232), .I0(n8119[4]), .I1(n442_adj_3765), 
            .CO(n30233));
    SB_CARRY mult_10_add_1225_18 (.CI(n30021), .I0(n7798[15]), .I1(GND_net), 
            .CO(n30022));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n29285), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_6_lut (.I0(GND_net), .I1(n8119[3]), .I2(n369_adj_3766), 
            .I3(n30231), .O(n8095[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n25020), .I1(n7798[14]), .I2(GND_net), 
            .I3(n30020), .O(n3054[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_7  (.CI(n29285), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n29286));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n29284), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3750_5_lut (.I0(GND_net), .I1(n8329[2]), .I2(n332_adj_3767), 
            .I3(n30438), .O(n8317[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_6 (.CI(n30231), .I0(n8119[3]), .I1(n369_adj_3766), 
            .CO(n30232));
    SB_CARRY mult_10_add_1225_17 (.CI(n30020), .I0(n7798[14]), .I1(GND_net), 
            .CO(n30021));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_6  (.CI(n29284), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n29285));
    SB_CARRY add_3750_5 (.CI(n30438), .I0(n8329[2]), .I1(n332_adj_3767), 
            .CO(n30439));
    SB_LUT4 add_3738_5_lut (.I0(GND_net), .I1(n8119[2]), .I2(n296_adj_3768), 
            .I3(n30230), .O(n8095[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n25020), .I1(n7798[13]), .I2(GND_net), 
            .I3(n30019), .O(n3054[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n29283), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_5 (.CI(n30230), .I0(n8119[2]), .I1(n296_adj_3768), 
            .CO(n30231));
    SB_CARRY mult_10_add_1225_16 (.CI(n30019), .I0(n7798[13]), .I1(GND_net), 
            .CO(n30020));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_5  (.CI(n29283), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n29284));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n29282), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_4_lut (.I0(GND_net), .I1(n8119[1]), .I2(n223_adj_3769), 
            .I3(n30229), .O(n8095[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n25020), .I1(n7798[12]), .I2(GND_net), 
            .I3(n30018), .O(n3054[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3738_4 (.CI(n30229), .I0(n8119[1]), .I1(n223_adj_3769), 
            .CO(n30230));
    SB_LUT4 add_3750_4_lut (.I0(GND_net), .I1(n8329[1]), .I2(n259_adj_3770), 
            .I3(n30437), .O(n8317[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n30018), .I0(n7798[12]), .I1(GND_net), 
            .CO(n30019));
    SB_LUT4 add_3738_3_lut (.I0(GND_net), .I1(n8119[0]), .I2(n150_adj_3771), 
            .I3(n30228), .O(n8095[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n25020), .I1(n7798[11]), .I2(GND_net), 
            .I3(n30017), .O(n3054[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_14 (.CI(n30017), .I0(n7798[11]), .I1(GND_net), 
            .CO(n30018));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_4  (.CI(n29282), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n29283));
    SB_CARRY add_3750_4 (.CI(n30437), .I0(n8329[1]), .I1(n259_adj_3770), 
            .CO(n30438));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n25020), .I1(n7798[10]), .I2(GND_net), 
            .I3(n30016), .O(n3054[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3738_3 (.CI(n30228), .I0(n8119[0]), .I1(n150_adj_3771), 
            .CO(n30229));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n29281), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n30016), .I0(n7798[10]), .I1(GND_net), 
            .CO(n30017));
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_3  (.CI(n29281), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n29282));
    SB_LUT4 \PID_CONTROLLER.integral_1202_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1202_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3750_3_lut (.I0(GND_net), .I1(n8329[0]), .I2(n186_adj_3772), 
            .I3(n30436), .O(n8317[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_2_lut (.I0(GND_net), .I1(n8_adj_3773), .I2(n77_adj_3774), 
            .I3(GND_net), .O(n8095[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n25020), .I1(n7798[9]), .I2(GND_net), 
            .I3(n30015), .O(n3054[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1202_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n29281));
    SB_CARRY add_3750_3 (.CI(n30436), .I0(n8329[0]), .I1(n186_adj_3772), 
            .CO(n30437));
    SB_CARRY add_3738_2 (.CI(GND_net), .I0(n8_adj_3773), .I1(n77_adj_3774), 
            .CO(n30228));
    SB_CARRY mult_10_add_1225_12 (.CI(n30015), .I0(n7798[9]), .I1(GND_net), 
            .CO(n30016));
    SB_LUT4 add_3750_2_lut (.I0(GND_net), .I1(n44_adj_3775), .I2(n113_adj_3776), 
            .I3(GND_net), .O(n8317[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_7_lut (.I0(GND_net), .I1(n37137), .I2(n490_adj_3777), 
            .I3(n30227), .O(n8062[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n25020), .I1(n7798[8]), .I2(GND_net), 
            .I3(n30014), .O(n3054[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3732_6_lut (.I0(GND_net), .I1(n8070[3]), .I2(n417_adj_3778), 
            .I3(n30226), .O(n8062[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_2 (.CI(GND_net), .I0(n44_adj_3775), .I1(n113_adj_3776), 
            .CO(n30436));
    SB_LUT4 add_3749_12_lut (.I0(GND_net), .I1(n8317[9]), .I2(GND_net), 
            .I3(n30435), .O(n8304[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n30014), .I0(n7798[8]), .I1(GND_net), 
            .CO(n30015));
    SB_CARRY add_3732_6 (.CI(n30226), .I0(n8070[3]), .I1(n417_adj_3778), 
            .CO(n30227));
    SB_LUT4 add_3749_11_lut (.I0(GND_net), .I1(n8317[8]), .I2(GND_net), 
            .I3(n30434), .O(n8304[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_5_lut (.I0(GND_net), .I1(n8070[2]), .I2(n344_adj_3779), 
            .I3(n30225), .O(n8062[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n25020), .I1(n7798[7]), .I2(GND_net), 
            .I3(n30013), .O(n3054[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3749_11 (.CI(n30434), .I0(n8317[8]), .I1(GND_net), .CO(n30435));
    SB_LUT4 add_3749_10_lut (.I0(GND_net), .I1(n8317[7]), .I2(GND_net), 
            .I3(n30433), .O(n8304[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_5 (.CI(n30225), .I0(n8070[2]), .I1(n344_adj_3779), 
            .CO(n30226));
    SB_CARRY mult_10_add_1225_10 (.CI(n30013), .I0(n7798[7]), .I1(GND_net), 
            .CO(n30014));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n25020), .I1(n7798[6]), .I2(GND_net), 
            .I3(n30012), .O(n3054[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3732_4_lut (.I0(GND_net), .I1(n8070[1]), .I2(n271_adj_3780), 
            .I3(n30224), .O(n8062[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n30012), .I0(n7798[6]), .I1(GND_net), 
            .CO(n30013));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n25020), .I1(n7798[5]), .I2(n512_adj_3781), 
            .I3(n30011), .O(n3054[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3749_10 (.CI(n30433), .I0(n8317[7]), .I1(GND_net), .CO(n30434));
    SB_CARRY add_3732_4 (.CI(n30224), .I0(n8070[1]), .I1(n271_adj_3780), 
            .CO(n30225));
    SB_LUT4 add_3732_3_lut (.I0(GND_net), .I1(n8070[0]), .I2(n198_adj_3782), 
            .I3(n30223), .O(n8062[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_3 (.CI(n30223), .I0(n8070[0]), .I1(n198_adj_3782), 
            .CO(n30224));
    SB_CARRY mult_10_add_1225_8 (.CI(n30011), .I0(n7798[5]), .I1(n512_adj_3781), 
            .CO(n30012));
    SB_LUT4 add_3749_9_lut (.I0(GND_net), .I1(n8317[6]), .I2(GND_net), 
            .I3(n30432), .O(n8304[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_2_lut (.I0(GND_net), .I1(n56_adj_3783), .I2(n125_adj_3784), 
            .I3(GND_net), .O(n8062[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n25020), .I1(n7798[4]), .I2(n439_adj_3785), 
            .I3(n30010), .O(n3054[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_7 (.CI(n30010), .I0(n7798[4]), .I1(n439_adj_3785), 
            .CO(n30011));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_3887[23]), .I3(n28752), .O(\PID_CONTROLLER.err_23__N_3379 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_3887[22]), .I3(n28751), .O(\PID_CONTROLLER.err_23__N_3379 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n28751), .I0(motor_state[22]), 
            .I1(n1_adj_3887[22]), .CO(n28752));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n25020), .I1(n7798[3]), .I2(n366_adj_3787), 
            .I3(n30009), .O(n3054[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_3887[21]), .I3(n28750), .O(\PID_CONTROLLER.err_23__N_3379 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n28750), .I0(motor_state[21]), 
            .I1(n1_adj_3887[21]), .CO(n28751));
    SB_CARRY add_3732_2 (.CI(GND_net), .I0(n56_adj_3783), .I1(n125_adj_3784), 
            .CO(n30223));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_3887[20]), .I3(n28749), .O(\PID_CONTROLLER.err_23__N_3379 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n30009), .I0(n7798[3]), .I1(n366_adj_3787), 
            .CO(n30010));
    SB_CARRY state_23__I_0_add_2_22 (.CI(n28749), .I0(motor_state[20]), 
            .I1(n1_adj_3887[20]), .CO(n28750));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n25020), .I1(n7798[2]), .I2(n293_adj_3790), 
            .I3(n30008), .O(n3054[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_3887[19]), .I3(n28748), .O(\PID_CONTROLLER.err_23__N_3379 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n30008), .I0(n7798[2]), .I1(n293_adj_3790), 
            .CO(n30009));
    SB_CARRY state_23__I_0_add_2_21 (.CI(n28748), .I0(motor_state[19]), 
            .I1(n1_adj_3887[19]), .CO(n28749));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_3887[18]), .I3(n28747), .O(\PID_CONTROLLER.err_23__N_3379 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n28747), .I0(motor_state[18]), 
            .I1(n1_adj_3887[18]), .CO(n28748));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_3887[17]), .I3(n28746), .O(\PID_CONTROLLER.err_23__N_3379 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n28746), .I0(motor_state[17]), 
            .I1(n1_adj_3887[17]), .CO(n28747));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_3887[16]), .I3(n28745), .O(\PID_CONTROLLER.err_23__N_3379 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n28745), .I0(motor_state[16]), 
            .I1(n1_adj_3887[16]), .CO(n28746));
    SB_CARRY add_3749_9 (.CI(n30432), .I0(n8317[6]), .I1(GND_net), .CO(n30433));
    SB_LUT4 add_3731_8_lut (.I0(GND_net), .I1(n8062[5]), .I2(n560_adj_3795), 
            .I3(n30222), .O(n8053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_3887[15]), .I3(n28744), .O(\PID_CONTROLLER.err_23__N_3379 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n28744), .I0(motor_state[15]), 
            .I1(n1_adj_3887[15]), .CO(n28745));
    SB_LUT4 add_3731_7_lut (.I0(GND_net), .I1(n8062[4]), .I2(n487_adj_3797), 
            .I3(n30221), .O(n8053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_3887[14]), .I3(n28743), .O(\PID_CONTROLLER.err_23__N_3379 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n28743), .I0(motor_state[14]), 
            .I1(n1_adj_3887[14]), .CO(n28744));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n25020), .I1(n7798[1]), .I2(n220_adj_3799), 
            .I3(n30007), .O(n3054[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_3887[13]), .I3(n28742), .O(\PID_CONTROLLER.err_23__N_3379 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n28742), .I0(motor_state[13]), 
            .I1(n1_adj_3887[13]), .CO(n28743));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_3887[12]), .I3(n28741), .O(\PID_CONTROLLER.err_23__N_3379 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n28741), .I0(motor_state[12]), 
            .I1(n1_adj_3887[12]), .CO(n28742));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_3887[11]), .I3(n28740), .O(\PID_CONTROLLER.err_23__N_3379 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n28740), .I0(motor_state[11]), 
            .I1(n1_adj_3887[11]), .CO(n28741));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_3887[10]), .I3(n28739), .O(\PID_CONTROLLER.err_23__N_3379 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n30007), .I0(n7798[1]), .I1(n220_adj_3799), 
            .CO(n30008));
    SB_LUT4 add_3749_8_lut (.I0(GND_net), .I1(n8317[5]), .I2(n548_adj_3804), 
            .I3(n30431), .O(n8304[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n28739), .I0(motor_state[10]), 
            .I1(n1_adj_3887[10]), .CO(n28740));
    SB_CARRY add_3731_7 (.CI(n30221), .I0(n8062[4]), .I1(n487_adj_3797), 
            .CO(n30222));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n25020), .I1(n7798[0]), .I2(n147_adj_3805), 
            .I3(n30006), .O(n3054[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_3887[9]), .I3(n28738), .O(\PID_CONTROLLER.err_23__N_3379 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n30006), .I0(n7798[0]), .I1(n147_adj_3805), 
            .CO(n30007));
    SB_CARRY state_23__I_0_add_2_11 (.CI(n28738), .I0(motor_state[9]), .I1(n1_adj_3887[9]), 
            .CO(n28739));
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_3887[8]), .I3(n28737), .O(\PID_CONTROLLER.err_23__N_3379 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3731_6_lut (.I0(GND_net), .I1(n8062[3]), .I2(n414_adj_3808), 
            .I3(n30220), .O(n8053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n25020), .I1(n5_adj_3809), .I2(n74_adj_3810), 
            .I3(GND_net), .O(n3054[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3731_6 (.CI(n30220), .I0(n8062[3]), .I1(n414_adj_3808), 
            .CO(n30221));
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_3809), .I1(n74_adj_3810), 
            .CO(n30006));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n28737), .I0(motor_state[8]), .I1(n1_adj_3887[8]), 
            .CO(n28738));
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_3887[7]), .I3(n28736), .O(\PID_CONTROLLER.err_23__N_3379 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3749_8 (.CI(n30431), .I0(n8317[5]), .I1(n548_adj_3804), 
            .CO(n30432));
    SB_LUT4 add_3731_5_lut (.I0(GND_net), .I1(n8062[2]), .I2(n341_adj_3812), 
            .I3(n30219), .O(n8053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n28736), .I0(motor_state[7]), .I1(n1_adj_3887[7]), 
            .CO(n28737));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_3887[6]), .I3(n28735), .O(\PID_CONTROLLER.err_23__N_3379 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n28735), .I0(motor_state[6]), .I1(n1_adj_3887[6]), 
            .CO(n28736));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_3887[5]), .I3(n28734), .O(\PID_CONTROLLER.err_23__N_3379 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n28734), .I0(motor_state[5]), .I1(n1_adj_3887[5]), 
            .CO(n28735));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_3887[4]), .I3(n28733), .O(\PID_CONTROLLER.err_23__N_3379 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n28733), .I0(motor_state[4]), .I1(n1_adj_3887[4]), 
            .CO(n28734));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_3887[3]), .I3(n28732), .O(\PID_CONTROLLER.err_23__N_3379 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n28732), .I0(motor_state[3]), .I1(n1_adj_3887[3]), 
            .CO(n28733));
    SB_CARRY add_3731_5 (.CI(n30219), .I0(n8062[2]), .I1(n341_adj_3812), 
            .CO(n30220));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_3887[2]), .I3(n28731), .O(\PID_CONTROLLER.err_23__N_3379 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n28731), .I0(motor_state[2]), .I1(n1_adj_3887[2]), 
            .CO(n28732));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_3887[1]), .I3(n28730), .O(\PID_CONTROLLER.err_23__N_3379 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n28730), .I0(motor_state[1]), .I1(n1_adj_3887[1]), 
            .CO(n28731));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_3887[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3379 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_3887[0]), 
            .CO(n28730));
    SB_LUT4 add_3749_7_lut (.I0(GND_net), .I1(n8317[4]), .I2(n475_adj_3820), 
            .I3(n30430), .O(n8304[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1_adj_3888[23]), 
            .I3(n28729), .O(n47_adj_3629)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[22]), 
            .I3(n28728), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3749_7 (.CI(n30430), .I0(n8317[4]), .I1(n475_adj_3820), 
            .CO(n30431));
    SB_LUT4 add_3731_4_lut (.I0(GND_net), .I1(n8062[1]), .I2(n268_adj_3823), 
            .I3(n30218), .O(n8053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28728), .I0(GND_net), .I1(n1_adj_3888[22]), 
            .CO(n28729));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[21]), 
            .I3(n28727), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28727), .I0(GND_net), .I1(n1_adj_3888[21]), 
            .CO(n28728));
    SB_LUT4 add_3749_6_lut (.I0(GND_net), .I1(n8317[3]), .I2(n402_adj_3825), 
            .I3(n30429), .O(n8304[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_4 (.CI(n30218), .I0(n8062[1]), .I1(n268_adj_3823), 
            .CO(n30219));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[20]), 
            .I3(n28726), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28726), .I0(GND_net), .I1(n1_adj_3888[20]), 
            .CO(n28727));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[19]), 
            .I3(n28725), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28725), .I0(GND_net), .I1(n1_adj_3888[19]), 
            .CO(n28726));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[18]), 
            .I3(n28724), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28724), .I0(GND_net), .I1(n1_adj_3888[18]), 
            .CO(n28725));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[17]), 
            .I3(n28723), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28723), .I0(GND_net), .I1(n1_adj_3888[17]), 
            .CO(n28724));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[16]), 
            .I3(n28722), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28722), .I0(GND_net), .I1(n1_adj_3888[16]), 
            .CO(n28723));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[15]), 
            .I3(n28721), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n28721), .I0(GND_net), .I1(n1_adj_3888[15]), 
            .CO(n28722));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[14]), 
            .I3(n28720), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n28720), .I0(GND_net), .I1(n1_adj_3888[14]), 
            .CO(n28721));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[13]), 
            .I3(n28719), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n28719), .I0(GND_net), .I1(n1_adj_3888[13]), 
            .CO(n28720));
    SB_CARRY add_3749_6 (.CI(n30429), .I0(n8317[3]), .I1(n402_adj_3825), 
            .CO(n30430));
    SB_LUT4 add_3731_3_lut (.I0(GND_net), .I1(n8062[0]), .I2(n195_adj_3834), 
            .I3(n30217), .O(n8053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_3 (.CI(n30217), .I0(n8062[0]), .I1(n195_adj_3834), 
            .CO(n30218));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[12]), 
            .I3(n28718), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n28718), .I0(GND_net), .I1(n1_adj_3888[12]), 
            .CO(n28719));
    SB_LUT4 add_3731_2_lut (.I0(GND_net), .I1(n53_adj_3836), .I2(n122_adj_3837), 
            .I3(GND_net), .O(n8053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[11]), 
            .I3(n28717), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_2 (.CI(GND_net), .I0(n53_adj_3836), .I1(n122_adj_3837), 
            .CO(n30217));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n28717), .I0(GND_net), .I1(n1_adj_3888[11]), 
            .CO(n28718));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[10]), 
            .I3(n28716), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n28716), .I0(GND_net), .I1(n1_adj_3888[10]), 
            .CO(n28717));
    SB_LUT4 add_3749_5_lut (.I0(GND_net), .I1(n8317[2]), .I2(n329_adj_3840), 
            .I3(n30428), .O(n8304[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3730_9_lut (.I0(GND_net), .I1(n8053[6]), .I2(GND_net), 
            .I3(n30216), .O(n8043[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[9]), 
            .I3(n28715), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n28715), .I0(GND_net), .I1(n1_adj_3888[9]), 
            .CO(n28716));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[8]), 
            .I3(n28714), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3730_8_lut (.I0(GND_net), .I1(n8053[5]), .I2(n557_adj_3843), 
            .I3(n30215), .O(n8043[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n28714), .I0(GND_net), .I1(n1_adj_3888[8]), 
            .CO(n28715));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[7]), 
            .I3(n28713), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n28713), .I0(GND_net), .I1(n1_adj_3888[7]), 
            .CO(n28714));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[6]), 
            .I3(n28712), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n28712), .I0(GND_net), .I1(n1_adj_3888[6]), 
            .CO(n28713));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[5]), 
            .I3(n28711), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n28711), .I0(GND_net), .I1(n1_adj_3888[5]), 
            .CO(n28712));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[4]), 
            .I3(n28710), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3749_5 (.CI(n30428), .I0(n8317[2]), .I1(n329_adj_3840), 
            .CO(n30429));
    SB_CARRY add_3730_8 (.CI(n30215), .I0(n8053[5]), .I1(n557_adj_3843), 
            .CO(n30216));
    SB_CARRY unary_minus_16_add_3_6 (.CI(n28710), .I0(GND_net), .I1(n1_adj_3888[4]), 
            .CO(n28711));
    SB_LUT4 add_3749_4_lut (.I0(GND_net), .I1(n8317[1]), .I2(n256_adj_3848), 
            .I3(n30427), .O(n8304[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[3]), 
            .I3(n28709), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n28709), .I0(GND_net), .I1(n1_adj_3888[3]), 
            .CO(n28710));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[2]), 
            .I3(n28708), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3730_7_lut (.I0(GND_net), .I1(n8053[4]), .I2(n484_adj_3851), 
            .I3(n30214), .O(n8043[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n28708), .I0(GND_net), .I1(n1_adj_3888[2]), 
            .CO(n28709));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3888[1]), 
            .I3(n28707), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n28707), .I0(GND_net), .I1(n1_adj_3888[1]), 
            .CO(n28708));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1_adj_3888[0]), 
            .I3(VCC_net), .O(n41179)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_3888[0]), 
            .CO(n28707));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n28706), .O(\PID_CONTROLLER.integral_23__N_3454 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n28705), .O(n45_adj_3684)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n28705), .I0(GND_net), .I1(n1[22]), 
            .CO(n28706));
    SB_CARRY add_3749_4 (.CI(n30427), .I0(n8317[1]), .I1(n256_adj_3848), 
            .CO(n30428));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n28704), .O(n43_adj_3681)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3730_7 (.CI(n30214), .I0(n8053[4]), .I1(n484_adj_3851), 
            .CO(n30215));
    SB_LUT4 add_654_25_lut (.I0(GND_net), .I1(n3054[23]), .I2(n3079[23]), 
            .I3(n28572), .O(duty_23__N_3478[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_654_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3730_6_lut (.I0(GND_net), .I1(n8053[3]), .I2(n411_adj_3858), 
            .I3(n30213), .O(n8043[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3749_3_lut (.I0(GND_net), .I1(n8317[0]), .I2(n183_adj_3859), 
            .I3(n30426), .O(n8304[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_6 (.CI(n30213), .I0(n8053[3]), .I1(n411_adj_3858), 
            .CO(n30214));
    SB_CARRY add_3749_3 (.CI(n30426), .I0(n8317[0]), .I1(n183_adj_3859), 
            .CO(n30427));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n28704), .I0(GND_net), .I1(n1[21]), 
            .CO(n28705));
    SB_LUT4 add_3730_5_lut (.I0(GND_net), .I1(n8053[2]), .I2(n338_adj_3860), 
            .I3(n30212), .O(n8043[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3749_2_lut (.I0(GND_net), .I1(n41_adj_3861), .I2(n110_adj_3862), 
            .I3(GND_net), .O(n8304[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3749_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_5 (.CI(n30212), .I0(n8053[2]), .I1(n338_adj_3860), 
            .CO(n30213));
    SB_CARRY add_3749_2 (.CI(GND_net), .I0(n41_adj_3861), .I1(n110_adj_3862), 
            .CO(n30426));
    SB_LUT4 add_3730_4_lut (.I0(GND_net), .I1(n8053[1]), .I2(n265_adj_3863), 
            .I3(n30211), .O(n8043[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_4 (.CI(n30211), .I0(n8053[1]), .I1(n265_adj_3863), 
            .CO(n30212));
    SB_LUT4 add_3748_13_lut (.I0(GND_net), .I1(n8304[10]), .I2(GND_net), 
            .I3(n30425), .O(n8290[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n28703), .O(n41_adj_3698)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3730_3_lut (.I0(GND_net), .I1(n8053[0]), .I2(n192_adj_3865), 
            .I3(n30210), .O(n8043[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_3 (.CI(n30210), .I0(n8053[0]), .I1(n192_adj_3865), 
            .CO(n30211));
    SB_LUT4 add_3730_2_lut (.I0(GND_net), .I1(n50_adj_3866), .I2(n119_adj_3867), 
            .I3(GND_net), .O(n8043[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_2 (.CI(GND_net), .I0(n50_adj_3866), .I1(n119_adj_3867), 
            .CO(n30210));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n28703), .I0(GND_net), .I1(n1[20]), 
            .CO(n28704));
    SB_LUT4 add_3748_12_lut (.I0(GND_net), .I1(n8304[9]), .I2(GND_net), 
            .I3(n30424), .O(n8290[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_10_lut (.I0(GND_net), .I1(n8043[7]), .I2(GND_net), 
            .I3(n30209), .O(n8032[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_9_lut (.I0(GND_net), .I1(n8043[6]), .I2(GND_net), 
            .I3(n30208), .O(n8032[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3748_12 (.CI(n30424), .I0(n8304[9]), .I1(GND_net), .CO(n30425));
    SB_CARRY add_3729_9 (.CI(n30208), .I0(n8043[6]), .I1(GND_net), .CO(n30209));
    SB_LUT4 add_3748_11_lut (.I0(GND_net), .I1(n8304[8]), .I2(GND_net), 
            .I3(n30423), .O(n8290[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3748_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_652_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256), 
            .I3(GND_net), .O(n3079[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3867));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3866));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3865));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3863));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3862));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3861));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_3860));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3859));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_3858));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256), 
            .I3(GND_net), .O(n3079[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_3851));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3848));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_3843));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3840));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3837));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23721_3_lut_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [21]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n28399));   // verilog/motorControl.v(42[26:37])
    defparam i23721_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3836));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3834));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3825));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3823));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3888[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3820));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3677));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34666_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n41519));
    defparam i34666_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34681_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n41534));
    defparam i34681_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_3812));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23678_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n28340), .I3(n8380[0]), .O(n4_adj_3868));   // verilog/motorControl.v(42[26:37])
    defparam i23678_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3809));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_3808));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n8380[0]), .I3(n28340), .O(n8374[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i23665_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n8374[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23665_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23667_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n28340));   // verilog/motorControl.v(42[26:37])
    defparam i23667_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mux_652_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256), 
            .I3(GND_net), .O(n3079[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3805));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3804));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23696_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8380[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23696_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3676));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3675));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23698_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n28374));   // verilog/motorControl.v(42[26:37])
    defparam i23698_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23647_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_3869), .I3(n8374[1]), .O(n6_adj_3870));   // verilog/motorControl.v(42[26:37])
    defparam i23647_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3799));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_840 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8374[1]), .I3(n4_adj_3869), .O(n8367[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_840.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_3797));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3674));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_841 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8374[0]), .I3(n28297), .O(n8367[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_841.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_3795));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3673));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23639_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n28297), .I3(n8374[0]), .O(n4_adj_3869));   // verilog/motorControl.v(42[26:37])
    defparam i23639_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23628_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n28297));   // verilog/motorControl.v(42[26:37])
    defparam i23628_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23626_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n8367[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23626_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_3790));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_3787));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3672));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3887[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_3785));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3784));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3783));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3782));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_3781));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3780));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3623));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_3779));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_3778));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_3871), .I1(\Kp[4] ), .I2(n8077[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8070[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 i23597_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8088[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23597_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_842 (.I0(n4_adj_3872), .I1(\Kp[3] ), .I2(n8083[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8077[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_842.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_3777));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_843 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_3873));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_843.LUT_INIT = 16'h9c50;
    SB_LUT4 i23533_4_lut (.I0(n8077[2]), .I1(\Kp[4] ), .I2(n6_adj_3871), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_3874));   // verilog/motorControl.v(42[17:23])
    defparam i23533_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_3875));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23564_4_lut (.I0(n8083[1]), .I1(\Kp[3] ), .I2(n4_adj_3872), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_3876));   // verilog/motorControl.v(42[17:23])
    defparam i23564_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23599_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n28267));   // verilog/motorControl.v(42[17:23])
    defparam i23599_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3876), .I1(n11_adj_3875), .I2(n8_adj_3874), 
            .I3(n12_adj_3873), .O(n18_adj_3877));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_3878));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_3878), .I1(n18_adj_3877), .I2(n28267), 
            .I3(n4_adj_3879), .O(n37137));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20320_2_lut_2_lut (.I0(n256), .I1(n6244[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3054[23]));   // verilog/motorControl.v(46[19:35])
    defparam i20320_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3776));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23587_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n28242), .I3(n8088[0]), .O(n4_adj_3879));   // verilog/motorControl.v(42[17:23])
    defparam i23587_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3775));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_844 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8088[0]), .I3(n28242), .O(n8083[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_844.LUT_INIT = 16'h8778;
    SB_LUT4 i23574_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8083[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23574_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_3774));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3773));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3772));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23576_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n28242));   // verilog/motorControl.v(42[17:23])
    defparam i23576_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_3771));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3770));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_3769));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23556_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n28208), .I3(n8083[0]), .O(n4_adj_3872));   // verilog/motorControl.v(42[17:23])
    defparam i23556_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_3768));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3767));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_845 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n8083[0]), .I3(n28208), .O(n8077[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_845.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_3766));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_3765));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3764));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23543_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n8077[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23543_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_3763));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3762));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20297_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25020));   // verilog/motorControl.v(46[19:35])
    defparam i20297_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_3761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3760));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23545_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n28208));   // verilog/motorControl.v(42[17:23])
    defparam i23545_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3759));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3758));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3757));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3756));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_3755));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_3754));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_3753));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3752));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3751));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3750));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23525_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_3880), .I3(n8077[1]), .O(n6_adj_3871));   // verilog/motorControl.v(42[17:23])
    defparam i23525_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_846 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8077[1]), .I3(n4_adj_3880), .O(n8070[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_846.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3749));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_847 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8077[0]), .I3(n28165), .O(n8070[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_847.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3748));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23517_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n28165), .I3(n8077[0]), .O(n4_adj_3880));   // verilog/motorControl.v(42[17:23])
    defparam i23517_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3747));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3746));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3745));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23504_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8070[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23504_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_3744));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23506_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n28165));   // verilog/motorControl.v(42[17:23])
    defparam i23506_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_3735));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3734));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3733));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3732));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_3731));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_3730));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3729));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_3728));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34760_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n41613));   // verilog/motorControl.v(46[19:35])
    defparam i34760_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_3727));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_3580));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3726));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i24_3_lut_3_lut (.I0(PWMLimit[23]), .I1(n256), .I2(n41237), 
            .I3(GND_net), .O(n3079[23]));   // verilog/motorControl.v(47[19:28])
    defparam mux_652_i24_3_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3572));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3562));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3724));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3723));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3722));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_3721));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3720));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3719));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_3718));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_3717));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3716));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_3715));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_3714));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3713));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3712));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_848 (.I0(n6_adj_3870), .I1(\Ki[4] ), .I2(n8374[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8367[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_848.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_3711));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3710));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_849 (.I0(n4_adj_3868), .I1(\Ki[3] ), .I2(n8380[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8374[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_849.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i93_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(GND_net), .I3(GND_net), .O(n137));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i140_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n207));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(GND_net), .I3(GND_net), .O(n68));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_850 (.I0(n28374), .I1(n207), .I2(n68), .I3(n137), 
            .O(n8380[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_851 (.I0(\Ki[1] ), .I1(\Ki[5] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_3881));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_851.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23686_4_lut (.I0(n8380[1]), .I1(\Ki[3] ), .I2(n4_adj_3868), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_3882));   // verilog/motorControl.v(42[26:37])
    defparam i23686_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_852 (.I0(\Ki[2] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral [21]), 
            .I3(\PID_CONTROLLER.integral [23]), .O(n7_adj_3883));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_852.LUT_INIT = 16'h93a0;
    SB_LUT4 i23655_4_lut (.I0(n8374[2]), .I1(\Ki[4] ), .I2(n6_adj_3870), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_3884));   // verilog/motorControl.v(42[26:37])
    defparam i23655_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23709_4_lut (.I0(n68), .I1(n207), .I2(n28374), .I3(n137), 
            .O(n4_adj_3885));   // verilog/motorControl.v(42[26:37])
    defparam i23709_4_lut.LUT_INIT = 16'hd4e8;
    SB_LUT4 i5_4_lut (.I0(n8_adj_3884), .I1(n7_adj_3883), .I2(n6_adj_3882), 
            .I3(n8_adj_3881), .O(n37855));   // verilog/motorControl.v(42[26:37])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_853 (.I0(\Ki[4] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n5_adj_3886));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_853.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_854 (.I0(n5_adj_3886), .I1(n37855), .I2(n4_adj_3885), 
            .I3(n28399), .O(n31074));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_854.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_3709));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3708));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3707));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34935_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n41789));   // verilog/motorControl.v(44[10:25])
    defparam i34935_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3634));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_3706));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_3705));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_3704));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_652_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256), 
            .I3(GND_net), .O(n3079[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_652_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256), 
            .I3(GND_net), .O(n3079[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_652_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3692));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3703));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3478[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3478[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3478[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3478[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3478[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3478[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3478[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3478[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3478[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3478[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3478[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3478[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3478[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3478[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3478[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3478[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3478[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3478[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3478[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3478[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3478[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3478[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3478[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3638));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34766_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n41619));
    defparam i34766_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_3636));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_3644));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34838_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n41692));
    defparam i34838_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_3630));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34600_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n41453));
    defparam i34600_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_3702));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3701));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3622));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    
endmodule
