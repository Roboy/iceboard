// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Oct 23 20:51:05 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_0, PIN_2_c_1, PIN_6_c_0, PIN_7_c_1, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c;
    wire [23:0]color;   // verilog/TinyFPGA_B.v(42[12:17])
    
    wire n25226;
    wire [7:0]blue;   // verilog/TinyFPGA_B.v(43[11:15])
    
    wire send_to_neopixels, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(108[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(109[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(146[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(147[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(148[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(149[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(150[22:24])
    
    wire n36049, n25225, n25224, n25223, n25222;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(153[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(154[22:30])
    
    wire n25221, n25220, n25219, n25218, n25217, n36056;
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(157[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(181[22:33])
    
    wire send_to_neopixels_N_191, n25216;
    wire [22:0]pwm_setpoint_22__N_17;
    
    wire n25215, PIN_13_N_65, n25214, n36160;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n34703, n34698, n34695, n34685, n34681, n34679, n34671, 
        n34669, n34667, n34643;
    wire [31:0]motor_state_23__N_66;
    wire [24:0]displacement_23__N_164;
    wire [23:0]displacement_23__N_40;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n15;
    wire [3:0]state_3__N_298;
    
    wire n25213, n25212, n25211, n25210, n25209, n25208, n25044, 
        n25043, n25207, n25042, n25041, n25040, n25206, n25205, 
        n29071, n25204, n35194, n25039, n35192, n25203, n25038, 
        n25202, n25201, n25200, n25199, n25198, n25037, n25036, 
        n29079, n25197, n2645, n2644, n25196, n25195, n25035, 
        n25194, n25034, n25193, n25033, n24749, n35441, n2643, 
        n25192, n25032, n2572, n2573, n25191, n25031, n25030, 
        n2642, n2641, n25190, n24748, n25189, n2640, n35437, n25188, 
        n25187, n2575, n2574, n2639, n2638, n2637, n2636, n2635, 
        n2634, n2633, n2632, n2631, n2630, n2629, n2628, n2627, 
        n2626, n2625, n2624, n2623, n2622, n2595, n2594, n2593, 
        n2592, n2591, n2590, n2589, n2588, n2587, n2586, n25186, 
        n22030, n25185, n25184, n25183, n25182, n25181, n29081, 
        n383, n382, n381, n380, n379, n378, n377, n376, n375, 
        n374, n373, n372, n371, n370, n369, n35174, n35172, 
        n2585, n24747;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n35166, n2584, n2583, n2582, n7, n15244, n3, n4, n5, 
        n6, n7_adj_3934, n8, n9, n10, n11, n12, n13, n14, 
        n15_adj_3935, n16, n17, n18, n19, n20, n21, n22, n23, 
        n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n36054;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n15475, n24746, n15472, n15469, n15466, n15463;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n15460, n25180, n24745, n35142, n24744, n2, n24743, n24742, 
        n22016, n2_adj_3936, n34633, n24741, n34631, n36052, n740, 
        n6_adj_3937, n24740, n34628, n34626, n24739, n35116, n25158, 
        n25157, n24738, n24737, n25156, n24736, n35463, n24735, 
        n25155, n24734, n15457, n15484, n15454, n15451, n25154, 
        n24733, n15448, n15445, n25005, n15493, n25153, n25004, 
        n25003, n25002, n25152, n15442, n2_adj_3938, n15490, n25001, 
        n25000, n24999, n24998, n24997, n25151, n24996, n24732, 
        n25150, n24995, n24731, n36018, n24730, n6_adj_3939, n24729, 
        n24728, n15439, n25149, n4_adj_3940, n15487, n25148, n24873, 
        n24872, n35082, n24871, n24870, n2_adj_3941, n25147, n15436, 
        n5_adj_3942, n24869, n24868, n21347, n25146, n24867, n25145, 
        n25144, n24866, n24865, n24864, n25143, n15433, n24863, 
        n24862, n25142, n25141, n24861, n25140, n15481, n35443, 
        n15430, n25139, n25138, n25137, n25136, n2581, n2580, 
        n24860, n2579, n35068, n25135, n25134, n24859, n24858, 
        n25133, n24857, n24856, n24855, n25132, n24854, n25131, 
        n25130, n25129, n15_adj_3943, n3761, n31259, n24853, n24852, 
        n24851, n36158, n25128, n25127, n34611, n34608, n15494, 
        n25126, n25125, n35052, n25124, n25123, n25122, n25121, 
        n25120, n34605, n35044, n18493, n35650, n34602, n35034, 
        n36022, n32471, n15387, n35010, n29083, n4573, n35467, 
        n17214, n17213, n17212, n17211, n17210, n17209, n17208, 
        n17207, n17206, n17205, n17204, n17203, n17202, n17201, 
        n17200, n17199, n17198, n17197, n17196, n17195, n17194, 
        n17193, n17192, n17191, n17190, n17189, n17188, n17187, 
        n17186, n17185, n17184, n17183, n17182, n17181, n17180, 
        n17179, n17178, n17177, n17176, n17175, n17174, n17173, 
        n17172, n17171, n17170, n17169, n17168, n17167, n17166, 
        n17165, n17164, n17163, n17162, n17161, n17160, n17159, 
        n17158, n17157, n17156, n17155, n17154, n17153, n17152, 
        n17151, n17150, n17149, n17148, n17147, n17146, n17145, 
        n17144, n17143, n17142, n17141, n17140, n17139, n17138, 
        n17137, n17136, n17135, n17134, n17133, n17132, n17131, 
        n17130, n17129, n17128, n17127, n17126, n17125, n17124, 
        n17123, n17122, n17121, n17120, n17119, n17118, n17117, 
        n17116, n17115, n17114, n17113, n17112, n17111, n17110, 
        n17109, n17108, n17107, n17106, n17105, n17104, n17103, 
        n17102, n17101, n17100, n17099, n17098, n17097, n17096, 
        n17095, n17094, n17093, n17092, n17091, n17090, n17089, 
        n17088, n17087, n17086, n17085, n17084, n17076, n17075, 
        n17074, n17073, n17072, n17071, n17070, n17069, n17068, 
        n17067, n17066, n17065, n17064, n17063, n17062, n17061, 
        n17060, n17059, n17058, n17057, n17056, n17055, n17054, 
        n17053, n17052, n17051, n17050, n17049, n17048, n17047, 
        n17046, n29087, n29089, n17040, n17039, n17038, n17037, 
        n17036, n17035, n17034, n17033, n17032, n17031, n17030, 
        n17029, n17028, n17027, n17026, n17025, n17024, n17023, 
        n17022, n17021, n17020, n17019, n17018, n17013, n249, 
        n248, n224, n35473, n34995, n99, n98, n97, n96, n95, 
        n94, n93, n92, n91, n90, n89, n88, n87, n86, n85, 
        n84, n83, n82, n81, n80, n79, n78, n77, n75, n74, 
        n73, n72, n71, n70, n69, n68, n67, n66, n65, n64, 
        n63, n62, n61, n60, n59, n58, n57, n56, n55, n54, 
        n53, n17006, n17005, n17004, n17003, n17002, n2578, n2577, 
        n2576, n17001, n2421, n925, n25_adj_3944, n24_adj_3945, 
        n23_adj_3946, n22_adj_3947, n21_adj_3948, n20_adj_3949, n19_adj_3950, 
        n18_adj_3951, n17_adj_3952, n16_adj_3953, n15_adj_3954, n14_adj_3955, 
        n13_adj_3956, n12_adj_3957, n11_adj_3958, n10_adj_3959, n9_adj_3960, 
        n8_adj_3961, n7_adj_3962, n6_adj_3963, n5_adj_3964, n4_adj_3965, 
        n3_adj_3966, n36156, n34991, n31114, n4_adj_3967, n17000, 
        n35660, n16999, n4335, n4334, n4333, n4332, n4331, n4330, 
        n4329, n4328, n4327, n4326, n4325, n4324, n4323, n4322, 
        n4321, n4320, n4319, n4318, n4317, n4316, n4315, n4314, 
        n4313, n4312, n15_adj_3968, n34588, quadA_debounced, quadB_debounced, 
        count_enable, n3_adj_3969, n4404, n34586, quadA_debounced_adj_3970, 
        quadB_debounced_adj_3971, count_enable_adj_3972, n25589, n25588, 
        n25587, n25586, n25585, n25584, n25583, n25582, n25581, 
        n25580, n25579, n25578, n25577, n25576, n25575, n25574, 
        n25573, n25572, n22044, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n25571, n25570, n25569, n25568, n34584, n25567, n8_adj_3973, 
        n25566, n25565, n25564, n25563, n25562;
    wire [2:0]r_SM_Main_2__N_3185;
    
    wire n25561, n16998, n25560, n25559, n25558, n25557, n16997, 
        n16996, n16995, n16994, n16993, n16992, n16991, n16990, 
        n25556, n25555, n25554, n34582, n919, n25553, n25552, 
        n25551, n25550, n25549, n25548, n35483, n25547;
    wire [2:0]r_SM_Main_2__N_3259;
    
    wire n25546, n25545, n25544, n16989, n15502, n16988, n16987, 
        n16986, n16985, n16984, n16983, n16982, n16981;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    wire [1:0]reg_B_adj_4409;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n3915, n6555, n4_adj_3976, n4_adj_3977, n35485, n4_adj_3978, 
        n16980, n15373, n25097, n8_adj_3979, n9_adj_3980, n10_adj_3981, 
        n11_adj_3982, n12_adj_3983, n13_adj_3984, n14_adj_3985, n15_adj_3986, 
        n16_adj_3987, n17_adj_3988, n18_adj_3989, n19_adj_3990, n20_adj_3991, 
        n21_adj_3992, n22_adj_3993, n23_adj_3994, n24_adj_3995, n25_adj_3996, 
        n384, n385, n386, n387, n388, n389, n390, n391, n392, 
        n393, n510, n533, n534, n558, n648, n649, n671, n672, 
        n35668, n783, n784, n785, n806, n807, n914, n915, n916, 
        n917, n918, n938, n939, n16770, n1043, n1044, n1045, 
        n1046, n1047, n1048, n1067, n1068, n35495, n1169, n1170, 
        n1171, n1172, n1173, n1174, n1175, n1193, n1194, n35497, 
        n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n1316, n1317, n34778, n34566, n6591, n6592, n6593, n6594, 
        n6595, n6596, n6597, n15395, n1412, n1413, n1414, n1415, 
        n1416, n1417, n1418, n1419, n1420, n1436, n1437, n8_adj_3997, 
        n37085, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
        n1536, n1537, n1538, n35715, n1553, n1554, n36097, n34774, 
        n12917, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
        n6622, n6623, n6624, n34564, n1643, n1644, n1645, n1646, 
        n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1667, 
        n1668, n35672, n34768, n25463, n1754, n1755, n1756, n1757, 
        n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
        n1778, n1779, n6550, n6551, n6552, n6553, n6554, n34761, 
        n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
        n1870, n1871, n1872, n1873, n1874, n1886, n1887, n6564, 
        n6563, n6562, n6561, n6560, n6658, n6659, n6660, n6661, 
        n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, 
        n6670, n6671, n25462, n6559, n34742, n1967, n1968, n1969, 
        n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
        n1978, n1979, n1980, n1991, n1992, n25461, n6682, n6683, 
        n6684, n6685, n6686, n6687, n6688, n6689, n6690, n25460, 
        n25459, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
        n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
        n2093, n2094, n6709, n34562, n2168, n2169, n2170, n2171, 
        n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
        n2180, n2181, n2182, n2183, n6574, n6573, n6572, n2192, 
        n2193, n25458, n6570, n6569, n6568, n6567, n6722, n6723, 
        n6724, n6725, n6726, n6727, n6728, n6729, n6750, n6772, 
        n6795, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
        n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
        n2279, n2280, n2288, n2289, n35507, n25457, n6584, n6583, 
        n6582, n6581, n6580, n6579, n6732, n6733, n6734, n6735, 
        n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
        n6744, n6745, n6746, n6747, n6748, n6749, n6578, n2357, 
        n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, 
        n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
        n2374, n2381, n2382, n6753, n6754, n6755, n6756, n6757, 
        n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
        n6766, n6767, n6768, n6769, n6770, n6771, n2447, n2448, 
        n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
        n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
        n2465, n2471, n2472, n6775, n6776, n6777, n6778, n6779, 
        n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, 
        n6788, n6789, n6790, n6791, n6792, n6793, n6794, n2534, 
        n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
        n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
        n2551, n2552, n2553, n2558, n2559, n35509, n6804, n6805, 
        n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
        n6814, n6815, n6816, n6817, n6818, n6819, n2618, n2619, 
        n2620, n2621, n2622_adj_3998, n2623_adj_3999, n2624_adj_4000, 
        n2625_adj_4001, n2626_adj_4002, n2627_adj_4003, n2628_adj_4004, 
        n2629_adj_4005, n2630_adj_4006, n2631_adj_4007, n2632_adj_4008, 
        n2633_adj_4009, n2634_adj_4010, n2635_adj_4011, n2636_adj_4012, 
        n2637_adj_4013, n2638_adj_4014, n2642_adj_4015, n2643_adj_4016, 
        n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
        n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
        n6842, n6843, n6844, n2699, n2700, n2701, n2702, n2703, 
        n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
        n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
        n2720, n2723, n2724, n2777, n2798, n2799, n2801, n2802, 
        n16979, n16978, n16977, n16976, n16975, n16974, n16973, 
        n16972, n16971, n16970, n16969, n16968, n6590, n6589, 
        n6588, n34718, n34713, n6610, n6609, n6608, n6607, n6606, 
        n6605, n6604, n6603, n6602, n6601, n6600, n6614, n25096, 
        n36041, n25095, n63_adj_4017, n34711, n5_adj_4018, n6639, 
        n6638, n6637, n6636, n6635, n6634, n6633, n6632, n6631, 
        n6630, n6629, n6628, n6627, n6672, n6655, n6654, n6653, 
        n6652, n6651, n6650, n6649, n6648, n6647, n6646, n6645, 
        n6644, n6643, n6681, n6680, n6679, n6678, n6677, n6676, 
        n6675, n6708, n6707, n6706, n6705, n6704, n6703, n6702, 
        n6701, n6700, n6699, n6698, n6697, n6696, n6695, n6694, 
        n6693, n6721, n6720, n6719, n6718, n6717, n6716, n17487, 
        n17486, n17485, n17484, n17483, n17482, n17481, n17479, 
        n29073, n29075, n34560, n35707, n16936, n29095, n29097, 
        n25094, n25093, n16923, n29105, n16918, n29107, n29109, 
        n16907, n16906, n16904, n16899, n29111, n35678, n29113, 
        n29115, n29117, n25092, n29119, n25091, n25090, n29121, 
        n25089, n25088, n25087, n16841, n16840, n16839, n29077, 
        n17467, n17466, n17465, n17464, n17463, n17462, n17461, 
        n17460, n17459, n17458, n17457, n17456, n17455, n17454, 
        n17453, n17452, n17451, n17450, n17449, n17448, n17447, 
        n34323, n17446, n17445, n17444, n17442, n17441, n34322, 
        n17440, n17439, n17438, n17437, n17436, n17435, n17434, 
        n17433, n17432, n17431, n17430, n17429, n17428, n17427, 
        n17426, n17425, n17424, n17423, n17422, n17421, n17420, 
        n6715, n6714, n25086, n6713, n25085, n25084, n35711, n25083, 
        n25082, n25081, n25080, n25079, n25078, n6803, n6802, 
        n6801, n6800, n6799, n6798, n6825, n6824, n6823, n6822, 
        n25077, n25076, n34321, n25075, n25371, n16600, n38, n39, 
        n40, n41, n42, n43, n44, n45, n34320, n29123, n25370, 
        n16835, n25369, n29125, n25368, n34319, n25367, n25366, 
        n25365, n29127, n6_adj_4019, n25364, n25074, n34318, n25363, 
        n25362, n25361, n34317, n34316, n29085, n29091, n29093, 
        n16771, n29129, n16825, n16824, n16823, n29131, n16819, 
        n16816, n34315, n34314, n34313, n16549, n25360, n34312, 
        n25359, n2_adj_4020, n3_adj_4021, n4_adj_4022, n5_adj_4023, 
        n6_adj_4024, n7_adj_4025, n8_adj_4026, n9_adj_4027, n10_adj_4028, 
        n11_adj_4029, n12_adj_4030, n13_adj_4031, n14_adj_4032, n15_adj_4033, 
        n16_adj_4034, n17_adj_4035, n18_adj_4036, n19_adj_4037, n20_adj_4038, 
        n21_adj_4039, n22_adj_4040, n23_adj_4041, n24_adj_4042, n25_adj_4043, 
        n2_adj_4044, n3_adj_4045, n4_adj_4046, n5_adj_4047, n6_adj_4048, 
        n7_adj_4049, n8_adj_4050, n9_adj_4051, n10_adj_4052, n11_adj_4053, 
        n12_adj_4054, n13_adj_4055, n14_adj_4056, n15_adj_4057, n16_adj_4058, 
        n17_adj_4059, n18_adj_4060, n19_adj_4061, n20_adj_4062, n21_adj_4063, 
        n22_adj_4064, n23_adj_4065, n24_adj_4066, n25_adj_4067, n25358, 
        n29133, n16527, n35682, n25357, n25356, n25355, n25354, 
        n25073, n29135, n16501, n34311, n25353, n46, n34310, n34309, 
        n29137, n25352, n34308, n44_adj_4068, n25351, n34307, n25350, 
        n42_adj_4069, n25349, n34306, n34305, n25348, n25347, n25346, 
        n25345, n25344, n25343, n40_adj_4070, n42_adj_4071, n44_adj_4072, 
        n45_adj_4073, n25342, n25341, n25340, n25339, n25338, n34304, 
        n25337, n25336, n38_adj_4074, n40_adj_4075, n42_adj_4076, 
        n43_adj_4077, n35929, n25335, n25334, n25333, n34303, n25332, 
        n36, n38_adj_4078, n40_adj_4079, n41_adj_4080, n36012, n34302, 
        n25072, n25331, n34301, n25330, n34, n36_adj_4081, n38_adj_4082, 
        n39_adj_4083, n41_adj_4084, n43_adj_4085, n35325, n45_adj_4086, 
        n35706, n25329, n34300, n25328, n32, n34_adj_4087, n37, 
        n39_adj_4088, n41_adj_4089, n35620, n43_adj_4090, n34298, 
        n25327, n30, n31, n32_adj_4091, n33, n34_adj_4092, n35, 
        n37_adj_4093, n39_adj_4094, n36014, n41_adj_4095, n42_adj_4096, 
        n43_adj_4097, n45_adj_4098, n25326, n25325, n25324, n28, 
        n29, n30_adj_4099, n31_adj_4100, n32_adj_4101, n33_adj_4102, 
        n35_adj_4103, n37_adj_4104, n35869, n39_adj_4105, n40_adj_4106, 
        n41_adj_4107, n43_adj_4108, n35867, n25323, n25322, n34296, 
        n34295, n25321, n26, n27, n28_adj_4109, n29_adj_4110, n30_adj_4111, 
        n31_adj_4112, n33_adj_4113, n35_adj_4114, n35865, n37_adj_4115, 
        n38_adj_4116, n39_adj_4117, n41_adj_4118, n36051, n34294, 
        n25320, n24_adj_4119, n25_adj_4120, n26_adj_4121, n27_adj_4122, 
        n28_adj_4123, n29_adj_4124, n30_adj_4125, n31_adj_4126, n32_adj_4127, 
        n33_adj_4128, n35_adj_4129, n36_adj_4130, n37_adj_4131, n39_adj_4132, 
        n41_adj_4133, n35720, n43_adj_4134, n44_adj_4135, n45_adj_4136, 
        n35722, n35684, n25319, n25318, n22_adj_4137, n23_adj_4138, 
        n24_adj_4139, n25_adj_4140, n26_adj_4141, n27_adj_4142, n28_adj_4143, 
        n29_adj_4144, n30_adj_4145, n31_adj_4146, n33_adj_4147, n34_adj_4148, 
        n35_adj_4149, n37_adj_4150, n39_adj_4151, n41_adj_4152, n42_adj_4153, 
        n43_adj_4154, n20_adj_4155, n21_adj_4156, n22_adj_4157, n23_adj_4158, 
        n24_adj_4159, n25_adj_4160, n26_adj_4161, n27_adj_4162, n28_adj_4163, 
        n29_adj_4164, n31_adj_4165, n32_adj_4166, n33_adj_4167, n35_adj_4168, 
        n37_adj_4169, n35857, n39_adj_4170, n41_adj_4171, n36079, 
        n36059, n25317, n18_adj_4172, n19_adj_4173, n20_adj_4174, 
        n21_adj_4175, n22_adj_4176, n23_adj_4177, n24_adj_4178, n25_adj_4179, 
        n26_adj_4180, n27_adj_4181, n29_adj_4182, n30_adj_4183, n31_adj_4184, 
        n33_adj_4185, n35_adj_4186, n37_adj_4187, n36061, n39_adj_4188, 
        n41_adj_4189, n42_adj_4190, n43_adj_4191, n45_adj_4192, n35577, 
        n6571, n34293, n25316, n16_adj_4193, n17_adj_4194, n18_adj_4195, 
        n19_adj_4196, n20_adj_4197, n21_adj_4198, n22_adj_4199, n23_adj_4200, 
        n25_adj_4201, n27_adj_4202, n28_adj_4203, n29_adj_4204, n31_adj_4205, 
        n33_adj_4206, n35_adj_4207, n36063, n37_adj_4208, n39_adj_4209, 
        n41_adj_4210, n35580, n43_adj_4211, n36128, n34292, n6585, 
        n34291, n25315, n14_adj_4212, n16_adj_4213, n17_adj_4214, 
        n18_adj_4215, n19_adj_4216, n20_adj_4217, n21_adj_4218, n22_adj_4219, 
        n23_adj_4220, n25_adj_4221, n26_adj_4222, n27_adj_4223, n29_adj_4224, 
        n31_adj_4225, n33_adj_4226, n35953, n35_adj_4227, n37_adj_4228, 
        n35841, n39_adj_4229, n40_adj_4230, n41_adj_4231, n43_adj_4232, 
        n45_adj_4233, n35955, n25314, n25313, n34525, n12_adj_4234, 
        n14_adj_4235, n15_adj_4236, n16_adj_4237, n17_adj_4238, n18_adj_4239, 
        n19_adj_4240, n20_adj_4241, n21_adj_4242, n23_adj_4243, n24_adj_4244, 
        n25_adj_4245, n27_adj_4246, n29_adj_4247, n31_adj_4248, n36067, 
        n33_adj_4249, n35_adj_4250, n35837, n37_adj_4251, n38_adj_4252, 
        n39_adj_4253, n41_adj_4254, n35621, n43_adj_4255, n35835, 
        n25312, n10_adj_4256, n12_adj_4257, n13_adj_4258, n14_adj_4259, 
        n15_adj_4260, n16_adj_4261, n17_adj_4262, n18_adj_4263, n19_adj_4264, 
        n21_adj_4265, n22_adj_4266, n23_adj_4267, n25_adj_4268, n27_adj_4269, 
        n29_adj_4270, n36069, n31_adj_4271, n33_adj_4272, n35831, 
        n35_adj_4273, n36_adj_4274, n37_adj_4275, n39_adj_4276, n41_adj_4277, 
        n36071, n36157, n34290, n25311, n8_adj_4278, n10_adj_4279, 
        n11_adj_4280, n12_adj_4281, n13_adj_4282, n14_adj_4283, n15_adj_4284, 
        n16_adj_4285, n17_adj_4286, n19_adj_4287, n20_adj_4288, n21_adj_4289, 
        n23_adj_4290, n25_adj_4291, n35827, n27_adj_4292, n29_adj_4293, 
        n31_adj_4294, n35825, n33_adj_4295, n34_adj_4296, n35_adj_4297, 
        n37_adj_4298, n39_adj_4299, n35769, n36073, n35771, n25310, 
        n25309, n34514, n6_adj_4300, n8_adj_4301, n9_adj_4302, n10_adj_4303, 
        n11_adj_4304, n12_adj_4305, n13_adj_4306, n14_adj_4307, n15_adj_4308, 
        n17_adj_4309, n19_adj_4310, n21_adj_4311, n23_adj_4312, n35775, 
        n25_adj_4313, n35821, n27_adj_4314, n29_adj_4315, n35819, 
        n31_adj_4316, n32_adj_4317, n33_adj_4318, n35_adj_4319, n37_adj_4320, 
        n39_adj_4321, n36075, n41_adj_4322, n42_adj_4323, n43_adj_4324, 
        n36016, n35815, n34511, n4_adj_4325, n6_adj_4326, n7_adj_4327, 
        n8_adj_4328, n9_adj_4329, n10_adj_4330, n11_adj_4331, n12_adj_4332, 
        n13_adj_4333, n15_adj_4334, n16_adj_4335, n17_adj_4336, n19_adj_4337, 
        n21_adj_4338, n35813, n23_adj_4339, n24_adj_4340, n25_adj_4341, 
        n27_adj_4342, n35811, n29_adj_4343, n30_adj_4344, n31_adj_4345, 
        n33_adj_4346, n35_adj_4347, n35791, n37_adj_4348, n39_adj_4349, 
        n40_adj_4350, n41_adj_4351, n43_adj_4352, n35812, n45_adj_4353, 
        n36043, n34289, n34288, n35625, n35624, n35686, n10_adj_4354, 
        n25308, n35692, n36035, n25307, n16687, n25306, n25071, 
        n25305, n25070, n6558, n6577, n6613, n36034, n6642, n25069, 
        n6712, n34506, n34504, n25284, n25283, n25068, n25282, 
        n34489, n34483, n34481, n34477, n34475, n25281, n25280, 
        n15501, n35578, n15478, n25279, n25278, n25277, n25276, 
        n34421, n25275, n25274, n35698, n25273, n25272, n25271, 
        n25270, n25269, n35700, n25268, n25267, n25266, n25265, 
        n25264, n35704, n4_adj_4355, n36863, n25263, n25262, n25261, 
        n25260, n25259, n34458, n25258, n25257, n34225, n35565, 
        n25256, n25255, n25254, n25253, n25252, n35709, n25251, 
        n25250, n35569, n25249, n25248, n25247, n25246, n25245, 
        n25244, n25243, n25242, n25241, n25240, n35931, n25239, 
        n25238, n25237, n25236, n25235, n25234, n34452, n25233, 
        n25232, n35575, n34450, n25231, n25230, n25229, n36055, 
        n29611, n25228, n25227, n15495, n34445, n13117, n35619, 
        n35618, n5_adj_4356, n29069, n34443, n34441, n34433, n19_adj_4357, 
        n34425, n29103, n34411, n34405, n34403, n34395, n34389, 
        n34381, n36154, n29225, n30199, n30957, n36152, n36150, 
        n36148, n36142, n36141, n36129, n36123, n36143, n36117, 
        n36115, n36151, n36149, n36147, n36145, n36098, n37539, 
        n36089, n36080, n36078, n36068, n34364, n36066, n36064, 
        n36062, n36060, n36017, n36015, n36013, n34360, n36005, 
        n36003, n36001, n36057, n35997, n35995, n35993, n30819, 
        n35991, n35989, n36858, n30817, n30813, n36159, n35959, 
        n35957, n36065, n35952, n35950, n35948, n35942, n36053, 
        n35930, n47, n31_adj_4358, n34358, n34356, n5_adj_4359, 
        n35883, n35872, n35870, n35866, n35852, n35848, n35847, 
        n35842, n35838, n35832, n31841, n35828, n35826, n35822, 
        n35820, n35814, n35788, n35786, n35778, n35774, n35766, 
        n35764, n35760, n35754, n35750, n29853, n6_adj_4360, n35337, 
        n35331, n35323, n34343, n34341, n35845, n35743, n35851;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 add_548_21_lut (.I0(duty[19]), .I1(n36858), .I2(n6), .I3(n24746), 
            .O(pwm_setpoint_22__N_17[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_21 (.CI(n24746), .I0(n36858), .I1(n6), .CO(n24747));
    SB_DFF h2_58 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_40[0]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_59 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF dir_63 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF send_to_neopixels_47 (.Q(send_to_neopixels), .C(LED_c), .D(send_to_neopixels_N_191));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_LUT4 i12743_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n12917), .I3(GND_net), .O(n17130));   // verilog/coms.v(126[12] 289[6])
    defparam i12743_3_lut.LUT_INIT = 16'hcaca;
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.timer({timer}), .GND_net(GND_net), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .n29069(n29069), .VCC_net(VCC_net), .bit_ctr({bit_ctr}), 
            .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), .n29137(n29137), 
            .n29135(n29135), .n29133(n29133), .n29131(n29131), .n29129(n29129), 
            .n29127(n29127), .n29125(n29125), .n29123(n29123), .n29121(n29121), 
            .n29119(n29119), .n29117(n29117), .n29115(n29115), .n29113(n29113), 
            .n29111(n29111), .n29109(n29109), .n29107(n29107), .n29105(n29105), 
            .n29103(n29103), .n29097(n29097), .n29095(n29095), .n29093(n29093), 
            .n29091(n29091), .n29089(n29089), .n29085(n29085), .n29083(n29083), 
            .n29071(n29071), .n29073(n29073), .n29075(n29075), .n34308(n34308), 
            .n19(n19_adj_4357), .n34303(n34303), .\state[0] (state[0]), 
            .\state[1] (state[1]), .start(start), .n34301(n34301), .n34295(n34295), 
            .n34294(n34294), .n34293(n34293), .n34307(n34307), .n34292(n34292), 
            .n34302(n34302), .n34288(n34288), .n34323(n34323), .n34322(n34322), 
            .n34320(n34320), .n34296(n34296), .n34319(n34319), .n34291(n34291), 
            .n34318(n34318), .n34290(n34290), .n34317(n34317), .\state_3__N_298[1] (state_3__N_298[1]), 
            .n15387(n15387), .n919(n919), .n4404(n4404), .\color[18] (color[18]), 
            .\color[19] (color[19]), .n34321(n34321), .\color[17] (color[17]), 
            .\color[16] (color[16]), .n34289(n34289), .n34316(n34316), 
            .n34305(n34305), .n34306(n34306), .n34315(n34315), .n34314(n34314), 
            .n34313(n34313), .n34304(n34304), .n34312(n34312), .n16527(n16527), 
            .n30957(n30957), .n34311(n34311), .PIN_8_c(PIN_8_c), .n29087(n29087), 
            .n16771(n16771), .n29081(n29081), .n17005(n17005), .n17004(n17004), 
            .n17003(n17003), .n17002(n17002), .n17001(n17001), .n17000(n17000), 
            .n16999(n16999), .n16998(n16998), .n16997(n16997), .n16996(n16996), 
            .n16995(n16995), .n16994(n16994), .n16993(n16993), .n16992(n16992), 
            .n16991(n16991), .n16990(n16990), .n16989(n16989), .n16988(n16988), 
            .n16987(n16987), .n16986(n16986), .n16985(n16985), .n16983(n16983), 
            .n16982(n16982), .n16981(n16981), .n16980(n16980), .n16979(n16979), 
            .n16978(n16978), .n16977(n16977), .n16976(n16976), .n16975(n16975), 
            .n16974(n16974), .n29079(n29079), .n16923(n16923), .n34310(n34310), 
            .n29077(n29077), .n34309(n34309), .n22030(n22030), .n29225(n29225), 
            .\color[22] (color[22]), .\color[23] (color[23]), .\color[21] (color[21]), 
            .\color[20] (color[20]), .n22016(n22016)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(55[10] 61[2])
    SB_LUT4 add_548_20_lut (.I0(duty[18]), .I1(n36858), .I2(n7_adj_3934), 
            .I3(n24745), .O(pwm_setpoint_22__N_17[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_3961), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_20 (.CI(n24745), .I0(n36858), .I1(n7_adj_3934), .CO(n24746));
    SB_LUT4 add_548_19_lut (.I0(duty[17]), .I1(n36858), .I2(n8), .I3(n24744), 
            .O(pwm_setpoint_22__N_17[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12744_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n12917), .I3(GND_net), .O(n17131));   // verilog/coms.v(126[12] 289[6])
    defparam i12744_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_19 (.CI(n24744), .I0(n36858), .I1(n8), .CO(n24745));
    SB_LUT4 div_43_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4077));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_548_18_lut (.I0(duty[16]), .I1(n36858), .I2(n9), .I3(n24743), 
            .O(pwm_setpoint_22__N_17[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i659_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_548_18 (.CI(n24743), .I0(n36858), .I1(n9), .CO(n24744));
    SB_LUT4 add_548_17_lut (.I0(duty[15]), .I1(n36858), .I2(n10), .I3(n24742), 
            .O(pwm_setpoint_22__N_17[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_17 (.CI(n24742), .I0(n36858), .I1(n10), .CO(n24743));
    SB_LUT4 add_548_16_lut (.I0(duty[14]), .I1(n36858), .I2(n11), .I3(n24741), 
            .O(pwm_setpoint_22__N_17[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_16 (.CI(n24741), .I0(n36858), .I1(n11), .CO(n24742));
    SB_LUT4 add_548_15_lut (.I0(duty[13]), .I1(n36858), .I2(n12), .I3(n24740), 
            .O(pwm_setpoint_22__N_17[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_15 (.CI(n24740), .I0(n36858), .I1(n12), .CO(n24741));
    SB_LUT4 add_548_14_lut (.I0(duty[12]), .I1(n36858), .I2(n13), .I3(n24739), 
            .O(pwm_setpoint_22__N_17[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_14 (.CI(n24739), .I0(n36858), .I1(n13), .CO(n24740));
    SB_LUT4 div_43_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4074));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_548_13_lut (.I0(duty[11]), .I1(n36858), .I2(n14), .I3(n24738), 
            .O(pwm_setpoint_22__N_17[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_13 (.CI(n24738), .I0(n36858), .I1(n14), .CO(n24739));
    SB_LUT4 add_548_12_lut (.I0(duty[10]), .I1(n36858), .I2(n15_adj_3935), 
            .I3(n24737), .O(pwm_setpoint_22__N_17[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_LessThan_657_i42_3_lut (.I0(n40_adj_4075), .I1(n96), 
            .I2(n43_adj_4077), .I3(GND_net), .O(n42_adj_4076));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30395_4_lut (.I0(n42_adj_4076), .I1(n38_adj_4074), .I2(n43_adj_4077), 
            .I3(n34774), .O(n36034));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30395_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30396_3_lut (.I0(n36034), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n36035));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30396_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut (.I0(n36035), .I1(n15445), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i20087_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4019), .I3(GND_net), 
            .O(n8_adj_3973));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20087_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i20079_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4355), .I3(GND_net), 
            .O(n6_adj_4019));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20079_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_43_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4073));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i20063_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3936));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20063_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_548_12 (.CI(n24737), .I0(n36858), .I1(n15_adj_3935), 
            .CO(n24738));
    SB_LUT4 div_43_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_3962), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4070));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_LessThan_570_i44_3_lut (.I0(n42_adj_4071), .I1(n96), 
            .I2(n45_adj_4073), .I3(GND_net), .O(n44_adj_4072));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30061_4_lut (.I0(n44_adj_4072), .I1(n40_adj_4070), .I2(n45_adj_4073), 
            .I3(n34778), .O(n35700));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30061_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1546 (.I0(n35700), .I1(n15442), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1546.LUT_INIT = 16'hceef;
    SB_LUT4 i20031_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3941));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20031_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20047_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_3940), .I3(GND_net), 
            .O(n6_adj_3939));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20047_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i12745_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n12917), .I3(GND_net), .O(n17132));   // verilog/coms.v(126[12] 289[6])
    defparam i12745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_3963), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4069));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i29985_3_lut (.I0(n42_adj_4069), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n35624));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29985_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i29986_3_lut (.I0(n35624), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n35625));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29986_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1547 (.I0(n35625), .I1(n15439), .I2(n96), .I3(n30819), 
            .O(n806));
    defparam i1_4_lut_adj_1547.LUT_INIT = 16'hefce;
    SB_LUT4 unary_minus_25_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20007_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3938));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20007_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12746_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n12917), .I3(GND_net), .O(n17133));   // verilog/coms.v(126[12] 289[6])
    defparam i12746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_3964), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12747_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n12917), .I3(GND_net), .O(n17134));   // verilog/coms.v(126[12] 289[6])
    defparam i12747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12748_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n12917), .I3(GND_net), .O(n17135));   // verilog/coms.v(126[12] 289[6])
    defparam i12748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12749_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n12917), .I3(GND_net), .O(n17136));   // verilog/coms.v(126[12] 289[6])
    defparam i12749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12750_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n12917), .I3(GND_net), .O(n17137));   // verilog/coms.v(126[12] 289[6])
    defparam i12750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12751_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n12917), .I3(GND_net), .O(n17138));   // verilog/coms.v(126[12] 289[6])
    defparam i12751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44_adj_4068));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30059_3_lut (.I0(n44_adj_4068), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n35698));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30059_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i12752_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n12917), .I3(GND_net), .O(n17139));   // verilog/coms.v(126[12] 289[6])
    defparam i12752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12753_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n12917), .I3(GND_net), .O(n17140));   // verilog/coms.v(126[12] 289[6])
    defparam i12753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1548 (.I0(n35698), .I1(n15436), .I2(n97), .I3(n30817), 
            .O(n671));
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'hefce;
    SB_LUT4 i19991_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i19991_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12754_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n12917), .I3(GND_net), .O(n17141));   // verilog/coms.v(126[12] 289[6])
    defparam i12754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_3965), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12755_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n12917), .I3(GND_net), .O(n17142));   // verilog/coms.v(126[12] 289[6])
    defparam i12755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1549 (.I0(n46), .I1(n15433), .I2(n98), .I3(n30813), 
            .O(n533));
    defparam i1_4_lut_adj_1549.LUT_INIT = 16'hefce;
    SB_LUT4 i12756_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n12917), .I3(GND_net), .O(n17143));   // verilog/coms.v(126[12] 289[6])
    defparam i12756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_3969));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1550 (.I0(n224), .I1(n99), .I2(n15430), .I3(n558), 
            .O(n5_adj_4356));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i1_4_lut_adj_1550.LUT_INIT = 16'h555d;
    SB_LUT4 div_43_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_3966), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29029_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n34225));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29029_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1551 (.I0(n34225), .I1(n15430), .I2(n99), .I3(n5_adj_4356), 
            .O(n392));
    defparam i1_4_lut_adj_1551.LUT_INIT = 16'hefce;
    SB_LUT4 i12757_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n12917), .I3(GND_net), .O(n17144));   // verilog/coms.v(126[12] 289[6])
    defparam i12757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n15490));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(n81), .I1(n15484), .I2(GND_net), .I3(GND_net), 
            .O(n15481));
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1553 (.I0(n84), .I1(n15475), .I2(GND_net), .I3(GND_net), 
            .O(n15472));
    defparam i1_2_lut_adj_1553.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12758_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n12917), .I3(GND_net), .O(n17145));   // verilog/coms.v(126[12] 289[6])
    defparam i12758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1554 (.I0(n87), .I1(n15466), .I2(GND_net), .I3(GND_net), 
            .O(n15463));
    defparam i1_2_lut_adj_1554.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12759_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n12917), .I3(GND_net), .O(n17146));   // verilog/coms.v(126[12] 289[6])
    defparam i12759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(n90), .I1(n15457), .I2(GND_net), .I3(GND_net), 
            .O(n15454));
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(n93), .I1(n15448), .I2(GND_net), .I3(GND_net), 
            .O(n15445));
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(n96), .I1(n15439), .I2(GND_net), .I3(GND_net), 
            .O(n15436));
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'hdddd;
    SB_LUT4 div_43_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_548_11_lut (.I0(duty[9]), .I1(n36858), .I2(n16), .I3(n24736), 
            .O(pwm_setpoint_22__N_17[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15430), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 i31226_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n36863));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i31226_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12807_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n12917), .I3(GND_net), .O(n17194));   // verilog/coms.v(126[12] 289[6])
    defparam i12807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12808_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n12917), .I3(GND_net), .O(n17195));   // verilog/coms.v(126[12] 289[6])
    defparam i12808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12809_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n12917), .I3(GND_net), .O(n17196));   // verilog/coms.v(126[12] 289[6])
    defparam i12809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12810_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n12917), .I3(GND_net), .O(n17197));   // verilog/coms.v(126[12] 289[6])
    defparam i12810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_72_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[0]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_25_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_71_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_66[0]), 
            .I2(n15), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_72_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[1]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_66[1]), 
            .I2(n15), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12811_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n12917), .I3(GND_net), .O(n17198));   // verilog/coms.v(126[12] 289[6])
    defparam i12811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[2]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_66[2]), 
            .I2(n15), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12812_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n12917), .I3(GND_net), .O(n17199));   // verilog/coms.v(126[12] 289[6])
    defparam i12812_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_11 (.CI(n24736), .I0(n36858), .I1(n16), .CO(n24737));
    SB_LUT4 mux_72_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[3]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_66[3]), 
            .I2(n15), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_548_10_lut (.I0(duty[8]), .I1(n36858), .I2(n17), .I3(n24735), 
            .O(pwm_setpoint_22__N_17[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12813_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n12917), .I3(GND_net), .O(n17200));   // verilog/coms.v(126[12] 289[6])
    defparam i12813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_65));   // verilog/TinyFPGA_B.v(164[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_548_10 (.CI(n24735), .I0(n36858), .I1(n17), .CO(n24736));
    SB_LUT4 i12814_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n12917), .I3(GND_net), .O(n17201));   // verilog/coms.v(126[12] 289[6])
    defparam i12814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12760_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n12917), .I3(GND_net), .O(n17147));   // verilog/coms.v(126[12] 289[6])
    defparam i12760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12761_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n12917), .I3(GND_net), .O(n17148));   // verilog/coms.v(126[12] 289[6])
    defparam i12761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12762_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n12917), .I3(GND_net), .O(n17149));   // verilog/coms.v(126[12] 289[6])
    defparam i12762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12763_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n12917), .I3(GND_net), .O(n17150));   // verilog/coms.v(126[12] 289[6])
    defparam i12763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12764_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n12917), .I3(GND_net), .O(n17151));   // verilog/coms.v(126[12] 289[6])
    defparam i12764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_548_9_lut (.I0(duty[7]), .I1(n36858), .I2(n18), .I3(n24734), 
            .O(pwm_setpoint_22__N_17[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12765_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n12917), .I3(GND_net), .O(n17152));   // verilog/coms.v(126[12] 289[6])
    defparam i12765_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_9 (.CI(n24734), .I0(n36858), .I1(n18), .CO(n24735));
    SB_LUT4 i12766_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n12917), .I3(GND_net), .O(n17153));   // verilog/coms.v(126[12] 289[6])
    defparam i12766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_548_8_lut (.I0(duty[6]), .I1(n36858), .I2(n19), .I3(n24733), 
            .O(pwm_setpoint_22__N_17[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_i637_3_lut_3_lut (.I0(n938), .I1(n6553), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12767_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n12917), .I3(GND_net), .O(n17154));   // verilog/coms.v(126[12] 289[6])
    defparam i12767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12768_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n12917), .I3(GND_net), .O(n17155));   // verilog/coms.v(126[12] 289[6])
    defparam i12768_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_8 (.CI(n24733), .I0(n36858), .I1(n19), .CO(n24734));
    SB_LUT4 add_548_7_lut (.I0(duty[5]), .I1(n36858), .I2(n20), .I3(n24732), 
            .O(pwm_setpoint_22__N_17[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_7 (.CI(n24732), .I0(n36858), .I1(n20), .CO(n24733));
    SB_LUT4 i12769_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n12917), .I3(GND_net), .O(n17156));   // verilog/coms.v(126[12] 289[6])
    defparam i12769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12770_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n12917), .I3(GND_net), .O(n17157));   // verilog/coms.v(126[12] 289[6])
    defparam i12770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12771_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n12917), .I3(GND_net), .O(n17158));   // verilog/coms.v(126[12] 289[6])
    defparam i12771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12772_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n12917), .I3(GND_net), .O(n17159));   // verilog/coms.v(126[12] 289[6])
    defparam i12772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12773_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n12917), .I3(GND_net), .O(n17160));   // verilog/coms.v(126[12] 289[6])
    defparam i12773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12774_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n12917), .I3(GND_net), .O(n17161));   // verilog/coms.v(126[12] 289[6])
    defparam i12774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12775_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n12917), .I3(GND_net), .O(n17162));   // verilog/coms.v(126[12] 289[6])
    defparam i12775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12776_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n12917), .I3(GND_net), .O(n17163));   // verilog/coms.v(126[12] 289[6])
    defparam i12776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12777_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n12917), .I3(GND_net), .O(n17164));   // verilog/coms.v(126[12] 289[6])
    defparam i12777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_548_6_lut (.I0(duty[4]), .I1(n36858), .I2(n21), .I3(n24731), 
            .O(pwm_setpoint_22__N_17[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12778_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n12917), .I3(GND_net), .O(n17165));   // verilog/coms.v(126[12] 289[6])
    defparam i12778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12779_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n12917), .I3(GND_net), .O(n17166));   // verilog/coms.v(126[12] 289[6])
    defparam i12779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12780_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n12917), 
            .I3(GND_net), .O(n17167));   // verilog/coms.v(126[12] 289[6])
    defparam i12780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12781_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n12917), 
            .I3(GND_net), .O(n17168));   // verilog/coms.v(126[12] 289[6])
    defparam i12781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12782_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n12917), 
            .I3(GND_net), .O(n17169));   // verilog/coms.v(126[12] 289[6])
    defparam i12782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12783_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n12917), 
            .I3(GND_net), .O(n17170));   // verilog/coms.v(126[12] 289[6])
    defparam i12783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12784_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n12917), 
            .I3(GND_net), .O(n17171));   // verilog/coms.v(126[12] 289[6])
    defparam i12784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12785_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n12917), 
            .I3(GND_net), .O(n17172));   // verilog/coms.v(126[12] 289[6])
    defparam i12785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12786_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n12917), 
            .I3(GND_net), .O(n17173));   // verilog/coms.v(126[12] 289[6])
    defparam i12786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12787_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n12917), 
            .I3(GND_net), .O(n17174));   // verilog/coms.v(126[12] 289[6])
    defparam i12787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12788_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n12917), 
            .I3(GND_net), .O(n17175));   // verilog/coms.v(126[12] 289[6])
    defparam i12788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12789_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n12917), 
            .I3(GND_net), .O(n17176));   // verilog/coms.v(126[12] 289[6])
    defparam i12789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 send_to_neopixels_I_0_1_lut (.I0(send_to_neopixels), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(send_to_neopixels_N_191));   // verilog/TinyFPGA_B.v(48[3] 52[6])
    defparam send_to_neopixels_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12790_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n12917), 
            .I3(GND_net), .O(n17177));   // verilog/coms.v(126[12] 289[6])
    defparam i12790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12791_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n12917), 
            .I3(GND_net), .O(n17178));   // verilog/coms.v(126[12] 289[6])
    defparam i12791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12792_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n12917), 
            .I3(GND_net), .O(n17179));   // verilog/coms.v(126[12] 289[6])
    defparam i12792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12793_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n12917), 
            .I3(GND_net), .O(n17180));   // verilog/coms.v(126[12] 289[6])
    defparam i12793_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_6 (.CI(n24731), .I0(n36858), .I1(n21), .CO(n24732));
    SB_LUT4 add_548_5_lut (.I0(duty[3]), .I1(n36858), .I2(n22), .I3(n24730), 
            .O(pwm_setpoint_22__N_17[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_5 (.CI(n24730), .I0(n36858), .I1(n22), .CO(n24731));
    SB_LUT4 add_548_4_lut (.I0(duty[2]), .I1(n36858), .I2(n23), .I3(n24729), 
            .O(pwm_setpoint_22__N_17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_548_4 (.CI(n24729), .I0(n36858), .I1(n23), .CO(n24730));
    SB_LUT4 add_548_3_lut (.I0(duty[1]), .I1(n36858), .I2(n24), .I3(n24728), 
            .O(pwm_setpoint_22__N_17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_3_lut.LUT_INIT = 16'h8BB8;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 mux_72_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[4]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_66[4]), 
            .I2(n15), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12794_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n12917), 
            .I3(GND_net), .O(n17181));   // verilog/coms.v(126[12] 289[6])
    defparam i12794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12795_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n12917), 
            .I3(GND_net), .O(n17182));   // verilog/coms.v(126[12] 289[6])
    defparam i12795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_72_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[5]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_66[5]), 
            .I2(n15), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_548_3 (.CI(n24728), .I0(n36858), .I1(n24), .CO(n24729));
    SB_LUT4 add_3176_25_lut (.I0(n249), .I1(n36863), .I2(n248), .I3(n25371), 
            .O(displacement_23__N_164[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3176_24_lut (.I0(n393), .I1(n36863), .I2(n392), .I3(n25370), 
            .O(displacement_23__N_164[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_164[23]), 
            .I2(n3_adj_3969), .I3(n24873), .O(displacement_23__N_40[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_24 (.CI(n25370), .I0(n36863), .I1(n392), .CO(n25371));
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_164[22]), 
            .I2(n3_adj_3969), .I3(n24872), .O(displacement_23__N_40[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_23_lut (.I0(n534), .I1(n36863), .I2(n533), .I3(n25369), 
            .O(displacement_23__N_164[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_23 (.CI(n25369), .I0(n36863), .I1(n533), .CO(n25370));
    SB_LUT4 add_3176_22_lut (.I0(n672), .I1(n36863), .I2(n671), .I3(n25368), 
            .O(displacement_23__N_164[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_22 (.CI(n25368), .I0(n36863), .I1(n671), .CO(n25369));
    SB_LUT4 add_548_2_lut (.I0(duty[0]), .I1(n36858), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_72_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[6]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3176_21_lut (.I0(n807), .I1(n36863), .I2(n806), .I3(n25367), 
            .O(displacement_23__N_164[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_21 (.CI(n25367), .I0(n36863), .I1(n806), .CO(n25368));
    SB_LUT4 add_3176_20_lut (.I0(n939), .I1(n36863), .I2(n938), .I3(n25366), 
            .O(displacement_23__N_164[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_20 (.CI(n25366), .I0(n36863), .I1(n938), .CO(n25367));
    SB_LUT4 add_3176_19_lut (.I0(n1068), .I1(n36863), .I2(n1067), .I3(n25365), 
            .O(displacement_23__N_164[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_19 (.CI(n25365), .I0(n36863), .I1(n1067), .CO(n25366));
    SB_LUT4 mux_71_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_66[6]), 
            .I2(n15), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3176_18_lut (.I0(n1194), .I1(n36863), .I2(n1193), .I3(n25364), 
            .O(displacement_23__N_164[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_i808_3_lut_3_lut (.I0(n1193), .I1(n6573), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n15395), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_3996));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_3995));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i807_3_lut_3_lut (.I0(n1193), .I1(n6572), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_3994));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_3993));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i805_3_lut_3_lut (.I0(n1193), .I1(n6570), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3176_18 (.CI(n25364), .I0(n36863), .I1(n1193), .CO(n25365));
    SB_LUT4 add_3176_17_lut (.I0(n1317), .I1(n36863), .I2(n1316), .I3(n25363), 
            .O(displacement_23__N_164[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_17 (.CI(n25363), .I0(n36863), .I1(n1316), .CO(n25364));
    SB_LUT4 mux_72_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[7]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3176_16_lut (.I0(n1437), .I1(n36863), .I2(n1436), .I3(n25362), 
            .O(displacement_23__N_164[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_71_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_66[7]), 
            .I2(n15), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i804_3_lut_3_lut (.I0(n1193), .I1(n6569), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i809_3_lut_3_lut (.I0(n1193), .I1(n6574), .I2(n375), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_3992));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[8]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_66[8]), 
            .I2(n15), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i803_3_lut_3_lut (.I0(n1193), .I1(n6568), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i806_3_lut_3_lut (.I0(n1193), .I1(n6571), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i802_3_lut_3_lut (.I0(n1193), .I1(n6567), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n24872), .I0(displacement_23__N_164[22]), 
            .I1(n3_adj_3969), .CO(n24873));
    SB_CARRY add_548_2 (.CI(VCC_net), .I0(n36858), .I1(n25), .CO(n24728));
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_164[21]), 
            .I2(n3_adj_3969), .I3(n24871), .O(displacement_23__N_40[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n24871), .I0(displacement_23__N_164[21]), 
            .I1(n3_adj_3969), .CO(n24872));
    SB_CARRY add_3176_16 (.CI(n25362), .I0(n36863), .I1(n1436), .CO(n25363));
    SB_LUT4 i1_2_lut_3_lut_adj_1558 (.I0(control_mode[0]), .I1(n15395), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_3943));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i1_2_lut_3_lut_adj_1558.LUT_INIT = 16'hefef;
    SB_LUT4 add_3176_15_lut (.I0(n1554), .I1(n36863), .I2(n1553), .I3(n25361), 
            .O(displacement_23__N_164[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_164[20]), 
            .I2(n3_adj_3969), .I3(n24870), .O(displacement_23__N_40[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_15 (.CI(n25361), .I0(n36863), .I1(n1553), .CO(n25362));
    SB_LUT4 add_3176_14_lut (.I0(n1668), .I1(n36863), .I2(n1667), .I3(n25360), 
            .O(displacement_23__N_164[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n24870), .I0(displacement_23__N_164[20]), 
            .I1(n3_adj_3969), .CO(n24871));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_164[19]), 
            .I2(n6_adj_3937), .I3(n24869), .O(displacement_23__N_40[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_14 (.CI(n25360), .I0(n36863), .I1(n1667), .CO(n25361));
    SB_LUT4 add_3176_13_lut (.I0(n1779), .I1(n36863), .I2(n1778), .I3(n25359), 
            .O(displacement_23__N_164[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n24869), .I0(displacement_23__N_164[19]), 
            .I1(n6_adj_3937), .CO(n24870));
    SB_CARRY add_3176_13 (.CI(n25359), .I0(n36863), .I1(n1778), .CO(n25360));
    SB_LUT4 mux_72_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[9]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3176_12_lut (.I0(n1887), .I1(n36863), .I2(n1886), .I3(n25358), 
            .O(displacement_23__N_164[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_12 (.CI(n25358), .I0(n36863), .I1(n1886), .CO(n25359));
    SB_LUT4 mux_71_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_66[9]), 
            .I2(n15), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4078));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 add_3176_11_lut (.I0(n1992), .I1(n36863), .I2(n1991), .I3(n25357), 
            .O(displacement_23__N_164[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_72_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[10]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3176_11 (.CI(n25357), .I0(n36863), .I1(n1991), .CO(n25358));
    SB_LUT4 add_3176_10_lut (.I0(n2094), .I1(n36863), .I2(n2093), .I3(n25356), 
            .O(displacement_23__N_164[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i29131_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n34768));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29131_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_CARRY add_3176_10 (.CI(n25356), .I0(n36863), .I1(n2093), .CO(n25357));
    SB_LUT4 add_3176_9_lut (.I0(n2193), .I1(n36863), .I2(n2192), .I3(n25355), 
            .O(displacement_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_71_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_66[10]), 
            .I2(n15), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3176_9 (.CI(n25355), .I0(n36863), .I1(n2192), .CO(n25356));
    SB_LUT4 div_43_i889_3_lut_3_lut (.I0(n1316), .I1(n6583), .I2(n1298), 
            .I3(GND_net), .O(n1418));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i891_3_lut_3_lut (.I0(n1316), .I1(n6585), .I2(n376), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i890_3_lut_3_lut (.I0(n1316), .I1(n6584), .I2(n1299), 
            .I3(GND_net), .O(n1419));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3176_8_lut (.I0(n2289), .I1(n36863), .I2(n2288), .I3(n25354), 
            .O(displacement_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_72_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[11]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_66[11]), 
            .I2(n15), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i887_3_lut_3_lut (.I0(n1316), .I1(n6581), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3176_8 (.CI(n25354), .I0(n36863), .I1(n2288), .CO(n25355));
    SB_LUT4 add_3176_7_lut (.I0(n2382), .I1(n36863), .I2(n2381), .I3(n25353), 
            .O(displacement_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 blue_1128_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(blue[7]), 
            .I3(n25463), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_7 (.CI(n25353), .I0(n36863), .I1(n2381), .CO(n25354));
    SB_LUT4 unary_minus_25_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i886_3_lut_3_lut (.I0(n1316), .I1(n6580), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_25_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i888_3_lut_3_lut (.I0(n1316), .I1(n6582), .I2(n1297), 
            .I3(GND_net), .O(n1417));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 blue_1128_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(blue[6]), 
            .I3(n25462), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_6_lut (.I0(n2472), .I1(n36863), .I2(n2471), .I3(n25352), 
            .O(displacement_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_6 (.CI(n25352), .I0(n36863), .I1(n2471), .CO(n25353));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_164[18]), 
            .I2(n7), .I3(n24868), .O(displacement_23__N_40[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_5_lut (.I0(n2559), .I1(n36863), .I2(n2558), .I3(n25351), 
            .O(displacement_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3176_5 (.CI(n25351), .I0(n36863), .I1(n2558), .CO(n25352));
    SB_LUT4 div_43_i885_3_lut_3_lut (.I0(n1316), .I1(n6579), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i884_3_lut_3_lut (.I0(n1316), .I1(n6578), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3176_4_lut (.I0(n2643_adj_4016), .I1(n36863), .I2(n2642_adj_4015), 
            .I3(n25350), .O(displacement_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY blue_1128_add_4_8 (.CI(n25462), .I0(GND_net), .I1(blue[6]), 
            .CO(n25463));
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n24868), .I0(displacement_23__N_164[18]), 
            .I1(n7), .CO(n24869));
    SB_CARRY add_3176_4 (.CI(n25350), .I0(n36863), .I1(n2642_adj_4015), 
            .CO(n25351));
    SB_LUT4 unary_minus_25_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 blue_1128_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(blue[5]), 
            .I3(n25461), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1128_add_4_7 (.CI(n25461), .I0(GND_net), .I1(blue[5]), 
            .CO(n25462));
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_3991));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3176_3_lut (.I0(n2724), .I1(n36863), .I2(n2723), .I3(n25349), 
            .O(displacement_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 blue_1128_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(blue[4]), 
            .I3(n25460), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_3 (.CI(n25349), .I0(n36863), .I1(n2723), .CO(n25350));
    SB_LUT4 add_3176_2_lut (.I0(n2802), .I1(n36863), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_3990));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3176_2 (.CI(VCC_net), .I0(n36863), .I1(n2801), .CO(n25349));
    SB_LUT4 add_3175_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n25348), 
            .O(n6822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1128_add_4_6 (.CI(n25460), .I0(GND_net), .I1(blue[4]), 
            .CO(n25461));
    SB_LUT4 add_3175_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n25347), 
            .O(n6823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_24 (.CI(n25347), .I0(n2700), .I1(n79), .CO(n25348));
    SB_LUT4 add_3175_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n25346), 
            .O(n6824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_23 (.CI(n25346), .I0(n2701), .I1(n80), .CO(n25347));
    SB_LUT4 add_3175_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n25345), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_22 (.CI(n25345), .I0(n2702), .I1(n81), .CO(n25346));
    SB_LUT4 add_3175_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n25344), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12815_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n12917), .I3(GND_net), .O(n17202));   // verilog/coms.v(126[12] 289[6])
    defparam i12815_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3175_21 (.CI(n25344), .I0(n2703), .I1(n82), .CO(n25345));
    SB_LUT4 i12816_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n12917), .I3(GND_net), .O(n17203));   // verilog/coms.v(126[12] 289[6])
    defparam i12816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3175_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n25343), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blue_1128_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(blue[3]), 
            .I3(n25459), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_20 (.CI(n25343), .I0(n2704), .I1(n83), .CO(n25344));
    SB_LUT4 unary_minus_25_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY blue_1128_add_4_5 (.CI(n25459), .I0(GND_net), .I1(blue[3]), 
            .CO(n25460));
    SB_LUT4 div_43_i883_3_lut_3_lut (.I0(n1316), .I1(n6577), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 blue_1128_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(blue[2]), 
            .I3(n25458), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29124_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n34761));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29124_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 add_3175_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n25342), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_19_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3175_19 (.CI(n25342), .I0(n2705), .I1(n84), .CO(n25343));
    SB_LUT4 add_3175_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n25341), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4081));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_CARRY add_3175_18 (.CI(n25341), .I0(n2706), .I1(n85), .CO(n25342));
    SB_LUT4 div_43_i970_3_lut_3_lut (.I0(n1436), .I1(n6596), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3175_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n25340), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i968_3_lut_3_lut (.I0(n1436), .I1(n6594), .I2(n1418), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_25_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i969_3_lut_3_lut (.I0(n1436), .I1(n6595), .I2(n1419), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3175_17 (.CI(n25340), .I0(n2707), .I1(n86), .CO(n25341));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_164[17]), 
            .I2(n8_adj_3979), .I3(n24867), .O(displacement_23__N_40[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3175_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n25339), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_16 (.CI(n25339), .I0(n2708), .I1(n87), .CO(n25340));
    SB_LUT4 add_3175_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n25338), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_15 (.CI(n25338), .I0(n2709), .I1(n88), .CO(n25339));
    SB_LUT4 add_3175_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n25337), 
            .O(n6833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_14 (.CI(n25337), .I0(n2710), .I1(n89), .CO(n25338));
    SB_LUT4 add_3175_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n25336), 
            .O(n6834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i967_3_lut_3_lut (.I0(n1436), .I1(n6593), .I2(n1417), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY blue_1128_add_4_4 (.CI(n25458), .I0(GND_net), .I1(blue[2]), 
            .CO(n25459));
    SB_CARRY add_3175_13 (.CI(n25336), .I0(n2711), .I1(n90), .CO(n25337));
    SB_LUT4 blue_1128_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(blue[1]), 
            .I3(n25457), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_3989));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3175_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n25335), 
            .O(n6835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_57 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_CARRY add_3175_12 (.CI(n25335), .I0(n2712), .I1(n91), .CO(n25336));
    SB_LUT4 mux_72_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[12]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3175_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n25334), 
            .O(n6836)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i964_3_lut_3_lut (.I0(n1436), .I1(n6590), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3175_11 (.CI(n25334), .I0(n2713), .I1(n92), .CO(n25335));
    SB_LUT4 add_3175_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n25333), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i963_3_lut_3_lut (.I0(n1436), .I1(n6589), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3175_10 (.CI(n25333), .I0(n2714), .I1(n93), .CO(n25334));
    SB_LUT4 div_43_i971_3_lut_3_lut (.I0(n1436), .I1(n6597), .I2(n377), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3175_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n25332), 
            .O(n6838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_9 (.CI(n25332), .I0(n2715), .I1(n94), .CO(n25333));
    SB_LUT4 add_3175_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n25331), 
            .O(n6839)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_8 (.CI(n25331), .I0(n2716), .I1(n95), .CO(n25332));
    SB_LUT4 mux_71_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_66[12]), 
            .I2(n15), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3175_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n25330), 
            .O(n6840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_7 (.CI(n25330), .I0(n2717), .I1(n96), .CO(n25331));
    SB_LUT4 div_43_i966_3_lut_3_lut (.I0(n1436), .I1(n6592), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3175_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n25329), 
            .O(n6841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i965_3_lut_3_lut (.I0(n1436), .I1(n6591), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3175_6 (.CI(n25329), .I0(n2718), .I1(n97), .CO(n25330));
    SB_LUT4 add_3175_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n25328), 
            .O(n6842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_40[23]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_CARRY add_3175_5 (.CI(n25328), .I0(n2719), .I1(n98), .CO(n25329));
    SB_LUT4 add_3175_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n25327), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_4 (.CI(n25327), .I0(n2720), .I1(n99), .CO(n25328));
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n24867), .I0(displacement_23__N_164[17]), 
            .I1(n8_adj_3979), .CO(n24868));
    SB_CARRY blue_1128_add_4_3 (.CI(n25457), .I0(GND_net), .I1(blue[1]), 
            .CO(n25458));
    SB_LUT4 add_3175_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n25326), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_3 (.CI(n25326), .I0(n390), .I1(n558), .CO(n25327));
    SB_CARRY add_3175_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n25326));
    SB_LUT4 add_3174_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n25325), 
            .O(n6798)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3174_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n25324), 
            .O(n6799)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i962_3_lut_3_lut (.I0(n1436), .I1(n6588), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3174_22 (.CI(n25324), .I0(n2619), .I1(n80), .CO(n25325));
    SB_LUT4 add_3174_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n25323), 
            .O(n6800)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_21 (.CI(n25323), .I0(n2620), .I1(n81), .CO(n25324));
    SB_LUT4 i29105_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n34742));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29105_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 add_3174_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n25322), 
            .O(n6801)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_20 (.CI(n25322), .I0(n2621), .I1(n82), .CO(n25323));
    SB_LUT4 add_3174_19_lut (.I0(GND_net), .I1(n2622_adj_3998), .I2(n83), 
            .I3(n25321), .O(n6802)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4087));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_CARRY add_3174_19 (.CI(n25321), .I0(n2622_adj_3998), .I1(n83), 
            .CO(n25322));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_164[16]), 
            .I2(n9_adj_3980), .I3(n24866), .O(displacement_23__N_40[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3174_18_lut (.I0(GND_net), .I1(n2623_adj_3999), .I2(n84), 
            .I3(n25320), .O(n6803)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n24866), .I0(displacement_23__N_164[16]), 
            .I1(n9_adj_3980), .CO(n24867));
    SB_CARRY add_3174_18 (.CI(n25320), .I0(n2623_adj_3999), .I1(n84), 
            .CO(n25321));
    SB_LUT4 add_3174_17_lut (.I0(GND_net), .I1(n2624_adj_4000), .I2(n85), 
            .I3(n25319), .O(n6804)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_17 (.CI(n25319), .I0(n2624_adj_4000), .I1(n85), 
            .CO(n25320));
    SB_LUT4 add_3174_16_lut (.I0(GND_net), .I1(n2625_adj_4001), .I2(n86), 
            .I3(n25318), .O(n6805)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_16 (.CI(n25318), .I0(n2625_adj_4001), .I1(n86), 
            .CO(n25319));
    SB_LUT4 add_3174_15_lut (.I0(GND_net), .I1(n2626_adj_4002), .I2(n87), 
            .I3(n25317), .O(n6806)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_15 (.CI(n25317), .I0(n2626_adj_4002), .I1(n87), 
            .CO(n25318));
    SB_LUT4 add_3174_14_lut (.I0(GND_net), .I1(n2627_adj_4003), .I2(n88), 
            .I3(n25316), .O(n6807)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_14 (.CI(n25316), .I0(n2627_adj_4003), .I1(n88), 
            .CO(n25317));
    SB_LUT4 add_3174_13_lut (.I0(GND_net), .I1(n2628_adj_4004), .I2(n89), 
            .I3(n25315), .O(n6808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blue_1128_add_4_2_lut (.I0(GND_net), .I1(send_to_neopixels), 
            .I2(blue[0]), .I3(GND_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1128_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_13 (.CI(n25315), .I0(n2628_adj_4004), .I1(n89), 
            .CO(n25316));
    SB_LUT4 add_3174_12_lut (.I0(GND_net), .I1(n2629_adj_4005), .I2(n90), 
            .I3(n25314), .O(n6809)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_12 (.CI(n25314), .I0(n2629_adj_4005), .I1(n90), 
            .CO(n25315));
    SB_LUT4 add_3174_11_lut (.I0(GND_net), .I1(n2630_adj_4006), .I2(n91), 
            .I3(n25313), .O(n6810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_11 (.CI(n25313), .I0(n2630_adj_4006), .I1(n91), 
            .CO(n25314));
    SB_LUT4 add_3174_10_lut (.I0(GND_net), .I1(n2631_adj_4007), .I2(n92), 
            .I3(n25312), .O(n6811)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_10 (.CI(n25312), .I0(n2631_adj_4007), .I1(n92), 
            .CO(n25313));
    SB_LUT4 add_3174_9_lut (.I0(GND_net), .I1(n2632_adj_4008), .I2(n93), 
            .I3(n25311), .O(n6812)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_3988));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_164[15]), 
            .I2(n10_adj_3981), .I3(n24865), .O(displacement_23__N_40[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_9 (.CI(n25311), .I0(n2632_adj_4008), .I1(n93), .CO(n25312));
    SB_LUT4 add_3174_8_lut (.I0(GND_net), .I1(n2633_adj_4009), .I2(n94), 
            .I3(n25310), .O(n6813)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_8 (.CI(n25310), .I0(n2633_adj_4009), .I1(n94), .CO(n25311));
    SB_LUT4 add_3174_7_lut (.I0(GND_net), .I1(n2634_adj_4010), .I2(n95), 
            .I3(n25309), .O(n6814)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_7 (.CI(n25309), .I0(n2634_adj_4010), .I1(n95), .CO(n25310));
    SB_LUT4 i12817_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n12917), .I3(GND_net), .O(n17204));   // verilog/coms.v(126[12] 289[6])
    defparam i12817_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n24865), .I0(displacement_23__N_164[15]), 
            .I1(n10_adj_3981), .CO(n24866));
    SB_LUT4 add_3174_6_lut (.I0(GND_net), .I1(n2635_adj_4011), .I2(n96), 
            .I3(n25308), .O(n6815)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_6 (.CI(n25308), .I0(n2635_adj_4011), .I1(n96), .CO(n25309));
    SB_CARRY blue_1128_add_4_2 (.CI(GND_net), .I0(send_to_neopixels), .I1(blue[0]), 
            .CO(n25457));
    SB_LUT4 i12818_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n12917), .I3(GND_net), .O(n17205));   // verilog/coms.v(126[12] 289[6])
    defparam i12818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3174_5_lut (.I0(GND_net), .I1(n2636_adj_4012), .I2(n97), 
            .I3(n25307), .O(n6816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_164[14]), 
            .I2(n11_adj_3982), .I3(n24864), .O(displacement_23__N_40[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_5 (.CI(n25307), .I0(n2636_adj_4012), .I1(n97), .CO(n25308));
    SB_LUT4 i12819_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n12917), .I3(GND_net), .O(n17206));   // verilog/coms.v(126[12] 289[6])
    defparam i12819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3174_4_lut (.I0(GND_net), .I1(n2637_adj_4013), .I2(n98), 
            .I3(n25306), .O(n6817)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_4 (.CI(n25306), .I0(n2637_adj_4013), .I1(n98), .CO(n25307));
    SB_LUT4 add_3174_3_lut (.I0(GND_net), .I1(n2638_adj_4014), .I2(n99), 
            .I3(n25305), .O(n6818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_3 (.CI(n25305), .I0(n2638_adj_4014), .I1(n99), .CO(n25306));
    SB_LUT4 mux_72_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[13]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12820_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n12917), .I3(GND_net), .O(n17207));   // verilog/coms.v(126[12] 289[6])
    defparam i12820_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n24864), .I0(displacement_23__N_164[14]), 
            .I1(n11_adj_3982), .CO(n24865));
    SB_LUT4 add_3174_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n6819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n25305));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_164[13]), 
            .I2(n12_adj_3983), .I3(n24863), .O(displacement_23__N_40[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n24863), .I0(displacement_23__N_164[13]), 
            .I1(n12_adj_3983), .CO(n24864));
    SB_LUT4 i12821_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n12917), .I3(GND_net), .O(n17208));   // verilog/coms.v(126[12] 289[6])
    defparam i12821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27_4_lut (.I0(n919), .I1(n15387), .I2(state[0]), .I3(state[1]), 
            .O(n19_adj_4357));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 mux_71_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_66[13]), 
            .I2(n15), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_164[12]), 
            .I2(n13_adj_3984), .I3(n24862), .O(displacement_23__N_40[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n24862), .I0(displacement_23__N_164[12]), 
            .I1(n13_adj_3984), .CO(n24863));
    SB_LUT4 i12796_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n12917), 
            .I3(GND_net), .O(n17183));   // verilog/coms.v(126[12] 289[6])
    defparam i12796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12822_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n12917), .I3(GND_net), .O(n17209));   // verilog/coms.v(126[12] 289[6])
    defparam i12822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12823_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n12917), .I3(GND_net), .O(n17210));   // verilog/coms.v(126[12] 289[6])
    defparam i12823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_164[11]), 
            .I2(n14_adj_3985), .I3(n24861), .O(displacement_23__N_40[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12824_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n12917), .I3(GND_net), .O(n17211));   // verilog/coms.v(126[12] 289[6])
    defparam i12824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12825_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n12917), .I3(GND_net), .O(n17212));   // verilog/coms.v(126[12] 289[6])
    defparam i12825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12826_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n12917), .I3(GND_net), .O(n17213));   // verilog/coms.v(126[12] 289[6])
    defparam i12826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12797_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n12917), 
            .I3(GND_net), .O(n17184));   // verilog/coms.v(126[12] 289[6])
    defparam i12797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12798_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n12917), 
            .I3(GND_net), .O(n17185));   // verilog/coms.v(126[12] 289[6])
    defparam i12798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12799_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n12917), 
            .I3(GND_net), .O(n17186));   // verilog/coms.v(126[12] 289[6])
    defparam i12799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12800_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n12917), 
            .I3(GND_net), .O(n17187));   // verilog/coms.v(126[12] 289[6])
    defparam i12800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12801_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n12917), 
            .I3(GND_net), .O(n17188));   // verilog/coms.v(126[12] 289[6])
    defparam i12801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12802_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n12917), 
            .I3(GND_net), .O(n17189));   // verilog/coms.v(126[12] 289[6])
    defparam i12802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12803_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n12917), 
            .I3(GND_net), .O(n17190));   // verilog/coms.v(126[12] 289[6])
    defparam i12803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_72_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[14]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_66[14]), 
            .I2(n15), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1048_3_lut_3_lut (.I0(n1553), .I1(n6609), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12827_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n12917), .I3(GND_net), .O(n17214));   // verilog/coms.v(126[12] 289[6])
    defparam i12827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1047_3_lut_3_lut (.I0(n1553), .I1(n6608), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1046_3_lut_3_lut (.I0(n1553), .I1(n6607), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_72_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[15]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_66[15]), 
            .I2(n15), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1045_3_lut_3_lut (.I0(n1553), .I1(n6606), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_3987));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[16]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n24861), .I0(displacement_23__N_164[11]), 
            .I1(n14_adj_3985), .CO(n24862));
    SB_LUT4 mux_71_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_66[16]), 
            .I2(n15), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1042_3_lut_3_lut (.I0(n1553), .I1(n6603), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_3986));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_3985));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_3984));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1041_3_lut_3_lut (.I0(n1553), .I1(n6602), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1049_3_lut_3_lut (.I0(n1553), .I1(n6610), .I2(n378), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_164[10]), 
            .I2(n15_adj_3986), .I3(n24860), .O(displacement_23__N_40[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_3983));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[17]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_66[17]), 
            .I2(n15), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n24860), .I0(displacement_23__N_164[10]), 
            .I1(n15_adj_3986), .CO(n24861));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_164[9]), 
            .I2(n16_adj_3987), .I3(n24859), .O(displacement_23__N_40[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1044_3_lut_3_lut (.I0(n1553), .I1(n6605), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_72_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[18]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_66[18]), 
            .I2(n15), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1043_3_lut_3_lut (.I0(n1553), .I1(n6604), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12804_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n12917), .I3(GND_net), .O(n17191));   // verilog/coms.v(126[12] 289[6])
    defparam i12804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1040_3_lut_3_lut (.I0(n1553), .I1(n6601), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1039_3_lut_3_lut (.I0(n1553), .I1(n6600), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_3982));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[19]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_66[19]), 
            .I2(n15), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1123_3_lut_3_lut (.I0(n1667), .I1(n6622), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1121_3_lut_3_lut (.I0(n1667), .I1(n6620), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12805_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n12917), .I3(GND_net), .O(n17192));   // verilog/coms.v(126[12] 289[6])
    defparam i12805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_72_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[20]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_66[20]), 
            .I2(n15), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1118_3_lut_3_lut (.I0(n1667), .I1(n6617), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1124_3_lut_3_lut (.I0(n1667), .I1(n6623), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_3981));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[21]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_66[21]), 
            .I2(n15), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1117_3_lut_3_lut (.I0(n1667), .I1(n6616), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_72_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[22]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_43_i1125_3_lut_3_lut (.I0(n1667), .I1(n6624), .I2(n379), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_66[22]), 
            .I2(n15), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1120_3_lut_3_lut (.I0(n1667), .I1(n6619), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_3980));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_4354));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4354), .I2(control_mode[2]), 
            .I3(GND_net), .O(n15395));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_43_i1119_3_lut_3_lut (.I0(n1667), .I1(n6618), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n15395), 
            .I3(GND_net), .O(n15_adj_3968));   // verilog/TinyFPGA_B.v(185[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_43_i1115_3_lut_3_lut (.I0(n1667), .I1(n6614), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1116_3_lut_3_lut (.I0(n1667), .I1(n6615), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_72_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_3968), .I3(n15_adj_3943), .O(motor_state_23__N_66[23]));   // verilog/TinyFPGA_B.v(185[5] 188[10])
    defparam mux_72_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_71_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_66[23]), 
            .I2(n15), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(184[5] 188[10])
    defparam mux_71_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1114_3_lut_3_lut (.I0(n1667), .I1(n6613), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1122_3_lut_3_lut (.I0(n1667), .I1(n6621), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1197_3_lut_3_lut (.I0(n1778), .I1(n6637), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_3979));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6826), 
            .I3(n2724), .O(n39_adj_4349));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6825), 
            .I3(n2724), .O(n41_adj_4351));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_i1187_3_lut_3_lut (.I0(n1778), .I1(n6627), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_3944), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6823), 
            .I3(n2724), .O(n45_adj_4353));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6824), 
            .I3(n2724), .O(n43_adj_4352));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6831), 
            .I3(n2724), .O(n29_adj_4343));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6830), 
            .I3(n2724), .O(n31_adj_4345));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6835), 
            .I3(n2724), .O(n21_adj_4338));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6834), 
            .I3(n2724), .O(n23_adj_4339));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6833), 
            .I3(n2724), .O(n25_adj_4341));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6837), 
            .I3(n2724), .O(n17_adj_4336));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6836), 
            .I3(n2724), .O(n19_adj_4337));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6842), 
            .I3(n2724), .O(n7_adj_4327));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6841), 
            .I3(n2724), .O(n9_adj_4329));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_i1196_3_lut_3_lut (.I0(n1778), .I1(n6636), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6827), 
            .I3(n2724), .O(n37_adj_4348));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6828), 
            .I3(n2724), .O(n35_adj_4347));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6840), 
            .I3(n2724), .O(n11_adj_4331));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_i1195_3_lut_3_lut (.I0(n1778), .I1(n6635), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6839), 
            .I3(n2724), .O(n13_adj_4333));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6838), 
            .I3(n2724), .O(n15_adj_4334));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6832), 
            .I3(n2724), .O(n27_adj_4342));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6829), 
            .I3(n2724), .O(n33_adj_4346));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_43_i1198_3_lut_3_lut (.I0(n1778), .I1(n6638), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28727_4_lut (.I0(n27_adj_4342), .I1(n15_adj_4334), .I2(n13_adj_4333), 
            .I3(n11_adj_4331), .O(n34364));
    defparam i28727_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4346), 
            .I3(GND_net), .O(n12_adj_4332));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i28719_2_lut (.I0(n33_adj_4346), .I1(n15_adj_4334), .I2(GND_net), 
            .I3(GND_net), .O(n34356));
    defparam i28719_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_43_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4333), 
            .I3(GND_net), .O(n10_adj_4330));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_LessThan_1830_i30_3_lut (.I0(n12_adj_4332), .I1(n83), 
            .I2(n35_adj_4347), .I3(GND_net), .O(n30_adj_4344));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1828_3_lut (.I0(n2720), .I1(n6843), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_43_i1194_3_lut_3_lut (.I0(n1778), .I1(n6634), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3173_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n25284), 
            .O(n6775)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28766_3_lut (.I0(n7_adj_4327), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n34403));
    defparam i28766_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 add_3173_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n25283), 
            .O(n6776)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_21 (.CI(n25283), .I0(n2535), .I1(n81), .CO(n25284));
    SB_LUT4 add_3173_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n25282), 
            .O(n6777)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_20 (.CI(n25282), .I0(n2536), .I1(n82), .CO(n25283));
    SB_LUT4 add_3173_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n25281), 
            .O(n6778)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1192_3_lut_3_lut (.I0(n1778), .I1(n6632), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3173_19 (.CI(n25281), .I0(n2537), .I1(n83), .CO(n25282));
    SB_LUT4 add_3173_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n25280), 
            .O(n6779)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_18 (.CI(n25280), .I0(n2538), .I1(n84), .CO(n25281));
    SB_LUT4 add_3173_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n25279), 
            .O(n6780)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_17 (.CI(n25279), .I0(n2539), .I1(n85), .CO(n25280));
    SB_LUT4 add_3173_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n25278), 
            .O(n6781)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_16 (.CI(n25278), .I0(n2540), .I1(n86), .CO(n25279));
    SB_LUT4 add_3173_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n25277), 
            .O(n6782)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_15 (.CI(n25277), .I0(n2541), .I1(n87), .CO(n25278));
    SB_LUT4 add_3173_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n25276), 
            .O(n6783)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_14 (.CI(n25276), .I0(n2542), .I1(n88), .CO(n25277));
    SB_LUT4 div_43_i1193_3_lut_3_lut (.I0(n1778), .I1(n6633), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n24859), .I0(displacement_23__N_164[9]), 
            .I1(n16_adj_3987), .CO(n24860));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_164[8]), 
            .I2(n17_adj_3988), .I3(n24858), .O(displacement_23__N_40[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3173_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n25275), 
            .O(n6784)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_13 (.CI(n25275), .I0(n2543), .I1(n89), .CO(n25276));
    SB_LUT4 div_43_i1199_3_lut_3_lut (.I0(n1778), .I1(n6639), .I2(n380), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3173_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n25274), 
            .O(n6785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29414_4_lut (.I0(n13_adj_4333), .I1(n11_adj_4331), .I2(n9_adj_4329), 
            .I3(n34403), .O(n35052));
    defparam i29414_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3173_12 (.CI(n25274), .I0(n2544), .I1(n90), .CO(n25275));
    SB_LUT4 i29406_4_lut (.I0(n19_adj_4337), .I1(n17_adj_4336), .I2(n15_adj_4334), 
            .I3(n35052), .O(n35044));
    defparam i29406_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3173_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n25273), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30244_4_lut (.I0(n25_adj_4341), .I1(n23_adj_4339), .I2(n21_adj_4338), 
            .I3(n35044), .O(n35883));
    defparam i30244_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29802_4_lut (.I0(n31_adj_4345), .I1(n29_adj_4343), .I2(n27_adj_4342), 
            .I3(n35883), .O(n35441));
    defparam i29802_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_43_i1191_3_lut_3_lut (.I0(n1778), .I1(n6631), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3173_11 (.CI(n25273), .I0(n2545), .I1(n91), .CO(n25274));
    SB_LUT4 i30379_4_lut (.I0(n37_adj_4348), .I1(n35_adj_4347), .I2(n33_adj_4346), 
            .I3(n35441), .O(n36018));
    defparam i30379_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3173_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n25272), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n24858), .I0(displacement_23__N_164[8]), 
            .I1(n17_adj_3988), .CO(n24859));
    SB_CARRY add_3173_10 (.CI(n25272), .I0(n2546), .I1(n92), .CO(n25273));
    SB_LUT4 add_3173_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n25271), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_9 (.CI(n25271), .I0(n2547), .I1(n93), .CO(n25272));
    SB_LUT4 add_3173_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n25270), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4352), 
            .I3(GND_net), .O(n16_adj_4335));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_3173_8 (.CI(n25270), .I0(n2548), .I1(n94), .CO(n25271));
    SB_LUT4 div_43_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4327), 
            .I3(GND_net), .O(n6_adj_4326));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_3173_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n25269), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_7 (.CI(n25269), .I0(n2549), .I1(n95), .CO(n25270));
    SB_LUT4 add_3173_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n25268), 
            .O(n6791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1190_3_lut_3_lut (.I0(n1778), .I1(n6630), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30174_3_lut (.I0(n6_adj_4326), .I1(n90), .I2(n21_adj_4338), 
            .I3(GND_net), .O(n35813));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30174_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3173_6 (.CI(n25268), .I0(n2550), .I1(n96), .CO(n25269));
    SB_LUT4 add_3173_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n25267), 
            .O(n6792)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1189_3_lut_3_lut (.I0(n1778), .I1(n6629), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3173_5 (.CI(n25267), .I0(n2551), .I1(n97), .CO(n25268));
    SB_LUT4 add_3173_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n25266), 
            .O(n6793)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1188_3_lut_3_lut (.I0(n1778), .I1(n6628), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_40[22]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_LUT4 div_43_i1270_3_lut_3_lut (.I0(n1886), .I1(n6654), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30175_3_lut (.I0(n35813), .I1(n89), .I2(n23_adj_4339), .I3(GND_net), 
            .O(n35814));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30175_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3173_4 (.CI(n25266), .I0(n2552), .I1(n98), .CO(n25267));
    SB_LUT4 add_3173_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n25265), 
            .O(n6794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1260_3_lut_3_lut (.I0(n1886), .I1(n6644), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3173_3 (.CI(n25265), .I0(n2553), .I1(n99), .CO(n25266));
    SB_LUT4 add_3173_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6795)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28744_4_lut (.I0(n21_adj_4338), .I1(n19_adj_4337), .I2(n17_adj_4336), 
            .I3(n9_adj_4329), .O(n34381));
    defparam i28744_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3173_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n25265));
    SB_LUT4 i29353_2_lut (.I0(n43_adj_4352), .I1(n19_adj_4337), .I2(GND_net), 
            .I3(GND_net), .O(n34991));
    defparam i29353_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_43_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4336), 
            .I3(GND_net), .O(n8_adj_4328));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_43_LessThan_1830_i24_3_lut (.I0(n16_adj_4335), .I1(n78), 
            .I2(n45_adj_4353), .I3(GND_net), .O(n24_adj_4340));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1259_3_lut_3_lut (.I0(n1886), .I1(n6643), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1258_3_lut_3_lut (.I0(n1886), .I1(n6642), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_164[7]), 
            .I2(n18_adj_3989), .I3(n24857), .O(displacement_23__N_40[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1269_3_lut_3_lut (.I0(n1886), .I1(n6653), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n24857), .I0(displacement_23__N_164[7]), 
            .I1(n18_adj_3989), .CO(n24858));
    SB_LUT4 div_43_i1267_3_lut_3_lut (.I0(n1886), .I1(n6651), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3172_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n25264), 
            .O(n6753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3172_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n25263), 
            .O(n6754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_20 (.CI(n25263), .I0(n2448), .I1(n82), .CO(n25264));
    SB_LUT4 i29357_4_lut (.I0(n43_adj_4352), .I1(n25_adj_4341), .I2(n23_adj_4339), 
            .I3(n34381), .O(n34995));
    defparam i29357_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30152_4_lut (.I0(n24_adj_4340), .I1(n8_adj_4328), .I2(n45_adj_4353), 
            .I3(n34991), .O(n35791));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30152_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30147_3_lut (.I0(n35814), .I1(n88), .I2(n25_adj_4341), .I3(GND_net), 
            .O(n35786));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30147_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1829_3_lut (.I0(n390), .I1(n6844), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3172_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n25262), 
            .O(n6755)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4325));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30172_3_lut (.I0(n4_adj_4325), .I1(n87), .I2(n27_adj_4342), 
            .I3(GND_net), .O(n35811));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30172_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30173_3_lut (.I0(n35811), .I1(n86), .I2(n29_adj_4343), .I3(GND_net), 
            .O(n35812));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30173_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28721_4_lut (.I0(n33_adj_4346), .I1(n31_adj_4345), .I2(n29_adj_4343), 
            .I3(n34364), .O(n34358));
    defparam i28721_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3172_19 (.CI(n25262), .I0(n2449), .I1(n83), .CO(n25263));
    SB_LUT4 add_3172_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n25261), 
            .O(n6756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_18 (.CI(n25261), .I0(n2450), .I1(n84), .CO(n25262));
    SB_LUT4 add_3172_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n25260), 
            .O(n6757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_17 (.CI(n25260), .I0(n2451), .I1(n85), .CO(n25261));
    SB_LUT4 add_3172_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n25259), 
            .O(n6758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_16 (.CI(n25259), .I0(n2452), .I1(n86), .CO(n25260));
    SB_LUT4 add_3172_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n25258), 
            .O(n6759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_15 (.CI(n25258), .I0(n2453), .I1(n87), .CO(n25259));
    SB_LUT4 add_3172_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n25257), 
            .O(n6760)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1268_3_lut_3_lut (.I0(n1886), .I1(n6652), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30436_4_lut (.I0(n30_adj_4344), .I1(n10_adj_4330), .I2(n35_adj_4347), 
            .I3(n34356), .O(n36075));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30436_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_43_i1265_3_lut_3_lut (.I0(n1886), .I1(n6649), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3172_14 (.CI(n25257), .I0(n2454), .I1(n88), .CO(n25258));
    SB_LUT4 i22_3_lut (.I0(bit_ctr[18]), .I1(n34315), .I2(n4404), .I3(GND_net), 
            .O(n29121));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1559 (.I0(bit_ctr[19]), .I1(n34316), .I2(n4404), 
            .I3(GND_net), .O(n29123));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1559.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1560 (.I0(bit_ctr[20]), .I1(n34317), .I2(n4404), 
            .I3(GND_net), .O(n29125));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1560.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1561 (.I0(bit_ctr[21]), .I1(n34318), .I2(n4404), 
            .I3(GND_net), .O(n29127));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1561.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1562 (.I0(bit_ctr[22]), .I1(n34319), .I2(n4404), 
            .I3(GND_net), .O(n29129));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1562.LUT_INIT = 16'hacac;
    SB_LUT4 i30149_3_lut (.I0(n35812), .I1(n85), .I2(n31_adj_4345), .I3(GND_net), 
            .O(n35788));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30149_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30510_4_lut (.I0(n35788), .I1(n36075), .I2(n35_adj_4347), 
            .I3(n34358), .O(n36149));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30510_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30511_3_lut (.I0(n36149), .I1(n82), .I2(n37_adj_4348), .I3(GND_net), 
            .O(n36150));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30511_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30476_3_lut (.I0(n36150), .I1(n81), .I2(n39_adj_4349), .I3(GND_net), 
            .O(n36115));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30476_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3172_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n25256), 
            .O(n6761)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_13 (.CI(n25256), .I0(n2455), .I1(n89), .CO(n25257));
    SB_LUT4 add_3172_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n25255), 
            .O(n6762)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28704_4_lut (.I0(n43_adj_4352), .I1(n41_adj_4351), .I2(n39_adj_4349), 
            .I3(n36018), .O(n34341));
    defparam i28704_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3172_12 (.CI(n25255), .I0(n2456), .I1(n90), .CO(n25256));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_164[6]), 
            .I2(n19_adj_3990), .I3(n24856), .O(displacement_23__N_40[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3172_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n25254), 
            .O(n6763)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30402_4_lut (.I0(n35786), .I1(n35791), .I2(n45_adj_4353), 
            .I3(n34995), .O(n36041));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30402_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_43_i1266_3_lut_3_lut (.I0(n1886), .I1(n6650), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30470_3_lut (.I0(n36115), .I1(n80), .I2(n41_adj_4351), .I3(GND_net), 
            .O(n40_adj_4350));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30470_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1807_3_lut (.I0(n2699), .I1(n6822), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30404_4_lut (.I0(n40_adj_4350), .I1(n36041), .I2(n45_adj_4353), 
            .I3(n34341), .O(n36043));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30404_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30405_3_lut (.I0(n36043), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30405_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3172_11 (.CI(n25254), .I0(n2457), .I1(n91), .CO(n25255));
    SB_LUT4 add_3172_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n25253), 
            .O(n6764)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_10 (.CI(n25253), .I0(n2458), .I1(n92), .CO(n25254));
    SB_LUT4 div_43_i1264_3_lut_3_lut (.I0(n1886), .I1(n6648), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3172_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n25252), 
            .O(n6765)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_9 (.CI(n25252), .I0(n2459), .I1(n93), .CO(n25253));
    SB_LUT4 add_3172_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n25251), 
            .O(n6766)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n24856), .I0(displacement_23__N_164[6]), 
            .I1(n19_adj_3990), .CO(n24857));
    SB_CARRY add_3172_8 (.CI(n25251), .I0(n2460), .I1(n94), .CO(n25252));
    SB_LUT4 add_3172_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n25250), 
            .O(n6767)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_7 (.CI(n25250), .I0(n2461), .I1(n95), .CO(n25251));
    SB_LUT4 add_3172_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n25249), 
            .O(n6768)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_6 (.CI(n25249), .I0(n2462), .I1(n96), .CO(n25250));
    SB_LUT4 add_3172_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n25248), 
            .O(n6769)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_5 (.CI(n25248), .I0(n2463), .I1(n97), .CO(n25249));
    SB_LUT4 add_3172_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n25247), 
            .O(n6770)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_4 (.CI(n25247), .I0(n2464), .I1(n98), .CO(n25248));
    SB_LUT4 add_3172_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n25246), 
            .O(n6771)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_3 (.CI(n25246), .I0(n2465), .I1(n99), .CO(n25247));
    SB_LUT4 add_3172_2_lut (.I0(GND_net), .I1(n387), .I2(n558), .I3(VCC_net), 
            .O(n6772)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_2 (.CI(VCC_net), .I0(n387), .I1(n558), .CO(n25246));
    SB_LUT4 add_3171_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n25245), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3171_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n25244), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_19 (.CI(n25244), .I0(n2358), .I1(n83), .CO(n25245));
    SB_LUT4 add_3171_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n25243), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_18 (.CI(n25243), .I0(n2359), .I1(n84), .CO(n25244));
    SB_LUT4 div_43_i1271_3_lut_3_lut (.I0(n1886), .I1(n6655), .I2(n381), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1263_3_lut_3_lut (.I0(n1886), .I1(n6647), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1777_i43_2_lut (.I0(n2701), .I1(n80), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4324));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1262_3_lut_3_lut (.I0(n1886), .I1(n6646), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1777_i41_2_lut (.I0(n2702), .I1(n81), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4322));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1777_i39_2_lut (.I0(n2703), .I1(n82), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4321));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_164[5]), 
            .I2(n20_adj_3991), .I3(n24855), .O(displacement_23__N_40[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3171_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n25242), 
            .O(n6735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n24855), .I0(displacement_23__N_164[5]), 
            .I1(n20_adj_3991), .CO(n24856));
    SB_LUT4 div_43_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_3945), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3171_17 (.CI(n25242), .I0(n2360), .I1(n85), .CO(n25243));
    SB_LUT4 add_3171_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n25241), 
            .O(n6736)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4316));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4318));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3171_16 (.CI(n25241), .I0(n2361), .I1(n86), .CO(n25242));
    SB_LUT4 add_3171_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n25240), 
            .O(n6737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4313));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4314));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4311));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4312));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_40[21]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_40[20]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_40[19]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_40[18]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_40[17]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_40[16]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_40[15]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_40[14]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_40[13]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_40[12]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_40[11]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_40[10]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_40[9]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_40[8]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_40[7]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_40[6]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_40[5]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_40[4]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_40[3]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_40[2]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_40[1]));   // verilog/TinyFPGA_B.v(205[10] 207[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[22]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[21]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[20]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[19]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[18]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[17]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[16]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[15]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[14]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[13]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[12]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[11]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[10]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[9]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[8]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[7]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[6]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[5]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[4]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[3]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[2]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[1]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_DFF blue_1128__i0 (.Q(blue[0]), .C(LED_c), .D(n45));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_LUT4 i12432_4_lut (.I0(n16687), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n16600), .O(n16819));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12432_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_43_i1261_3_lut_3_lut (.I0(n1886), .I1(n6645), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12429_4_lut (.I0(n16687), .I1(r_Bit_Index[2]), .I2(n4573), 
            .I3(n16600), .O(n16816));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12429_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_43_i1340_3_lut_3_lut (.I0(n1991), .I1(n6671), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1563 (.I0(bit_ctr[23]), .I1(n34320), .I2(n4404), 
            .I3(GND_net), .O(n29131));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1563.LUT_INIT = 16'hacac;
    SB_CARRY add_3171_15 (.CI(n25240), .I0(n2362), .I1(n87), .CO(n25241));
    SB_LUT4 add_3171_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n25239), 
            .O(n6738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_164[4]), 
            .I2(n21_adj_3992), .I3(n24854), .O(displacement_23__N_40[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n24854), .I0(displacement_23__N_164[4]), 
            .I1(n21_adj_3992), .CO(n24855));
    SB_LUT4 div_43_i1332_3_lut_3_lut (.I0(n1991), .I1(n6663), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1331_3_lut_3_lut (.I0(n1991), .I1(n6662), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i638_3_lut_3_lut (.I0(n938), .I1(n6554), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4302));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1330_3_lut_3_lut (.I0(n1991), .I1(n6661), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1564 (.I0(bit_ctr[1]), .I1(n34321), .I2(n4404), 
            .I3(GND_net), .O(n29133));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1564.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1565 (.I0(bit_ctr[24]), .I1(n34322), .I2(n4404), 
            .I3(GND_net), .O(n29135));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1565.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1566 (.I0(bit_ctr[25]), .I1(n34323), .I2(n4404), 
            .I3(GND_net), .O(n29137));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1566.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_164[3]), 
            .I2(n22_adj_3993), .I3(n24853), .O(displacement_23__N_40[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n24853), .I0(displacement_23__N_164[3]), 
            .I1(n22_adj_3993), .CO(n24854));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_164[2]), 
            .I2(n23_adj_3994), .I3(n24852), .O(displacement_23__N_40[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n24852), .I0(displacement_23__N_164[2]), 
            .I1(n23_adj_3994), .CO(n24853));
    SB_CARRY add_3171_14 (.CI(n25239), .I0(n2363), .I1(n88), .CO(n25240));
    SB_LUT4 div_43_i1328_3_lut_3_lut (.I0(n1991), .I1(n6659), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3171_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n25238), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_164[1]), 
            .I2(n24_adj_3995), .I3(n24851), .O(displacement_23__N_40[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_13 (.CI(n25238), .I0(n2364), .I1(n89), .CO(n25239));
    SB_LUT4 add_3171_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n25237), 
            .O(n6740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n24851), .I0(displacement_23__N_164[1]), 
            .I1(n24_adj_3995), .CO(n24852));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_164[0]), 
            .I2(n25_adj_3996), .I3(VCC_net), .O(displacement_23__N_40[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_12 (.CI(n25237), .I0(n2365), .I1(n90), .CO(n25238));
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_164[0]), 
            .I1(n25_adj_3996), .CO(n24851));
    SB_LUT4 add_3171_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n25236), 
            .O(n6741)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_11 (.CI(n25236), .I0(n2366), .I1(n91), .CO(n25237));
    SB_LUT4 div_43_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4320));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3171_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n25235), 
            .O(n6742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_10 (.CI(n25235), .I0(n2367), .I1(n92), .CO(n25236));
    SB_LUT4 add_3171_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n25234), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1329_3_lut_3_lut (.I0(n1991), .I1(n6660), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3171_9 (.CI(n25234), .I0(n2368), .I1(n93), .CO(n25235));
    SB_LUT4 add_3171_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n25233), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_8 (.CI(n25233), .I0(n2369), .I1(n94), .CO(n25234));
    SB_LUT4 add_3171_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n25232), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_7 (.CI(n25232), .I0(n2370), .I1(n95), .CO(n25233));
    SB_LUT4 add_3171_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n25231), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_6 (.CI(n25231), .I0(n2371), .I1(n96), .CO(n25232));
    SB_LUT4 add_3171_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n25230), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_5 (.CI(n25230), .I0(n2372), .I1(n97), .CO(n25231));
    SB_LUT4 add_3171_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n25229), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_4 (.CI(n25229), .I0(n2373), .I1(n98), .CO(n25230));
    SB_LUT4 add_3171_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n25228), 
            .O(n6749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_3 (.CI(n25228), .I0(n2374), .I1(n99), .CO(n25229));
    SB_LUT4 div_43_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4304));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3171_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4310));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3171_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n25228));
    SB_LUT4 div_43_i1327_3_lut_3_lut (.I0(n1991), .I1(n6658), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3170_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n25227), 
            .O(n6712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n25226), 
            .O(n6713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_18 (.CI(n25226), .I0(n2265), .I1(n84), .CO(n25227));
    SB_LUT4 add_3170_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n25225), 
            .O(n6714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_17 (.CI(n25225), .I0(n2266), .I1(n85), .CO(n25226));
    SB_LUT4 div_43_i1338_3_lut_3_lut (.I0(n1991), .I1(n6669), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3170_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n25224), 
            .O(n6715)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_16 (.CI(n25224), .I0(n2267), .I1(n86), .CO(n25225));
    SB_LUT4 add_3170_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n25223), 
            .O(n6716)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4319));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3170_15 (.CI(n25223), .I0(n2268), .I1(n87), .CO(n25224));
    SB_LUT4 add_3170_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n25222), 
            .O(n6717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4306));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3170_14 (.CI(n25222), .I0(n2269), .I1(n88), .CO(n25223));
    SB_LUT4 add_3170_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n25221), 
            .O(n6718)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_13 (.CI(n25221), .I0(n2270), .I1(n89), .CO(n25222));
    SB_LUT4 div_43_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4308));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3170_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n25220), 
            .O(n6719)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4309));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3170_12 (.CI(n25220), .I0(n2271), .I1(n90), .CO(n25221));
    SB_LUT4 i13033_3_lut (.I0(encoder0_position[1]), .I1(n2644), .I2(count_enable), 
            .I3(GND_net), .O(n17420));   // quad.v(35[10] 41[6])
    defparam i13033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3170_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n25219), 
            .O(n6720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4315));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13034_3_lut (.I0(encoder0_position[2]), .I1(n2643), .I2(count_enable), 
            .I3(GND_net), .O(n17421));   // quad.v(35[10] 41[6])
    defparam i13034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13035_3_lut (.I0(encoder0_position[3]), .I1(n2642), .I2(count_enable), 
            .I3(GND_net), .O(n17422));   // quad.v(35[10] 41[6])
    defparam i13035_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3170_11 (.CI(n25219), .I0(n2272), .I1(n91), .CO(n25220));
    SB_LUT4 add_3170_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n25218), 
            .O(n6721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_10 (.CI(n25218), .I0(n2273), .I1(n92), .CO(n25219));
    SB_LUT4 i13036_3_lut (.I0(encoder0_position[4]), .I1(n2641), .I2(count_enable), 
            .I3(GND_net), .O(n17423));   // quad.v(35[10] 41[6])
    defparam i13036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28806_4_lut (.I0(n29_adj_4315), .I1(n17_adj_4309), .I2(n15_adj_4308), 
            .I3(n13_adj_4306), .O(n34443));
    defparam i28806_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13037_3_lut (.I0(encoder0_position[5]), .I1(n2640), .I2(count_enable), 
            .I3(GND_net), .O(n17424));   // quad.v(35[10] 41[6])
    defparam i13037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3935));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_25_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_25_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_25_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_25_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_25_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1339_3_lut_3_lut (.I0(n1991), .I1(n6670), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13038_3_lut (.I0(encoder0_position[6]), .I1(n2639), .I2(count_enable), 
            .I3(GND_net), .O(n17425));   // quad.v(35[10] 41[6])
    defparam i13038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1337_3_lut_3_lut (.I0(n1991), .I1(n6668), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13039_3_lut (.I0(encoder0_position[7]), .I1(n2638), .I2(count_enable), 
            .I3(GND_net), .O(n17426));   // quad.v(35[10] 41[6])
    defparam i13039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13040_3_lut (.I0(encoder0_position[8]), .I1(n2637), .I2(count_enable), 
            .I3(GND_net), .O(n17427));   // quad.v(35[10] 41[6])
    defparam i13040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1777_i32_3_lut (.I0(n14_adj_4307), .I1(n83), 
            .I2(n37_adj_4320), .I3(GND_net), .O(n32_adj_4317));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13041_3_lut (.I0(encoder0_position[9]), .I1(n2636), .I2(count_enable), 
            .I3(GND_net), .O(n17428));   // quad.v(35[10] 41[6])
    defparam i13041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29396_4_lut (.I0(n11_adj_4304), .I1(n9_adj_4302), .I2(n2719), 
            .I3(n98), .O(n35034));
    defparam i29396_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i13042_3_lut (.I0(encoder0_position[10]), .I1(n2635), .I2(count_enable), 
            .I3(GND_net), .O(n17429));   // quad.v(35[10] 41[6])
    defparam i13042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29804_4_lut (.I0(n17_adj_4309), .I1(n15_adj_4308), .I2(n13_adj_4306), 
            .I3(n35034), .O(n35443));
    defparam i29804_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i13043_3_lut (.I0(encoder0_position[11]), .I1(n2634), .I2(count_enable), 
            .I3(GND_net), .O(n17430));   // quad.v(35[10] 41[6])
    defparam i13043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29798_4_lut (.I0(n23_adj_4312), .I1(n21_adj_4311), .I2(n19_adj_4310), 
            .I3(n35443), .O(n35437));
    defparam i29798_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28706_4_lut (.I0(n29_adj_4315), .I1(n27_adj_4314), .I2(n25_adj_4313), 
            .I3(n35437), .O(n34343));
    defparam i28706_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3170_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n25217), 
            .O(n6722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13044_3_lut (.I0(encoder0_position[12]), .I1(n2633), .I2(count_enable), 
            .I3(GND_net), .O(n17431));   // quad.v(35[10] 41[6])
    defparam i13044_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3170_9 (.CI(n25217), .I0(n2274), .I1(n93), .CO(n25218));
    SB_LUT4 i13045_3_lut (.I0(encoder0_position[13]), .I1(n2632), .I2(count_enable), 
            .I3(GND_net), .O(n17432));   // quad.v(35[10] 41[6])
    defparam i13045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29834_4_lut (.I0(n35_adj_4319), .I1(n33_adj_4318), .I2(n31_adj_4316), 
            .I3(n34343), .O(n35473));
    defparam i29834_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13046_3_lut (.I0(encoder0_position[14]), .I1(n2631), .I2(count_enable), 
            .I3(GND_net), .O(n17433));   // quad.v(35[10] 41[6])
    defparam i13046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13047_3_lut (.I0(encoder0_position[15]), .I1(n2630), .I2(count_enable), 
            .I3(GND_net), .O(n17434));   // quad.v(35[10] 41[6])
    defparam i13047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13048_3_lut (.I0(encoder0_position[16]), .I1(n2629), .I2(count_enable), 
            .I3(GND_net), .O(n17435));   // quad.v(35[10] 41[6])
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13049_3_lut (.I0(encoder0_position[17]), .I1(n2628), .I2(count_enable), 
            .I3(GND_net), .O(n17436));   // quad.v(35[10] 41[6])
    defparam i13049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30182_3_lut (.I0(n8_adj_4301), .I1(n90), .I2(n23_adj_4312), 
            .I3(GND_net), .O(n35821));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30182_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13050_3_lut (.I0(encoder0_position[18]), .I1(n2627), .I2(count_enable), 
            .I3(GND_net), .O(n17437));   // quad.v(35[10] 41[6])
    defparam i13050_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i30183_3_lut (.I0(n35821), .I1(n89), .I2(n25_adj_4313), .I3(GND_net), 
            .O(n35822));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30183_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13051_3_lut (.I0(encoder0_position[19]), .I1(n2626), .I2(count_enable), 
            .I3(GND_net), .O(n17438));   // quad.v(35[10] 41[6])
    defparam i13051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29372_4_lut (.I0(n25_adj_4313), .I1(n23_adj_4312), .I2(n21_adj_4311), 
            .I3(n34360), .O(n35010));
    defparam i29372_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_43_i1336_3_lut_3_lut (.I0(n1991), .I1(n6667), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3170_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n25216), 
            .O(n6723)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_8 (.CI(n25216), .I0(n2275), .I1(n94), .CO(n25217));
    SB_LUT4 i13052_3_lut (.I0(encoder0_position[20]), .I1(n2625), .I2(count_enable), 
            .I3(GND_net), .O(n17439));   // quad.v(35[10] 41[6])
    defparam i13052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3170_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n25215), 
            .O(n6724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24_3_lut (.I0(n34288), .I1(bit_ctr[26]), .I2(n4404), .I3(GND_net), 
            .O(n29069));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13053_3_lut (.I0(encoder0_position[21]), .I1(n2624), .I2(count_enable), 
            .I3(GND_net), .O(n17440));   // quad.v(35[10] 41[6])
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3170_7 (.CI(n25215), .I0(n2276), .I1(n95), .CO(n25216));
    SB_LUT4 i30136_3_lut (.I0(n10_adj_4303), .I1(n91), .I2(n21_adj_4311), 
            .I3(GND_net), .O(n35775));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30136_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13054_3_lut (.I0(encoder0_position[22]), .I1(n2623), .I2(count_enable), 
            .I3(GND_net), .O(n17441));   // quad.v(35[10] 41[6])
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30135_3_lut (.I0(n35822), .I1(n88), .I2(n27_adj_4314), .I3(GND_net), 
            .O(n35774));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30135_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4300));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30180_3_lut (.I0(n6_adj_4300), .I1(n87), .I2(n29_adj_4315), 
            .I3(GND_net), .O(n35819));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30180_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3170_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n25214), 
            .O(n6725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_6 (.CI(n25214), .I0(n2277), .I1(n96), .CO(n25215));
    SB_LUT4 add_3170_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n25213), 
            .O(n6726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_5 (.CI(n25213), .I0(n2278), .I1(n97), .CO(n25214));
    SB_LUT4 add_3170_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n25212), 
            .O(n6727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_4 (.CI(n25212), .I0(n2279), .I1(n98), .CO(n25213));
    SB_LUT4 i13055_3_lut (.I0(encoder0_position[23]), .I1(n2622), .I2(count_enable), 
            .I3(GND_net), .O(n17442));   // quad.v(35[10] 41[6])
    defparam i13055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3170_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n25211), 
            .O(n6728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30181_3_lut (.I0(n35819), .I1(n86), .I2(n31_adj_4316), .I3(GND_net), 
            .O(n35820));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30181_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28796_4_lut (.I0(n35_adj_4319), .I1(n33_adj_4318), .I2(n31_adj_4316), 
            .I3(n34443), .O(n34433));
    defparam i28796_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30434_4_lut (.I0(n32_adj_4317), .I1(n12_adj_4305), .I2(n37_adj_4320), 
            .I3(n34425), .O(n36073));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30434_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30139_3_lut (.I0(n35820), .I1(n85), .I2(n33_adj_4318), .I3(GND_net), 
            .O(n35778));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30139_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3170_3 (.CI(n25211), .I0(n2280), .I1(n99), .CO(n25212));
    SB_LUT4 add_3170_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n25211));
    SB_LUT4 add_3169_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n25210), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3169_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n25209), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_17 (.CI(n25209), .I0(n2169), .I1(n85), .CO(n25210));
    SB_LUT4 add_3169_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n25208), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_16 (.CI(n25208), .I0(n2170), .I1(n86), .CO(n25209));
    SB_LUT4 div_43_i1335_3_lut_3_lut (.I0(n1991), .I1(n6666), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30508_4_lut (.I0(n35778), .I1(n36073), .I2(n37_adj_4320), 
            .I3(n34433), .O(n36147));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30508_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30509_3_lut (.I0(n36147), .I1(n82), .I2(n39_adj_4321), .I3(GND_net), 
            .O(n36148));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30509_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30478_3_lut (.I0(n36148), .I1(n81), .I2(n41_adj_4322), .I3(GND_net), 
            .O(n36117));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30478_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3169_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n25207), 
            .O(n6696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_15 (.CI(n25207), .I0(n2171), .I1(n87), .CO(n25208));
    SB_LUT4 add_3169_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n25206), 
            .O(n6697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_14 (.CI(n25206), .I0(n2172), .I1(n88), .CO(n25207));
    SB_LUT4 add_3169_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n25205), 
            .O(n6698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30383_4_lut (.I0(n41_adj_4322), .I1(n39_adj_4321), .I2(n37_adj_4320), 
            .I3(n35473), .O(n36022));
    defparam i30383_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3169_13 (.CI(n25205), .I0(n2173), .I1(n89), .CO(n25206));
    SB_LUT4 add_3169_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n25204), 
            .O(n6699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_12 (.CI(n25204), .I0(n2174), .I1(n90), .CO(n25205));
    SB_LUT4 i30176_4_lut (.I0(n35774), .I1(n35775), .I2(n27_adj_4314), 
            .I3(n35010), .O(n35815));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30176_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3169_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n25203), 
            .O(n6700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_11 (.CI(n25203), .I0(n2175), .I1(n91), .CO(n25204));
    SB_LUT4 add_3169_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n25202), 
            .O(n6701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_10 (.CI(n25202), .I0(n2176), .I1(n92), .CO(n25203));
    SB_LUT4 add_3169_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n25201), 
            .O(n6702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30468_3_lut (.I0(n36117), .I1(n80), .I2(n43_adj_4324), .I3(GND_net), 
            .O(n42_adj_4323));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30468_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3169_9 (.CI(n25201), .I0(n2177), .I1(n93), .CO(n25202));
    SB_LUT4 i30375_4_lut (.I0(n42_adj_4323), .I1(n35815), .I2(n43_adj_4324), 
            .I3(n36022), .O(n36014));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30375_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3169_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n25200), 
            .O(n6703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30376_3_lut (.I0(n36014), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n36015));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30376_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY add_3169_8 (.CI(n25200), .I0(n2178), .I1(n94), .CO(n25201));
    SB_LUT4 add_3169_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n25199), 
            .O(n6704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_7 (.CI(n25199), .I0(n2179), .I1(n95), .CO(n25200));
    SB_LUT4 add_3169_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n25198), 
            .O(n6705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_6 (.CI(n25198), .I0(n2180), .I1(n96), .CO(n25199));
    SB_LUT4 add_3169_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n25197), 
            .O(n6706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_5 (.CI(n25197), .I0(n2181), .I1(n97), .CO(n25198));
    SB_LUT4 add_3169_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n25196), 
            .O(n6707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_4 (.CI(n25196), .I0(n2182), .I1(n98), .CO(n25197));
    SB_LUT4 div_43_i1334_3_lut_3_lut (.I0(n1991), .I1(n6665), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1974_4_lut (.I0(n36015), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1974_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 add_3169_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n25195), 
            .O(n6708)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_3 (.CI(n25195), .I0(n2183), .I1(n99), .CO(n25196));
    SB_LUT4 add_3169_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n25195));
    SB_LUT4 add_3168_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n25194), 
            .O(n6675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1341_3_lut_3_lut (.I0(n1991), .I1(n6672), .I2(n382), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3168_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n25193), 
            .O(n6676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1333_3_lut_3_lut (.I0(n1991), .I1(n6664), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i35_2_lut (.I0(n2624_adj_4000), .I1(n85), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4297));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1722_i39_2_lut (.I0(n2622_adj_3998), .I1(n83), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4299));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_16 (.CI(n25193), .I0(n2070), .I1(n86), .CO(n25194));
    SB_LUT4 div_43_LessThan_1722_i33_2_lut (.I0(n2625_adj_4001), .I1(n86), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4295));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3168_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n25192), 
            .O(n6677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_15 (.CI(n25192), .I0(n2071), .I1(n87), .CO(n25193));
    SB_LUT4 add_3168_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n25191), 
            .O(n6678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_14 (.CI(n25191), .I0(n2072), .I1(n88), .CO(n25192));
    SB_LUT4 add_3168_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n25190), 
            .O(n6679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_13 (.CI(n25190), .I0(n2073), .I1(n89), .CO(n25191));
    SB_LUT4 div_43_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_3946), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1408_3_lut_3_lut (.I0(n2093), .I1(n6689), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i37_2_lut (.I0(n2623_adj_3999), .I1(n84), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4298));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3168_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n25189), 
            .O(n6680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_12 (.CI(n25189), .I0(n2074), .I1(n90), .CO(n25190));
    SB_LUT4 add_3168_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n25188), 
            .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1722_i27_2_lut (.I0(n2628_adj_4004), .I1(n89), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4292));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1722_i29_2_lut (.I0(n2627_adj_4003), .I1(n88), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4293));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_11 (.CI(n25188), .I0(n2075), .I1(n91), .CO(n25189));
    SB_LUT4 div_43_i1397_3_lut_3_lut (.I0(n2093), .I1(n6678), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1401_3_lut_3_lut (.I0(n2093), .I1(n6682), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i11_2_lut (.I0(n2636_adj_4012), .I1(n97), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4280));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1722_i23_2_lut (.I0(n2630_adj_4006), .I1(n91), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4290));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3168_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n25187), 
            .O(n6682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1400_3_lut_3_lut (.I0(n2093), .I1(n6681), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i25_2_lut (.I0(n2629_adj_4005), .I1(n90), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4291));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(n5_adj_4018), .I1(n63_adj_4017), .I2(n2421), 
            .I3(n18493), .O(n6_adj_4360));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'heaaa;
    SB_CARRY add_3168_10 (.CI(n25187), .I0(n2076), .I1(n92), .CO(n25188));
    SB_LUT4 i3_4_lut (.I0(n3761), .I1(n6_adj_4360), .I2(n15501), .I3(n37539), 
            .O(n8_adj_3997));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut.LUT_INIT = 16'hcfce;
    SB_LUT4 i4_4_lut_adj_1568 (.I0(n18493), .I1(n8_adj_3997), .I2(n15494), 
            .I3(n5_adj_4359), .O(n37085));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1568.LUT_INIT = 16'hefcf;
    SB_LUT4 div_43_LessThan_1722_i13_2_lut (.I0(n2635_adj_4011), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4282));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1399_3_lut_3_lut (.I0(n2093), .I1(n6680), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3168_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n25186), 
            .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1396_3_lut_3_lut (.I0(n2093), .I1(n6677), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1395_3_lut_3_lut (.I0(n2093), .I1(n6676), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i15_2_lut (.I0(n2634_adj_4010), .I1(n95), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4284));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_9 (.CI(n25186), .I0(n2077), .I1(n93), .CO(n25187));
    SB_LUT4 div_43_i1398_3_lut_3_lut (.I0(n2093), .I1(n6679), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1394_3_lut_3_lut (.I0(n2093), .I1(n6675), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1405_3_lut_3_lut (.I0(n2093), .I1(n6686), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1404_3_lut_3_lut (.I0(n2093), .I1(n6685), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3168_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n25185), 
            .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1722_i17_2_lut (.I0(n2633_adj_4009), .I1(n94), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4286));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13057_3_lut (.I0(encoder1_position[1]), .I1(n2594), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17444));   // quad.v(35[10] 41[6])
    defparam i13057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13058_3_lut (.I0(encoder1_position[2]), .I1(n2593), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17445));   // quad.v(35[10] 41[6])
    defparam i13058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13059_3_lut (.I0(encoder1_position[3]), .I1(n2592), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17446));   // quad.v(35[10] 41[6])
    defparam i13059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13060_3_lut (.I0(encoder1_position[4]), .I1(n2591), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17447));   // quad.v(35[10] 41[6])
    defparam i13060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13061_3_lut (.I0(encoder1_position[5]), .I1(n2590), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17448));   // quad.v(35[10] 41[6])
    defparam i13061_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3168_8 (.CI(n25185), .I0(n2078), .I1(n94), .CO(n25186));
    SB_LUT4 i13062_3_lut (.I0(encoder1_position[6]), .I1(n2589), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17449));   // quad.v(35[10] 41[6])
    defparam i13062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(encoder1_position[7]), .I1(n2588), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17450));   // quad.v(35[10] 41[6])
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13064_3_lut (.I0(encoder1_position[8]), .I1(n2587), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17451));   // quad.v(35[10] 41[6])
    defparam i13064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3168_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n25184), 
            .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_7 (.CI(n25184), .I0(n2079), .I1(n95), .CO(n25185));
    SB_LUT4 add_3168_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n25183), 
            .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13065_3_lut (.I0(encoder1_position[9]), .I1(n2586), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17452));   // quad.v(35[10] 41[6])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1722_i19_2_lut (.I0(n2632_adj_4008), .I1(n93), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4287));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1407_3_lut_3_lut (.I0(n2093), .I1(n6688), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1722_i31_2_lut (.I0(n2626_adj_4002), .I1(n87), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4294));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_6 (.CI(n25183), .I0(n2080), .I1(n96), .CO(n25184));
    SB_LUT4 add_3168_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n25182), 
            .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13066_3_lut (.I0(encoder1_position[10]), .I1(n2585), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17453));   // quad.v(35[10] 41[6])
    defparam i13066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13067_3_lut (.I0(encoder1_position[11]), .I1(n2584), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17454));   // quad.v(35[10] 41[6])
    defparam i13067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13068_3_lut (.I0(encoder1_position[12]), .I1(n2583), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17455));   // quad.v(35[10] 41[6])
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13069_3_lut (.I0(encoder1_position[13]), .I1(n2582), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17456));   // quad.v(35[10] 41[6])
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13070_3_lut (.I0(encoder1_position[14]), .I1(n2581), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17457));   // quad.v(35[10] 41[6])
    defparam i13070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13071_3_lut (.I0(encoder1_position[15]), .I1(n2580), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17458));   // quad.v(35[10] 41[6])
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1722_i21_2_lut (.I0(n2631_adj_4007), .I1(n92), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4289));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1724_1_lut (.I0(n2642_adj_4015), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643_adj_4016));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1406_3_lut_3_lut (.I0(n2093), .I1(n6687), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i28768_4_lut (.I0(n31_adj_4294), .I1(n19_adj_4287), .I2(n17_adj_4286), 
            .I3(n15_adj_4284), .O(n34405));
    defparam i28768_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13072_3_lut (.I0(encoder1_position[16]), .I1(n2579), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17459));   // quad.v(35[10] 41[6])
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29444_4_lut (.I0(n13_adj_4282), .I1(n11_adj_4280), .I2(n2637_adj_4013), 
            .I3(n98), .O(n35082));
    defparam i29444_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i13073_3_lut (.I0(encoder1_position[17]), .I1(n2578), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17460));   // quad.v(35[10] 41[6])
    defparam i13073_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3168_5 (.CI(n25182), .I0(n2081), .I1(n97), .CO(n25183));
    SB_LUT4 i13074_3_lut (.I0(encoder1_position[18]), .I1(n2577), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17461));   // quad.v(35[10] 41[6])
    defparam i13074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13075_3_lut (.I0(encoder1_position[19]), .I1(n2576), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17462));   // quad.v(35[10] 41[6])
    defparam i13075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13076_3_lut (.I0(encoder1_position[20]), .I1(n2575), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17463));   // quad.v(35[10] 41[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13077_3_lut (.I0(encoder1_position[21]), .I1(n2574), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17464));   // quad.v(35[10] 41[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13078_3_lut (.I0(encoder1_position[22]), .I1(n2573), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17465));   // quad.v(35[10] 41[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3168_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n25181), 
            .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1409_3_lut_3_lut (.I0(n2093), .I1(n6690), .I2(n383), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3168_4 (.CI(n25181), .I0(n2082), .I1(n98), .CO(n25182));
    SB_LUT4 add_3168_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n25180), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_3 (.CI(n25180), .I0(n2083), .I1(n99), .CO(n25181));
    SB_LUT4 add_3168_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13079_3_lut (.I0(encoder1_position[23]), .I1(n2572), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n17466));   // quad.v(35[10] 41[6])
    defparam i13079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13080_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n31114), 
            .I3(GND_net), .O(n17467));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13080_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3168_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n25180));
    SB_LUT4 i24_3_lut_adj_1569 (.I0(n34291), .I1(bit_ctr[8]), .I2(n4404), 
            .I3(GND_net), .O(n29075));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1569.LUT_INIT = 16'hcaca;
    SB_LUT4 i29828_4_lut (.I0(n19_adj_4287), .I1(n17_adj_4286), .I2(n15_adj_4284), 
            .I3(n35082), .O(n35467));
    defparam i29828_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24_3_lut_adj_1570 (.I0(n34290), .I1(bit_ctr[7]), .I2(n4404), 
            .I3(GND_net), .O(n29073));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1570.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1571 (.I0(n34289), .I1(bit_ctr[6]), .I2(n4404), 
            .I3(GND_net), .O(n29071));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1571.LUT_INIT = 16'hcaca;
    SB_LUT4 i13092_3_lut (.I0(quadA_debounced_adj_3970), .I1(reg_B_adj_4409[1]), 
            .I2(n31841), .I3(GND_net), .O(n17479));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1403_3_lut_3_lut (.I0(n2093), .I1(n6684), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1402_3_lut_3_lut (.I0(n2093), .I1(n6683), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1572 (.I0(bit_ctr[30]), .I1(n34295), .I2(n4404), 
            .I3(GND_net), .O(n29083));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1572.LUT_INIT = 16'hacac;
    SB_LUT4 i13094_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n925), .I3(GND_net), .O(n17481));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13095_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n925), .I3(GND_net), .O(n17482));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13096_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n925), .I3(GND_net), .O(n17483));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13097_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n925), .I3(GND_net), .O(n17484));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13098_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n925), .I3(GND_net), .O(n17485));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13099_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n925), .I3(GND_net), .O(n17486));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29824_4_lut (.I0(n25_adj_4291), .I1(n23_adj_4290), .I2(n21_adj_4289), 
            .I3(n35467), .O(n35463));
    defparam i29824_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i13100_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n925), .I3(GND_net), .O(n17487));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1573 (.I0(bit_ctr[9]), .I1(n34296), .I2(n4404), 
            .I3(GND_net), .O(n29085));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1573.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1574 (.I0(bit_ctr[31]), .I1(n34301), .I2(n4404), 
            .I3(GND_net), .O(n29089));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1574.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1575 (.I0(bit_ctr[2]), .I1(n34302), .I2(n4404), 
            .I3(GND_net), .O(n29091));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1575.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1576 (.I0(bit_ctr[3]), .I1(n34303), .I2(n4404), 
            .I3(GND_net), .O(n29093));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1576.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1577 (.I0(bit_ctr[4]), .I1(n34304), .I2(n4404), 
            .I3(GND_net), .O(n29095));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1577.LUT_INIT = 16'hacac;
    SB_LUT4 i28774_4_lut (.I0(n31_adj_4294), .I1(n29_adj_4293), .I2(n27_adj_4292), 
            .I3(n35463), .O(n34411));
    defparam i28774_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i22_3_lut_adj_1578 (.I0(bit_ctr[0]), .I1(n34305), .I2(n4404), 
            .I3(GND_net), .O(n29097));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1578.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638_adj_4014), 
            .I3(n558), .O(n8_adj_4278));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_i1471_3_lut_3_lut (.I0(n2192), .I1(n6705), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1579 (.I0(bit_ctr[5]), .I1(n34306), .I2(n4404), 
            .I3(GND_net), .O(n29103));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1579.LUT_INIT = 16'hacac;
    SB_LUT4 i30186_3_lut (.I0(n8_adj_4278), .I1(n87), .I2(n31_adj_4294), 
            .I3(GND_net), .O(n35825));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30186_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30187_3_lut (.I0(n35825), .I1(n86), .I2(n33_adj_4295), .I3(GND_net), 
            .O(n35826));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30187_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1459_3_lut_3_lut (.I0(n2192), .I1(n6693), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1580 (.I0(bit_ctr[10]), .I1(n34307), .I2(n4404), 
            .I3(GND_net), .O(n29105));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1580.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1581 (.I0(bit_ctr[11]), .I1(n34308), .I2(n4404), 
            .I3(GND_net), .O(n29107));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1581.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1582 (.I0(bit_ctr[12]), .I1(n34309), .I2(n4404), 
            .I3(GND_net), .O(n29109));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1582.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1583 (.I0(bit_ctr[13]), .I1(n34310), .I2(n4404), 
            .I3(GND_net), .O(n29111));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1583.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1722_i34_3_lut (.I0(n16_adj_4285), .I1(n83), 
            .I2(n39_adj_4299), .I3(GND_net), .O(n34_adj_4296));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28758_4_lut (.I0(n37_adj_4298), .I1(n35_adj_4297), .I2(n33_adj_4295), 
            .I3(n34405), .O(n34395));
    defparam i28758_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i22_3_lut_adj_1584 (.I0(bit_ctr[14]), .I1(n34311), .I2(n4404), 
            .I3(GND_net), .O(n29113));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1584.LUT_INIT = 16'hacac;
    SB_LUT4 i30432_4_lut (.I0(n34_adj_4296), .I1(n14_adj_4283), .I2(n39_adj_4299), 
            .I3(n34389), .O(n36071));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30432_4_lut.LUT_INIT = 16'haaac;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i22_3_lut_adj_1585 (.I0(bit_ctr[15]), .I1(n34312), .I2(n4404), 
            .I3(GND_net), .O(n29115));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1585.LUT_INIT = 16'hacac;
    SB_LUT4 add_3167_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n25158), 
            .O(n6658)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n25157), 
            .O(n6659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_15 (.CI(n25157), .I0(n1968), .I1(n87), .CO(n25158));
    SB_LUT4 div_43_i1470_3_lut_3_lut (.I0(n2192), .I1(n6704), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1467_3_lut_3_lut (.I0(n2192), .I1(n6701), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3167_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n25156), 
            .O(n6660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_14 (.CI(n25156), .I0(n1969), .I1(n88), .CO(n25157));
    SB_LUT4 add_3167_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n25155), 
            .O(n6661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_13 (.CI(n25155), .I0(n1970), .I1(n89), .CO(n25156));
    SB_LUT4 div_43_i1465_3_lut_3_lut (.I0(n2192), .I1(n6699), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3167_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n25154), 
            .O(n6662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_12 (.CI(n25154), .I0(n1971), .I1(n90), .CO(n25155));
    SB_LUT4 add_3167_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n25153), 
            .O(n6663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_11 (.CI(n25153), .I0(n1972), .I1(n91), .CO(n25154));
    SB_LUT4 add_3167_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n25152), 
            .O(n6664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_10 (.CI(n25152), .I0(n1973), .I1(n92), .CO(n25153));
    SB_LUT4 add_3167_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n25151), 
            .O(n6665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_9 (.CI(n25151), .I0(n1974), .I1(n93), .CO(n25152));
    SB_LUT4 add_3167_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n25150), 
            .O(n6666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_8 (.CI(n25150), .I0(n1975), .I1(n94), .CO(n25151));
    SB_LUT4 add_3167_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n25149), 
            .O(n6667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30127_3_lut (.I0(n35826), .I1(n85), .I2(n35_adj_4297), .I3(GND_net), 
            .O(n35766));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30127_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1475_3_lut_3_lut (.I0(n2192), .I1(n6709), .I2(n384), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30188_3_lut (.I0(n10_adj_4279), .I1(n90), .I2(n25_adj_4291), 
            .I3(GND_net), .O(n35827));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30188_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3167_7 (.CI(n25149), .I0(n1976), .I1(n95), .CO(n25150));
    SB_LUT4 add_3167_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n25148), 
            .O(n6668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_6 (.CI(n25148), .I0(n1977), .I1(n96), .CO(n25149));
    SB_LUT4 add_3167_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n25147), 
            .O(n6669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1586 (.I0(bit_ctr[16]), .I1(n34313), .I2(n4404), 
            .I3(GND_net), .O(n29117));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1586.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1463_3_lut_3_lut (.I0(n2192), .I1(n6697), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3167_5 (.CI(n25147), .I0(n1978), .I1(n97), .CO(n25148));
    SB_LUT4 i30189_3_lut (.I0(n35827), .I1(n89), .I2(n27_adj_4292), .I3(GND_net), 
            .O(n35828));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30189_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29430_4_lut (.I0(n27_adj_4292), .I1(n25_adj_4291), .I2(n23_adj_4290), 
            .I3(n34421), .O(n35068));
    defparam i29430_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_43_LessThan_1722_i20_3_lut (.I0(n12_adj_4281), .I1(n91), 
            .I2(n23_adj_4290), .I3(GND_net), .O(n20_adj_4288));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30125_3_lut (.I0(n35828), .I1(n88), .I2(n29_adj_4293), .I3(GND_net), 
            .O(n35764));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30125_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i22_3_lut_adj_1587 (.I0(bit_ctr[17]), .I1(n34314), .I2(n4404), 
            .I3(GND_net), .O(n29119));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1587.LUT_INIT = 16'hacac;
    SB_LUT4 i30011_4_lut (.I0(n37_adj_4298), .I1(n35_adj_4297), .I2(n33_adj_4295), 
            .I3(n34411), .O(n35650));
    defparam i30011_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_43_i1462_3_lut_3_lut (.I0(n2192), .I1(n6696), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3167_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n25146), 
            .O(n6670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_4 (.CI(n25146), .I0(n1979), .I1(n98), .CO(n25147));
    SB_LUT4 add_3167_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n25145), 
            .O(n6671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_i1461_3_lut_3_lut (.I0(n2192), .I1(n6695), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1464_3_lut_3_lut (.I0(n2192), .I1(n6698), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3167_3 (.CI(n25145), .I0(n1980), .I1(n99), .CO(n25146));
    SB_LUT4 add_3167_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n25145));
    SB_LUT4 add_3166_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n25144), 
            .O(n6642)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3166_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n25143), 
            .O(n6643)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30506_4_lut (.I0(n35766), .I1(n36071), .I2(n39_adj_4299), 
            .I3(n34395), .O(n36145));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30506_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3166_14 (.CI(n25143), .I0(n1863), .I1(n88), .CO(n25144));
    SB_LUT4 add_3166_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n25142), 
            .O(n6644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_13 (.CI(n25142), .I0(n1864), .I1(n89), .CO(n25143));
    SB_LUT4 add_3166_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n25141), 
            .O(n6645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30130_4_lut (.I0(n35764), .I1(n20_adj_4288), .I2(n29_adj_4293), 
            .I3(n35068), .O(n35769));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30130_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3166_12 (.CI(n25141), .I0(n1865), .I1(n90), .CO(n25142));
    SB_LUT4 i30520_4_lut (.I0(n35769), .I1(n36145), .I2(n39_adj_4299), 
            .I3(n35650), .O(n36159));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30520_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30521_3_lut (.I0(n36159), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n36160));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30521_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3166_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n25140), 
            .O(n6646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_11 (.CI(n25140), .I0(n1866), .I1(n91), .CO(n25141));
    SB_LUT4 i30515_3_lut (.I0(n36160), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n36154));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30515_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3166_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n25139), 
            .O(n6647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_10 (.CI(n25139), .I0(n1867), .I1(n92), .CO(n25140));
    SB_LUT4 i30132_3_lut (.I0(n36154), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n35771));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30132_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3166_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n25138), 
            .O(n6648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(n35771), .I1(n15490), .I2(n79), .I3(n2618), 
            .O(n2642_adj_4015));
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_i1460_3_lut_3_lut (.I0(n2192), .I1(n6694), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3166_9 (.CI(n25138), .I0(n1868), .I1(n93), .CO(n25139));
    SB_LUT4 add_3166_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n25137), 
            .O(n6649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_8 (.CI(n25137), .I0(n1869), .I1(n94), .CO(n25138));
    SB_LUT4 add_3166_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n25136), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_7 (.CI(n25136), .I0(n1870), .I1(n95), .CO(n25137));
    SB_LUT4 div_43_i1474_3_lut_3_lut (.I0(n2192), .I1(n6708), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3166_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n25135), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_6 (.CI(n25135), .I0(n1871), .I1(n96), .CO(n25136));
    SB_LUT4 add_3166_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n25134), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_5 (.CI(n25134), .I0(n1872), .I1(n97), .CO(n25135));
    SB_LUT4 add_3166_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n25133), 
            .O(n6653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4275));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1472_3_lut_3_lut (.I0(n2192), .I1(n6706), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4277));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3166_4 (.CI(n25133), .I0(n1873), .I1(n98), .CO(n25134));
    SB_LUT4 div_43_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4273));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3166_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n25132), 
            .O(n6654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_3 (.CI(n25132), .I0(n1874), .I1(n99), .CO(n25133));
    SB_LUT4 add_3166_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6655)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n25132));
    SB_LUT4 add_3165_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n25131), 
            .O(n6627)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3165_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n25130), 
            .O(n6628)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_13 (.CI(n25130), .I0(n1755), .I1(n89), .CO(n25131));
    SB_LUT4 add_3165_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n25129), 
            .O(n6629)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_12 (.CI(n25129), .I0(n1756), .I1(n90), .CO(n25130));
    SB_LUT4 add_3165_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n25128), 
            .O(n6630)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_11 (.CI(n25128), .I0(n1757), .I1(n91), .CO(n25129));
    SB_LUT4 add_3165_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n25127), 
            .O(n6631)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_3947), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3165_10 (.CI(n25127), .I0(n1758), .I1(n92), .CO(n25128));
    SB_LUT4 add_3165_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n25126), 
            .O(n6632)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_9 (.CI(n25126), .I0(n1759), .I1(n93), .CO(n25127));
    SB_LUT4 add_3165_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n25125), 
            .O(n6633)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_8 (.CI(n25125), .I0(n1760), .I1(n94), .CO(n25126));
    SB_LUT4 add_3165_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n25124), 
            .O(n6634)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_7 (.CI(n25124), .I0(n1761), .I1(n95), .CO(n25125));
    SB_LUT4 add_3165_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n25123), 
            .O(n6635)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_6 (.CI(n25123), .I0(n1762), .I1(n96), .CO(n25124));
    SB_LUT4 add_3165_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n25122), 
            .O(n6636)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_5 (.CI(n25122), .I0(n1763), .I1(n97), .CO(n25123));
    SB_LUT4 add_3165_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n25121), 
            .O(n6637)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_4 (.CI(n25121), .I0(n1764), .I1(n98), .CO(n25122));
    SB_LUT4 div_43_i1473_3_lut_3_lut (.I0(n2192), .I1(n6707), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4276));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3165_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n25120), 
            .O(n6638)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_3 (.CI(n25120), .I0(n1765), .I1(n99), .CO(n25121));
    SB_LUT4 add_3165_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6639)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n25120));
    SB_LUT4 div_43_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4270));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1469_3_lut_3_lut (.I0(n2192), .I1(n6703), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1468_3_lut_3_lut (.I0(n2192), .I1(n6702), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4271));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_DFF blue_1128__i1 (.Q(blue[1]), .C(LED_c), .D(n44));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_LUT4 div_43_i1466_3_lut_3_lut (.I0(n2192), .I1(n6700), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1528_3_lut_3_lut (.I0(n2288), .I1(n6718), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1522_3_lut_3_lut (.I0(n2288), .I1(n6712), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1525_3_lut_3_lut (.I0(n2288), .I1(n6715), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1523_3_lut_3_lut (.I0(n2288), .I1(n6713), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1526_3_lut_3_lut (.I0(n2288), .I1(n6716), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1527_3_lut_3_lut (.I0(n2288), .I1(n6717), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3164_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n25097), 
            .O(n6613)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3164_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n25096), 
            .O(n6614)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_12 (.CI(n25096), .I0(n1644), .I1(n90), .CO(n25097));
    SB_LUT4 add_3164_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n25095), 
            .O(n6615)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_11 (.CI(n25095), .I0(n1645), .I1(n91), .CO(n25096));
    SB_LUT4 add_3164_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n25094), 
            .O(n6616)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_10 (.CI(n25094), .I0(n1646), .I1(n92), .CO(n25095));
    SB_LUT4 add_3164_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n25093), 
            .O(n6617)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_9 (.CI(n25093), .I0(n1647), .I1(n93), .CO(n25094));
    SB_LUT4 add_3164_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n25092), 
            .O(n6618)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_8 (.CI(n25092), .I0(n1648), .I1(n94), .CO(n25093));
    SB_LUT4 div_43_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4267));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3164_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n25091), 
            .O(n6619)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_7 (.CI(n25091), .I0(n1649), .I1(n95), .CO(n25092));
    SB_LUT4 add_3164_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n25090), 
            .O(n6620)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_6 (.CI(n25090), .I0(n1650), .I1(n96), .CO(n25091));
    SB_LUT4 add_3164_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n25089), 
            .O(n6621)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_5 (.CI(n25089), .I0(n1651), .I1(n97), .CO(n25090));
    SB_LUT4 add_3164_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n25088), 
            .O(n6622)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_4 (.CI(n25088), .I0(n1652), .I1(n98), .CO(n25089));
    SB_LUT4 add_3164_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n25087), 
            .O(n6623)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_3 (.CI(n25087), .I0(n1653), .I1(n99), .CO(n25088));
    SB_LUT4 add_3164_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6624)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n25087));
    SB_LUT4 add_3163_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n25086), 
            .O(n6600)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3163_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n25085), 
            .O(n6601)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_11 (.CI(n25085), .I0(n1530), .I1(n91), .CO(n25086));
    SB_LUT4 add_3163_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n25084), 
            .O(n6602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_10 (.CI(n25084), .I0(n1531), .I1(n92), .CO(n25085));
    SB_LUT4 add_3163_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n25083), 
            .O(n6603)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_9 (.CI(n25083), .I0(n1532), .I1(n93), .CO(n25084));
    SB_LUT4 add_3163_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n25082), 
            .O(n6604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_8 (.CI(n25082), .I0(n1533), .I1(n94), .CO(n25083));
    SB_LUT4 add_3163_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n25081), 
            .O(n6605)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_7 (.CI(n25081), .I0(n1534), .I1(n95), .CO(n25082));
    SB_LUT4 add_3163_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n25080), 
            .O(n6606)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_6 (.CI(n25080), .I0(n1535), .I1(n96), .CO(n25081));
    SB_LUT4 add_3163_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n25079), 
            .O(n6607)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_5 (.CI(n25079), .I0(n1536), .I1(n97), .CO(n25080));
    SB_LUT4 add_3163_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n25078), 
            .O(n6608)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_4 (.CI(n25078), .I0(n1537), .I1(n98), .CO(n25079));
    SB_LUT4 add_3163_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n25077), 
            .O(n6609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_3 (.CI(n25077), .I0(n1538), .I1(n99), .CO(n25078));
    SB_LUT4 add_3163_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n25077));
    SB_LUT4 add_3162_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n25076), 
            .O(n6588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3162_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n25075), 
            .O(n6589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_10 (.CI(n25075), .I0(n1413), .I1(n92), .CO(n25076));
    SB_LUT4 add_3162_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n25074), 
            .O(n6590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_9 (.CI(n25074), .I0(n1414), .I1(n93), .CO(n25075));
    SB_LUT4 add_3162_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n25073), 
            .O(n6591)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_8 (.CI(n25073), .I0(n1415), .I1(n94), .CO(n25074));
    SB_LUT4 add_3162_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n25072), 
            .O(n6592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_7 (.CI(n25072), .I0(n1416), .I1(n95), .CO(n25073));
    SB_LUT4 add_3162_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n25071), 
            .O(n6593)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_6 (.CI(n25071), .I0(n1417), .I1(n96), .CO(n25072));
    SB_LUT4 add_3162_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n25070), 
            .O(n6594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_5 (.CI(n25070), .I0(n1418), .I1(n97), .CO(n25071));
    SB_LUT4 add_3162_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n25069), 
            .O(n6595)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_4 (.CI(n25069), .I0(n1419), .I1(n98), .CO(n25070));
    SB_LUT4 add_3162_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n25068), 
            .O(n6596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_3 (.CI(n25068), .I0(n1420), .I1(n99), .CO(n25069));
    SB_LUT4 add_3162_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6597)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n25068));
    SB_LUT4 add_3161_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n25044), 
            .O(n6577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3161_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n25043), 
            .O(n6578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_9 (.CI(n25043), .I0(n1293), .I1(n93), .CO(n25044));
    SB_LUT4 add_3161_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n25042), 
            .O(n6579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_8 (.CI(n25042), .I0(n1294), .I1(n94), .CO(n25043));
    SB_LUT4 add_3161_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n25041), 
            .O(n6580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_7 (.CI(n25041), .I0(n1295), .I1(n95), .CO(n25042));
    SB_LUT4 add_3161_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n25040), 
            .O(n6581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_6 (.CI(n25040), .I0(n1296), .I1(n96), .CO(n25041));
    SB_LUT4 add_3161_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n25039), 
            .O(n6582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_5 (.CI(n25039), .I0(n1297), .I1(n97), .CO(n25040));
    SB_LUT4 add_3161_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n25038), 
            .O(n6583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_4 (.CI(n25038), .I0(n1298), .I1(n98), .CO(n25039));
    SB_LUT4 add_3161_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n25037), 
            .O(n6584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_3 (.CI(n25037), .I0(n1299), .I1(n99), .CO(n25038));
    SB_LUT4 add_3161_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n25037));
    SB_LUT4 add_3160_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n25036), 
            .O(n6567)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3160_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n25035), 
            .O(n6568)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_8 (.CI(n25035), .I0(n1170), .I1(n94), .CO(n25036));
    SB_LUT4 add_3160_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n25034), 
            .O(n6569)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_7 (.CI(n25034), .I0(n1171), .I1(n95), .CO(n25035));
    SB_LUT4 add_3160_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n25033), 
            .O(n6570)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_6 (.CI(n25033), .I0(n1172), .I1(n96), .CO(n25034));
    SB_LUT4 add_3160_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n25032), 
            .O(n6571)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_5 (.CI(n25032), .I0(n1173), .I1(n97), .CO(n25033));
    SB_LUT4 add_3160_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n25031), 
            .O(n6572)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_4 (.CI(n25031), .I0(n1174), .I1(n98), .CO(n25032));
    SB_LUT4 add_3160_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n25030), 
            .O(n6573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_3 (.CI(n25030), .I0(n1175), .I1(n99), .CO(n25031));
    SB_LUT4 add_3160_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6574)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n25030));
    SB_LUT4 add_3159_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n25005), 
            .O(n6558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3159_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n25004), 
            .O(n6559)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_7 (.CI(n25004), .I0(n1044), .I1(n95), .CO(n25005));
    SB_LUT4 add_3159_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n25003), 
            .O(n6560)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_6 (.CI(n25003), .I0(n1045), .I1(n96), .CO(n25004));
    SB_LUT4 add_3159_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n25002), 
            .O(n6561)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_5 (.CI(n25002), .I0(n1046), .I1(n97), .CO(n25003));
    SB_LUT4 add_3159_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n25001), 
            .O(n6562)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_4 (.CI(n25001), .I0(n1047), .I1(n98), .CO(n25002));
    SB_LUT4 add_3159_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n25000), 
            .O(n6563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_3 (.CI(n25000), .I0(n1048), .I1(n99), .CO(n25001));
    SB_LUT4 add_3159_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6564)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n25000));
    SB_LUT4 add_3158_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n24999), 
            .O(n6550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3158_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n24998), 
            .O(n6551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_6 (.CI(n24998), .I0(n915), .I1(n96), .CO(n24999));
    SB_LUT4 add_3158_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n24997), 
            .O(n6552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_5 (.CI(n24997), .I0(n916), .I1(n97), .CO(n24998));
    SB_LUT4 div_43_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4268));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3158_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n24996), 
            .O(n6553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4269));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1537_3_lut_3_lut (.I0(n2288), .I1(n6727), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3158_4 (.CI(n24996), .I0(n917), .I1(n98), .CO(n24997));
    SB_LUT4 div_43_i1536_3_lut_3_lut (.I0(n2288), .I1(n6726), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1524_3_lut_3_lut (.I0(n2288), .I1(n6714), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3158_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n24995), 
            .O(n6554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_3 (.CI(n24995), .I0(n918), .I1(n99), .CO(n24996));
    SB_LUT4 add_3158_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n6555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n24995));
    SB_LUT4 div_43_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4258));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4260));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1532_3_lut_3_lut (.I0(n2288), .I1(n6722), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4262));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1531_3_lut_3_lut (.I0(n2288), .I1(n6721), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1530_3_lut_3_lut (.I0(n2288), .I1(n6720), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4264));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4265));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4272));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1539_3_lut_3_lut (.I0(n2288), .I1(n6729), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1529_3_lut_3_lut (.I0(n2288), .I1(n6719), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1534_3_lut_3_lut (.I0(n2288), .I1(n6724), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i28813_4_lut (.I0(n33_adj_4272), .I1(n21_adj_4265), .I2(n19_adj_4264), 
            .I3(n17_adj_4262), .O(n34450));
    defparam i28813_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29478_4_lut (.I0(n15_adj_4260), .I1(n13_adj_4258), .I2(n2552), 
            .I3(n98), .O(n35116));
    defparam i29478_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i29846_4_lut (.I0(n21_adj_4265), .I1(n19_adj_4264), .I2(n17_adj_4262), 
            .I3(n35116), .O(n35485));
    defparam i29846_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29844_4_lut (.I0(n27_adj_4269), .I1(n25_adj_4268), .I2(n23_adj_4267), 
            .I3(n35485), .O(n35483));
    defparam i29844_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_43_i1535_3_lut_3_lut (.I0(n2288), .I1(n6725), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1533_3_lut_3_lut (.I0(n2288), .I1(n6723), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i28815_4_lut (.I0(n33_adj_4272), .I1(n31_adj_4271), .I2(n29_adj_4270), 
            .I3(n35483), .O(n34452));
    defparam i28815_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_i1538_3_lut_3_lut (.I0(n2288), .I1(n6728), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1595_3_lut_3_lut (.I0(n2381), .I1(n6744), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4256));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30192_3_lut (.I0(n10_adj_4256), .I1(n87), .I2(n33_adj_4272), 
            .I3(GND_net), .O(n35831));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30192_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30193_3_lut (.I0(n35831), .I1(n86), .I2(n35_adj_4273), .I3(GND_net), 
            .O(n35832));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30193_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1583_3_lut_3_lut (.I0(n2381), .I1(n6732), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1584_3_lut_3_lut (.I0(n2381), .I1(n6733), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1587_3_lut_3_lut (.I0(n2381), .I1(n6736), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i36_3_lut (.I0(n18_adj_4263), .I1(n83), 
            .I2(n41_adj_4277), .I3(GND_net), .O(n36_adj_4274));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1588_3_lut_3_lut (.I0(n2381), .I1(n6737), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1585_3_lut_3_lut (.I0(n2381), .I1(n6734), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i28808_4_lut (.I0(n39_adj_4276), .I1(n37_adj_4275), .I2(n35_adj_4273), 
            .I3(n34450), .O(n34445));
    defparam i28808_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_i1586_3_lut_3_lut (.I0(n2381), .I1(n6735), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30430_4_lut (.I0(n36_adj_4274), .I1(n16_adj_4261), .I2(n41_adj_4277), 
            .I3(n34441), .O(n36069));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30430_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30121_3_lut (.I0(n35832), .I1(n85), .I2(n37_adj_4275), .I3(GND_net), 
            .O(n35760));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30121_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1601_3_lut_3_lut (.I0(n2381), .I1(n6750), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1596_3_lut_3_lut (.I0(n2381), .I1(n6745), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1665_i22_3_lut (.I0(n14_adj_4259), .I1(n91), 
            .I2(n25_adj_4268), .I3(GND_net), .O(n22_adj_4266));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1592_3_lut_3_lut (.I0(n2381), .I1(n6741), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1600_3_lut_3_lut (.I0(n2381), .I1(n6749), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1599_3_lut_3_lut (.I0(n2381), .I1(n6748), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30428_4_lut (.I0(n22_adj_4266), .I1(n12_adj_4257), .I2(n25_adj_4268), 
            .I3(n34458), .O(n36067));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30428_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30429_3_lut (.I0(n36067), .I1(n90), .I2(n27_adj_4269), .I3(GND_net), 
            .O(n36068));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30429_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1598_3_lut_3_lut (.I0(n2381), .I1(n6747), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30350_3_lut (.I0(n36068), .I1(n89), .I2(n29_adj_4270), .I3(GND_net), 
            .O(n35989));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30350_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1591_3_lut_3_lut (.I0(n2381), .I1(n6740), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30021_4_lut (.I0(n39_adj_4276), .I1(n37_adj_4275), .I2(n35_adj_4273), 
            .I3(n34452), .O(n35660));
    defparam i30021_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_43_i1590_3_lut_3_lut (.I0(n2381), .I1(n6739), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1597_3_lut_3_lut (.I0(n2381), .I1(n6746), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30504_4_lut (.I0(n35760), .I1(n36069), .I2(n41_adj_4277), 
            .I3(n34445), .O(n36143));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30504_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_43_i1589_3_lut_3_lut (.I0(n2381), .I1(n6738), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1594_3_lut_3_lut (.I0(n2381), .I1(n6743), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1593_3_lut_3_lut (.I0(n2381), .I1(n6742), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30320_3_lut (.I0(n35989), .I1(n88), .I2(n31_adj_4271), .I3(GND_net), 
            .O(n35959));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30320_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1655_3_lut_3_lut (.I0(n2471), .I1(n6766), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1642_3_lut_3_lut (.I0(n2471), .I1(n6753), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1644_3_lut_3_lut (.I0(n2471), .I1(n6755), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30518_4_lut (.I0(n35959), .I1(n36143), .I2(n41_adj_4277), 
            .I3(n35660), .O(n36157));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30518_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_25_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30519_3_lut (.I0(n36157), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n36158));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30519_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_43_i1643_3_lut_3_lut (.I0(n2471), .I1(n6754), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30517_3_lut (.I0(n36158), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n36156));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30517_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_43_i1647_3_lut_3_lut (.I0(n2471), .I1(n6758), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1589 (.I0(n36156), .I1(n15487), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1589.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_i1645_3_lut_3_lut (.I0(n2471), .I1(n6756), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4253));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1648_3_lut_3_lut (.I0(n2471), .I1(n6759), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4251));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4255));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4254));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1661_3_lut_3_lut (.I0(n2471), .I1(n6772), .I2(n387), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_3948), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1646_3_lut_3_lut (.I0(n2471), .I1(n6757), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4248));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4249));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1650_3_lut_3_lut (.I0(n2471), .I1(n6761), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1651_3_lut_3_lut (.I0(n2471), .I1(n6762), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1656_3_lut_3_lut (.I0(n2471), .I1(n6767), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4236));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1659_3_lut_3_lut (.I0(n2471), .I1(n6770), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    GND i1 (.Y(GND_net));
    SB_LUT4 div_43_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4238));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1658_3_lut_3_lut (.I0(n2471), .I1(n6769), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i639_3_lut_3_lut (.I0(n938), .I1(n6555), .I2(n373), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1654_3_lut_3_lut (.I0(n2471), .I1(n6765), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4245));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i635_3_lut_3_lut (.I0(n938), .I1(n6551), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4246));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4247));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1653_3_lut_3_lut (.I0(n2471), .I1(n6764), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1652_3_lut_3_lut (.I0(n2471), .I1(n6763), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1649_3_lut_3_lut (.I0(n2471), .I1(n6760), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1657_3_lut_3_lut (.I0(n2471), .I1(n6768), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4250));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1660_3_lut_3_lut (.I0(n2471), .I1(n6771), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4240));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4242));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4243));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28844_4_lut (.I0(n35_adj_4250), .I1(n23_adj_4243), .I2(n21_adj_4242), 
            .I3(n19_adj_4240), .O(n34481));
    defparam i28844_4_lut.LUT_INIT = 16'haaab;
    SB_DFF blue_1128__i2 (.Q(blue[2]), .C(LED_c), .D(n43));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF blue_1128__i3 (.Q(blue[3]), .C(LED_c), .D(n42));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF blue_1128__i4 (.Q(blue[4]), .C(LED_c), .D(n41));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF blue_1128__i5 (.Q(blue[5]), .C(LED_c), .D(n40));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF blue_1128__i6 (.Q(blue[6]), .C(LED_c), .D(n39));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF blue_1128__i7 (.Q(blue[7]), .C(LED_c), .D(n38));   // verilog/TinyFPGA_B.v(51[13:19])
    SB_DFF color_16__55 (.Q(color[16]), .C(LED_c), .D(n17006));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_LUT4 i29504_4_lut (.I0(n17_adj_4238), .I1(n15_adj_4236), .I2(n2464), 
            .I3(n98), .O(n35142));
    defparam i29504_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i29858_4_lut (.I0(n23_adj_4243), .I1(n21_adj_4242), .I2(n19_adj_4240), 
            .I3(n35142), .O(n35497));
    defparam i29858_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF color_17__54 (.Q(color[17]), .C(LED_c), .D(n16984));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_LUT4 i29856_4_lut (.I0(n29_adj_4247), .I1(n27_adj_4246), .I2(n25_adj_4245), 
            .I3(n35497), .O(n35495));
    defparam i29856_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF color_23__48 (.Q(color[23]), .C(LED_c), .D(n16973));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_DFF color_18__53 (.Q(color[18]), .C(LED_c), .D(n16972));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_DFF color_19__52 (.Q(color[19]), .C(LED_c), .D(n16971));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_DFF color_20__51 (.Q(color[20]), .C(LED_c), .D(n16970));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_DFF color_21__50 (.Q(color[21]), .C(LED_c), .D(n16969));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_DFF color_22__49 (.Q(color[22]), .C(LED_c), .D(n16968));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    SB_LUT4 div_43_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4044), .I3(n25589), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_43_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4045), .I3(n25588), .O(n3_adj_3966)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_24 (.CI(n25588), .I0(GND_net), .I1(n3_adj_4045), 
            .CO(n25589));
    SB_LUT4 div_43_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4046), .I3(n25587), .O(n4_adj_3965)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_23 (.CI(n25587), .I0(GND_net), .I1(n4_adj_4046), 
            .CO(n25588));
    SB_LUT4 div_43_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4047), .I3(n25586), .O(n5_adj_3964)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_22 (.CI(n25586), .I0(GND_net), .I1(n5_adj_4047), 
            .CO(n25587));
    SB_LUT4 div_43_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4048), .I3(n25585), .O(n6_adj_3963)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_21 (.CI(n25585), .I0(GND_net), .I1(n6_adj_4048), 
            .CO(n25586));
    SB_LUT4 div_43_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4049), .I3(n25584), .O(n7_adj_3962)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_20 (.CI(n25584), .I0(GND_net), .I1(n7_adj_4049), 
            .CO(n25585));
    SB_LUT4 div_43_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4050), .I3(n25583), .O(n8_adj_3961)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_19 (.CI(n25583), .I0(GND_net), .I1(n8_adj_4050), 
            .CO(n25584));
    SB_LUT4 div_43_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4051), .I3(n25582), .O(n9_adj_3960)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_18 (.CI(n25582), .I0(GND_net), .I1(n9_adj_4051), 
            .CO(n25583));
    SB_LUT4 div_43_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4052), .I3(n25581), .O(n10_adj_3959)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_17 (.CI(n25581), .I0(GND_net), .I1(n10_adj_4052), 
            .CO(n25582));
    SB_LUT4 div_43_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4053), .I3(n25580), .O(n11_adj_3958)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_16 (.CI(n25580), .I0(GND_net), .I1(n11_adj_4053), 
            .CO(n25581));
    SB_LUT4 div_43_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4054), .I3(n25579), .O(n12_adj_3957)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_15 (.CI(n25579), .I0(GND_net), .I1(n12_adj_4054), 
            .CO(n25580));
    SB_LUT4 div_43_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4055), .I3(n25578), .O(n13_adj_3956)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_14 (.CI(n25578), .I0(GND_net), .I1(n13_adj_4055), 
            .CO(n25579));
    SB_LUT4 div_43_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4056), .I3(n25577), .O(n14_adj_3955)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_13 (.CI(n25577), .I0(GND_net), .I1(n14_adj_4056), 
            .CO(n25578));
    SB_LUT4 div_43_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4057), .I3(n25576), .O(n15_adj_3954)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_12 (.CI(n25576), .I0(GND_net), .I1(n15_adj_4057), 
            .CO(n25577));
    SB_LUT4 div_43_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4058), .I3(n25575), .O(n16_adj_3953)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_11 (.CI(n25575), .I0(GND_net), .I1(n16_adj_4058), 
            .CO(n25576));
    SB_LUT4 i28846_4_lut (.I0(n35_adj_4250), .I1(n33_adj_4249), .I2(n31_adj_4248), 
            .I3(n35495), .O(n34483));
    defparam i28846_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4059), .I3(n25574), .O(n17_adj_3952)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_43_LessThan_1606_i12_4_lut (.I0(n387), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4234));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY div_43_unary_minus_2_add_3_10 (.CI(n25574), .I0(GND_net), .I1(n17_adj_4059), 
            .CO(n25575));
    SB_LUT4 div_43_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4060), .I3(n25573), .O(n18_adj_3951)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_9 (.CI(n25573), .I0(GND_net), .I1(n18_adj_4060), 
            .CO(n25574));
    SB_LUT4 div_43_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4061), .I3(n25572), .O(n19_adj_3950)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_8 (.CI(n25572), .I0(GND_net), .I1(n19_adj_4061), 
            .CO(n25573));
    SB_LUT4 div_43_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4062), .I3(n25571), .O(n20_adj_3949)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_7 (.CI(n25571), .I0(GND_net), .I1(n20_adj_4062), 
            .CO(n25572));
    SB_LUT4 div_43_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4063), .I3(n25570), .O(n21_adj_3948)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_6 (.CI(n25570), .I0(GND_net), .I1(n21_adj_4063), 
            .CO(n25571));
    SB_LUT4 div_43_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4064), .I3(n25569), .O(n22_adj_3947)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_5 (.CI(n25569), .I0(GND_net), .I1(n22_adj_4064), 
            .CO(n25570));
    SB_LUT4 div_43_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4065), .I3(n25568), .O(n23_adj_3946)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_4 (.CI(n25568), .I0(GND_net), .I1(n23_adj_4065), 
            .CO(n25569));
    SB_LUT4 div_43_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4066), .I3(n25567), .O(n24_adj_3945)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_3 (.CI(n25567), .I0(GND_net), .I1(n24_adj_4066), 
            .CO(n25568));
    SB_LUT4 div_43_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4067), .I3(VCC_net), .O(n25_adj_3944)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4067), 
            .CO(n25567));
    SB_LUT4 div_43_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4020), .I3(n25566), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_43_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4021), .I3(n25565), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_24 (.CI(n25565), .I0(GND_net), .I1(n3_adj_4021), 
            .CO(n25566));
    SB_LUT4 div_43_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4022), .I3(n25564), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_23 (.CI(n25564), .I0(GND_net), .I1(n4_adj_4022), 
            .CO(n25565));
    SB_LUT4 div_43_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4023), .I3(n25563), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_22 (.CI(n25563), .I0(GND_net), .I1(n5_adj_4023), 
            .CO(n25564));
    SB_LUT4 div_43_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4024), .I3(n25562), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30198_3_lut (.I0(n12_adj_4234), .I1(n87), .I2(n35_adj_4250), 
            .I3(GND_net), .O(n35837));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30198_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_43_unary_minus_4_add_3_21 (.CI(n25562), .I0(GND_net), .I1(n6_adj_4024), 
            .CO(n25563));
    SB_LUT4 div_43_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4025), .I3(n25561), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_20 (.CI(n25561), .I0(GND_net), .I1(n7_adj_4025), 
            .CO(n25562));
    SB_LUT4 div_43_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4026), .I3(n25560), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_19 (.CI(n25560), .I0(GND_net), .I1(n8_adj_4026), 
            .CO(n25561));
    SB_LUT4 div_43_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4027), .I3(n25559), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_18 (.CI(n25559), .I0(GND_net), .I1(n9_adj_4027), 
            .CO(n25560));
    SB_LUT4 div_43_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4028), .I3(n25558), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_17 (.CI(n25558), .I0(GND_net), .I1(n10_adj_4028), 
            .CO(n25559));
    SB_LUT4 div_43_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4029), .I3(n25557), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_16 (.CI(n25557), .I0(GND_net), .I1(n11_adj_4029), 
            .CO(n25558));
    SB_LUT4 div_43_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4030), .I3(n25556), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_15 (.CI(n25556), .I0(GND_net), .I1(n12_adj_4030), 
            .CO(n25557));
    SB_LUT4 div_43_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4031), .I3(n25555), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_14 (.CI(n25555), .I0(GND_net), .I1(n13_adj_4031), 
            .CO(n25556));
    SB_LUT4 div_43_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4032), .I3(n25554), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_13 (.CI(n25554), .I0(GND_net), .I1(n14_adj_4032), 
            .CO(n25555));
    SB_LUT4 div_43_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4033), .I3(n25553), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_12 (.CI(n25553), .I0(GND_net), .I1(n15_adj_4033), 
            .CO(n25554));
    SB_LUT4 div_43_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4034), .I3(n25552), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_11 (.CI(n25552), .I0(GND_net), .I1(n16_adj_4034), 
            .CO(n25553));
    SB_LUT4 div_43_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4035), .I3(n25551), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_10 (.CI(n25551), .I0(GND_net), .I1(n17_adj_4035), 
            .CO(n25552));
    SB_LUT4 div_43_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4036), .I3(n25550), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_9 (.CI(n25550), .I0(GND_net), .I1(n18_adj_4036), 
            .CO(n25551));
    SB_LUT4 div_43_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4037), .I3(n25549), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_8 (.CI(n25549), .I0(GND_net), .I1(n19_adj_4037), 
            .CO(n25550));
    SB_LUT4 div_43_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4038), .I3(n25548), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_7 (.CI(n25548), .I0(GND_net), .I1(n20_adj_4038), 
            .CO(n25549));
    SB_LUT4 div_43_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4039), .I3(n25547), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_6 (.CI(n25547), .I0(GND_net), .I1(n21_adj_4039), 
            .CO(n25548));
    SB_LUT4 div_43_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4040), .I3(n25546), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_5 (.CI(n25546), .I0(GND_net), .I1(n22_adj_4040), 
            .CO(n25547));
    SB_LUT4 div_43_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4041), .I3(n25545), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_4 (.CI(n25545), .I0(GND_net), .I1(n23_adj_4041), 
            .CO(n25546));
    SB_LUT4 div_43_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4042), .I3(n25544), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_3 (.CI(n25544), .I0(GND_net), .I1(n24_adj_4042), 
            .CO(n25545));
    SB_LUT4 div_43_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4043), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_43_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_43_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4043), 
            .CO(n25544));
    SB_LUT4 div_43_LessThan_1606_i38_3_lut (.I0(n20_adj_4241), .I1(n83), 
            .I2(n43_adj_4255), .I3(GND_net), .O(n38_adj_4252));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30199_3_lut (.I0(n35837), .I1(n86), .I2(n37_adj_4251), .I3(GND_net), 
            .O(n35838));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30199_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28840_4_lut (.I0(n41_adj_4254), .I1(n39_adj_4253), .I2(n37_adj_4251), 
            .I3(n34481), .O(n34477));
    defparam i28840_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30196_4_lut (.I0(n38_adj_4252), .I1(n18_adj_4239), .I2(n43_adj_4255), 
            .I3(n34475), .O(n35835));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30196_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30115_3_lut (.I0(n35838), .I1(n85), .I2(n39_adj_4253), .I3(GND_net), 
            .O(n35754));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30115_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1606_i24_3_lut (.I0(n16_adj_4237), .I1(n91), 
            .I2(n27_adj_4246), .I3(GND_net), .O(n24_adj_4244));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_548_24_lut (.I0(duty[22]), .I1(n36858), .I2(n3), .I3(n24749), 
            .O(pwm_setpoint_22__N_17[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i30426_4_lut (.I0(n24_adj_4244), .I1(n14_adj_4235), .I2(n27_adj_4246), 
            .I3(n34489), .O(n36065));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30426_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30427_3_lut (.I0(n36065), .I1(n90), .I2(n29_adj_4247), .I3(GND_net), 
            .O(n36066));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30427_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30352_3_lut (.I0(n36066), .I1(n89), .I2(n31_adj_4248), .I3(GND_net), 
            .O(n35991));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30352_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1712_3_lut_3_lut (.I0(n2558), .I1(n6788), .I2(n2547), 
            .I3(GND_net), .O(n2631_adj_4007));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_548_23_lut (.I0(duty[21]), .I1(n36858), .I2(n4), .I3(n24748), 
            .O(pwm_setpoint_22__N_17[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i30029_4_lut (.I0(n41_adj_4254), .I1(n39_adj_4253), .I2(n37_adj_4251), 
            .I3(n34483), .O(n35668));
    defparam i30029_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30450_4_lut (.I0(n35754), .I1(n35835), .I2(n43_adj_4255), 
            .I3(n34477), .O(n36089));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30450_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_43_i1700_3_lut_3_lut (.I0(n2558), .I1(n6776), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30318_3_lut (.I0(n35991), .I1(n88), .I2(n33_adj_4249), .I3(GND_net), 
            .O(n35957));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30318_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30512_4_lut (.I0(n35957), .I1(n36089), .I2(n43_adj_4255), 
            .I3(n35668), .O(n36151));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30512_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30513_3_lut (.I0(n36151), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n36152));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30513_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1590 (.I0(n36152), .I1(n15484), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1590.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4231));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_17[0]));   // verilog/TinyFPGA_B.v(118[10] 131[6])
    SB_LUT4 div_43_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4233));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4229));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1699_3_lut_3_lut (.I0(n2558), .I1(n6775), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_3949), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_548_23 (.CI(n24748), .I0(n36858), .I1(n4), .CO(n24749));
    SB_LUT4 add_548_22_lut (.I0(duty[20]), .I1(n36858), .I2(n5), .I3(n24747), 
            .O(pwm_setpoint_22__N_17[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_43_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4223));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1702_3_lut_3_lut (.I0(n2558), .I1(n6778), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_548_22 (.CI(n24747), .I0(n36858), .I1(n5), .CO(n24748));
    SB_LUT4 div_43_i1701_3_lut_3_lut (.I0(n2558), .I1(n6777), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4224));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4225));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4232));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1705_3_lut_3_lut (.I0(n2558), .I1(n6781), .I2(n2540), 
            .I3(GND_net), .O(n2624_adj_4000));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4214));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4216));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1703_3_lut_3_lut (.I0(n2558), .I1(n6779), .I2(n2538), 
            .I3(GND_net), .O(n2622_adj_3998));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1706_3_lut_3_lut (.I0(n2558), .I1(n6782), .I2(n2541), 
            .I3(GND_net), .O(n2625_adj_4001));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4218));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4220));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4221));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1719_3_lut_3_lut (.I0(n2558), .I1(n6795), .I2(n388), 
            .I3(GND_net), .O(n2638_adj_4014));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4226));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4227));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4228));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28874_4_lut (.I0(n37_adj_4228), .I1(n25_adj_4221), .I2(n23_adj_4220), 
            .I3(n21_adj_4218), .O(n34511));
    defparam i28874_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29528_4_lut (.I0(n19_adj_4216), .I1(n17_adj_4214), .I2(n2373), 
            .I3(n98), .O(n35166));
    defparam i29528_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i29870_4_lut (.I0(n25_adj_4221), .I1(n23_adj_4220), .I2(n21_adj_4218), 
            .I3(n35166), .O(n35509));
    defparam i29870_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29868_4_lut (.I0(n31_adj_4225), .I1(n29_adj_4224), .I2(n27_adj_4223), 
            .I3(n35509), .O(n35507));
    defparam i29868_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28877_4_lut (.I0(n37_adj_4228), .I1(n35_adj_4227), .I2(n33_adj_4226), 
            .I3(n35507), .O(n34514));
    defparam i28877_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4212));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30202_3_lut (.I0(n14_adj_4212), .I1(n87), .I2(n37_adj_4228), 
            .I3(GND_net), .O(n35841));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30202_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30203_3_lut (.I0(n35841), .I1(n86), .I2(n39_adj_4229), .I3(GND_net), 
            .O(n35842));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30203_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1545_i40_3_lut (.I0(n22_adj_4219), .I1(n83), 
            .I2(n45_adj_4233), .I3(GND_net), .O(n40_adj_4230));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28869_4_lut (.I0(n43_adj_4232), .I1(n41_adj_4231), .I2(n39_adj_4229), 
            .I3(n34511), .O(n34506));
    defparam i28869_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29941_4_lut (.I0(n40_adj_4230), .I1(n20_adj_4217), .I2(n45_adj_4233), 
            .I3(n34504), .O(n35580));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29941_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30111_3_lut (.I0(n35842), .I1(n85), .I2(n41_adj_4231), .I3(GND_net), 
            .O(n35750));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30111_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1704_3_lut_3_lut (.I0(n2558), .I1(n6780), .I2(n2539), 
            .I3(GND_net), .O(n2623_adj_3999));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1545_i26_3_lut (.I0(n18_adj_4215), .I1(n91), 
            .I2(n29_adj_4224), .I3(GND_net), .O(n26_adj_4222));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30424_4_lut (.I0(n26_adj_4222), .I1(n16_adj_4213), .I2(n29_adj_4224), 
            .I3(n34525), .O(n36063));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30424_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30425_3_lut (.I0(n36063), .I1(n90), .I2(n31_adj_4225), .I3(GND_net), 
            .O(n36064));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30425_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30354_3_lut (.I0(n36064), .I1(n89), .I2(n33_adj_4226), .I3(GND_net), 
            .O(n35993));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30354_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30033_4_lut (.I0(n43_adj_4232), .I1(n41_adj_4231), .I2(n39_adj_4229), 
            .I3(n34514), .O(n35672));
    defparam i30033_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30314_4_lut (.I0(n35750), .I1(n35580), .I2(n45_adj_4233), 
            .I3(n34506), .O(n35953));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30314_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30313_3_lut (.I0(n35993), .I1(n88), .I2(n35_adj_4227), .I3(GND_net), 
            .O(n35952));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30313_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30316_4_lut (.I0(n35952), .I1(n35953), .I2(n45_adj_4233), 
            .I3(n35672), .O(n35955));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30316_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(n35955), .I1(n15481), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_i1709_3_lut_3_lut (.I0(n2558), .I1(n6785), .I2(n2544), 
            .I3(GND_net), .O(n2628_adj_4004));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4208));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4211));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4210));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4209));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_3950), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4205));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4206));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1708_3_lut_3_lut (.I0(n2558), .I1(n6784), .I2(n2543), 
            .I3(GND_net), .O(n2627_adj_4003));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4207));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4202));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4204));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1717_3_lut_3_lut (.I0(n2558), .I1(n6793), .I2(n2552), 
            .I3(GND_net), .O(n2636_adj_4012));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1718_3_lut_3_lut (.I0(n2558), .I1(n6794), .I2(n2553), 
            .I3(GND_net), .O(n2637_adj_4013));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4196));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1715_3_lut_3_lut (.I0(n2558), .I1(n6791), .I2(n2550), 
            .I3(GND_net), .O(n2634_adj_4010));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4198));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4200));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4201));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1707_3_lut_3_lut (.I0(n2558), .I1(n6783), .I2(n2542), 
            .I3(GND_net), .O(n2626_adj_4002));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4194));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28929_4_lut (.I0(n23_adj_4200), .I1(n21_adj_4198), .I2(n19_adj_4196), 
            .I3(n17_adj_4194), .O(n34566));
    defparam i28929_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28925_4_lut (.I0(n29_adj_4204), .I1(n27_adj_4202), .I2(n25_adj_4201), 
            .I3(n34566), .O(n34562));
    defparam i28925_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30039_4_lut (.I0(n35_adj_4207), .I1(n33_adj_4206), .I2(n31_adj_4205), 
            .I3(n34562), .O(n35678));
    defparam i30039_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_43_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4193));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_i1716_3_lut_3_lut (.I0(n2558), .I1(n6792), .I2(n2551), 
            .I3(GND_net), .O(n2635_adj_4011));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30208_3_lut (.I0(n16_adj_4193), .I1(n87), .I2(n39_adj_4209), 
            .I3(GND_net), .O(n35847));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30208_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30209_3_lut (.I0(n35847), .I1(n86), .I2(n41_adj_4210), .I3(GND_net), 
            .O(n35848));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30209_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29534_4_lut (.I0(n41_adj_4210), .I1(n39_adj_4209), .I2(n27_adj_4202), 
            .I3(n34564), .O(n35172));
    defparam i29534_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29939_3_lut (.I0(n22_adj_4199), .I1(n93), .I2(n27_adj_4202), 
            .I3(GND_net), .O(n35578));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29939_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30104_3_lut (.I0(n35848), .I1(n85), .I2(n43_adj_4211), .I3(GND_net), 
            .O(n35743));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30104_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1482_i28_3_lut (.I0(n20_adj_4197), .I1(n91), 
            .I2(n31_adj_4205), .I3(GND_net), .O(n28_adj_4203));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30422_4_lut (.I0(n28_adj_4203), .I1(n18_adj_4195), .I2(n31_adj_4205), 
            .I3(n34560), .O(n36061));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30422_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_43_i1711_3_lut_3_lut (.I0(n2558), .I1(n6787), .I2(n2546), 
            .I3(GND_net), .O(n2630_adj_4006));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30423_3_lut (.I0(n36061), .I1(n90), .I2(n33_adj_4206), .I3(GND_net), 
            .O(n36062));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30423_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30356_3_lut (.I0(n36062), .I1(n89), .I2(n35_adj_4207), .I3(GND_net), 
            .O(n35995));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30356_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29536_4_lut (.I0(n41_adj_4210), .I1(n39_adj_4209), .I2(n37_adj_4208), 
            .I3(n35678), .O(n35174));
    defparam i29536_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30206_4_lut (.I0(n35743), .I1(n35578), .I2(n43_adj_4211), 
            .I3(n35172), .O(n35845));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30206_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30311_3_lut (.I0(n35995), .I1(n88), .I2(n37_adj_4208), .I3(GND_net), 
            .O(n35950));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30311_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30440_4_lut (.I0(n35950), .I1(n35845), .I2(n43_adj_4211), 
            .I3(n35174), .O(n36079));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30440_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_43_i1710_3_lut_3_lut (.I0(n2558), .I1(n6786), .I2(n2545), 
            .I3(GND_net), .O(n2629_adj_4005));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30441_3_lut (.I0(n36079), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n36080));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30441_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n36080), .I1(n15478), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'hceef;
    SB_LUT4 i12806_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n12917), .I3(GND_net), .O(n17193));   // verilog/coms.v(126[12] 289[6])
    defparam i12806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1713_3_lut_3_lut (.I0(n2558), .I1(n6789), .I2(n2548), 
            .I3(GND_net), .O(n2632_adj_4008));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4188));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1714_3_lut_3_lut (.I0(n2558), .I1(n6790), .I2(n2549), 
            .I3(GND_net), .O(n2633_adj_4009));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4192));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4191));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4185));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4186));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4187));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4189));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4182));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4184));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_3951), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4175));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4177));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4179));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4181));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4173));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28951_4_lut (.I0(n25_adj_4179), .I1(n23_adj_4177), .I2(n21_adj_4175), 
            .I3(n19_adj_4173), .O(n34588));
    defparam i28951_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28947_4_lut (.I0(n31_adj_4184), .I1(n29_adj_4182), .I2(n27_adj_4181), 
            .I3(n34588), .O(n34584));
    defparam i28947_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30043_4_lut (.I0(n37_adj_4187), .I1(n35_adj_4186), .I2(n33_adj_4185), 
            .I3(n34584), .O(n35682));
    defparam i30043_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_43_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4172));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30212_3_lut (.I0(n18_adj_4172), .I1(n87), .I2(n41_adj_4189), 
            .I3(GND_net), .O(n35851));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30212_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30213_3_lut (.I0(n35851), .I1(n86), .I2(n43_adj_4191), .I3(GND_net), 
            .O(n35852));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30213_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29554_4_lut (.I0(n43_adj_4191), .I1(n41_adj_4189), .I2(n29_adj_4182), 
            .I3(n34586), .O(n35192));
    defparam i29554_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_43_LessThan_1417_i26_3_lut (.I0(n24_adj_4178), .I1(n93), 
            .I2(n29_adj_4182), .I3(GND_net), .O(n26_adj_4180));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30100_3_lut (.I0(n35852), .I1(n85), .I2(n45_adj_4192), .I3(GND_net), 
            .O(n42_adj_4190));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30100_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1417_i30_3_lut (.I0(n22_adj_4176), .I1(n91), 
            .I2(n33_adj_4185), .I3(GND_net), .O(n30_adj_4183));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30420_4_lut (.I0(n30_adj_4183), .I1(n20_adj_4174), .I2(n33_adj_4185), 
            .I3(n34582), .O(n36059));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30420_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30421_3_lut (.I0(n36059), .I1(n90), .I2(n35_adj_4186), .I3(GND_net), 
            .O(n36060));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30421_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30358_3_lut (.I0(n36060), .I1(n89), .I2(n37_adj_4187), .I3(GND_net), 
            .O(n35997));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30358_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29556_4_lut (.I0(n43_adj_4191), .I1(n41_adj_4189), .I2(n39_adj_4188), 
            .I3(n35682), .O(n35194));
    defparam i29556_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29936_4_lut (.I0(n42_adj_4190), .I1(n26_adj_4180), .I2(n45_adj_4192), 
            .I3(n35192), .O(n35575));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29936_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30309_3_lut (.I0(n35997), .I1(n88), .I2(n39_adj_4188), .I3(GND_net), 
            .O(n35948));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30309_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29938_4_lut (.I0(n35948), .I1(n35575), .I2(n45_adj_4192), 
            .I3(n35194), .O(n35577));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29938_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1593 (.I0(n35577), .I1(n15475), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1593.LUT_INIT = 16'hceef;
    SB_LUT4 unary_minus_25_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24_3_lut_adj_1594 (.I0(n34292), .I1(bit_ctr[27]), .I2(n4404), 
            .I3(GND_net), .O(n29077));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1594.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_25_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4171));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 unary_minus_25_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12436_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n15244), 
            .I3(n21347), .O(n16823));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12436_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 div_43_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4170));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12437_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n21347), 
            .I3(n15373), .O(n16824));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12437_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_43_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4169));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12438_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n15244), 
            .I3(n4_adj_3976), .O(n16825));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12438_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12448_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_3976), 
            .I3(n15373), .O(n16835));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12448_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12452_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n15244), 
            .I3(n4_adj_3977), .O(n16839));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12452_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12453_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_3977), 
            .I3(n15373), .O(n16840));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12453_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_43_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4168));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_3952), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4165));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4167));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4043));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4042));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4041));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4040));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4039));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4164));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4038));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4037));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4036));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4158));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4035));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4160));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4162));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4034));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4033));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4156));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4032));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28974_4_lut (.I0(n27_adj_4162), .I1(n25_adj_4160), .I2(n23_adj_4158), 
            .I3(n21_adj_4156), .O(n34611));
    defparam i28974_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28968_4_lut (.I0(n33_adj_4167), .I1(n31_adj_4165), .I2(n29_adj_4164), 
            .I3(n34611), .O(n34605));
    defparam i28968_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i12454_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n15244), 
            .I3(n4_adj_3978), .O(n16841));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12454_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12512_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n16899));   // verilog/coms.v(126[12] 289[6])
    defparam i12512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4031));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4155));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4030));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1350_i28_3_lut (.I0(n26_adj_4161), .I1(n93), 
            .I2(n31_adj_4165), .I3(GND_net), .O(n28_adj_4163));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4029));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12517_3_lut (.I0(encoder0_position[0]), .I1(n2645), .I2(count_enable), 
            .I3(GND_net), .O(n16904));   // quad.v(35[10] 41[6])
    defparam i12517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1595 (.I0(n31_adj_4358), .I1(n30199), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3942));
    defparam i1_2_lut_adj_1595.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(n5_adj_3942), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n32471), .I3(n13117), .O(n47));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'h8caf;
    SB_LUT4 i1_4_lut_adj_1597 (.I0(\FRAME_MATCHER.state [3]), .I1(n47), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n15493), .O(n29611));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1597.LUT_INIT = 16'hccce;
    SB_LUT4 div_43_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4028));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12519_3_lut (.I0(encoder1_position[0]), .I1(n2595), .I2(count_enable_adj_3972), 
            .I3(GND_net), .O(n16906));   // quad.v(35[10] 41[6])
    defparam i12519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1350_i32_3_lut (.I0(n24_adj_4159), .I1(n91), 
            .I2(n35_adj_4168), .I3(GND_net), .O(n32_adj_4166));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12520_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n31114), 
            .I3(GND_net), .O(n16907));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30416_4_lut (.I0(n32_adj_4166), .I1(n22_adj_4157), .I2(n35_adj_4168), 
            .I3(n34602), .O(n36055));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30416_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_43_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4027));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4026));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30417_3_lut (.I0(n36055), .I1(n90), .I2(n37_adj_4169), .I3(GND_net), 
            .O(n36056));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30417_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4025));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4024));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30362_3_lut (.I0(n36056), .I1(n89), .I2(n39_adj_4170), .I3(GND_net), 
            .O(n36001));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30362_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30045_4_lut (.I0(n39_adj_4170), .I1(n37_adj_4169), .I2(n35_adj_4168), 
            .I3(n34605), .O(n35684));
    defparam i30045_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_43_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4023));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30418_4_lut (.I0(n28_adj_4163), .I1(n20_adj_4155), .I2(n31_adj_4165), 
            .I3(n34608), .O(n36057));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30418_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30303_3_lut (.I0(n36001), .I1(n88), .I2(n41_adj_4171), .I3(GND_net), 
            .O(n35942));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30303_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30489_4_lut (.I0(n35942), .I1(n36057), .I2(n41_adj_4171), 
            .I3(n35684), .O(n36128));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30489_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30490_3_lut (.I0(n36128), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n36129));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30490_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30439_3_lut (.I0(n36129), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n36078));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30439_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_43_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4022));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4021));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1598 (.I0(n36078), .I1(n15472), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1598.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4020));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12531_3_lut (.I0(quadB_debounced_adj_3971), .I1(reg_B_adj_4409[0]), 
            .I2(n31841), .I3(GND_net), .O(n16918));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12531_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4067));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4066));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4154));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4152));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4151));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4150));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_3953), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4065));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4064));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4063));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4062));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4061));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12536_4_lut (.I0(n30957), .I1(state[1]), .I2(state_3__N_298[1]), 
            .I3(n16527), .O(n16923));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12536_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i12549_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n925), .I3(GND_net), .O(n16936));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4060));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4059));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4058));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4146));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3185[2]), 
            .I3(r_SM_Main[0]), .O(n16501));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 div_43_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4147));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4057));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4149));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n16501), 
            .I3(rx_data_ready), .O(n29853));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 div_43_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4056));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22_3_lut_adj_1599 (.I0(bit_ctr[28]), .I1(n34293), .I2(n4404), 
            .I3(GND_net), .O(n29079));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1599.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4140));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4055));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4142));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4144));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4054));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4138));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4053));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28996_4_lut (.I0(n29_adj_4144), .I1(n27_adj_4142), .I2(n25_adj_4140), 
            .I3(n23_adj_4138), .O(n34633));
    defparam i28996_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28991_4_lut (.I0(n35_adj_4149), .I1(n33_adj_4147), .I2(n31_adj_4146), 
            .I3(n34633), .O(n34628));
    defparam i28991_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4052));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4137));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_LessThan_1281_i30_3_lut (.I0(n28_adj_4143), .I1(n93), 
            .I2(n33_adj_4147), .I3(GND_net), .O(n30_adj_4145));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4051));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1281_i34_3_lut (.I0(n26_adj_4141), .I1(n91), 
            .I2(n37_adj_4150), .I3(GND_net), .O(n34_adj_4148));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30414_4_lut (.I0(n34_adj_4148), .I1(n24_adj_4139), .I2(n37_adj_4150), 
            .I3(n34626), .O(n36053));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30414_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30415_3_lut (.I0(n36053), .I1(n90), .I2(n39_adj_4151), .I3(GND_net), 
            .O(n36054));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30415_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30364_3_lut (.I0(n36054), .I1(n89), .I2(n41_adj_4152), .I3(GND_net), 
            .O(n36003));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30364_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4050));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30047_4_lut (.I0(n41_adj_4152), .I1(n39_adj_4151), .I2(n37_adj_4150), 
            .I3(n34628), .O(n35686));
    defparam i30047_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30218_4_lut (.I0(n30_adj_4145), .I1(n22_adj_4137), .I2(n33_adj_4147), 
            .I3(n34631), .O(n35857));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30218_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_43_i634_3_lut_3_lut (.I0(n938), .I1(n6550), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30299_3_lut (.I0(n36003), .I1(n88), .I2(n43_adj_4154), .I3(GND_net), 
            .O(n42_adj_4153));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30299_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4049));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30377_4_lut (.I0(n42_adj_4153), .I1(n35857), .I2(n43_adj_4154), 
            .I3(n35686), .O(n36016));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30377_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30378_3_lut (.I0(n36016), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n36017));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30378_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_43_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4048));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1600 (.I0(n36017), .I1(n15469), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1600.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4047));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4046));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_i1769_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6813), .I2(n2633_adj_4009), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4045));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4044));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12581_3_lut (.I0(color[22]), .I1(blue[6]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16968));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4136));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12582_3_lut (.I0(color[21]), .I1(blue[5]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16969));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1754_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6798), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4134));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12583_3_lut (.I0(color[20]), .I1(blue[4]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16970));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12584_3_lut (.I0(color[19]), .I1(blue[3]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16971));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12585_3_lut (.I0(color[18]), .I1(blue[2]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16972));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12586_3_lut (.I0(color[23]), .I1(blue[7]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16973));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4133));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4132));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12587_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n29225), .I3(GND_net), .O(n16974));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12588_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n29225), .I3(GND_net), .O(n16975));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12589_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n29225), .I3(GND_net), .O(n16976));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12590_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n29225), .I3(GND_net), .O(n16977));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1755_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6799), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_3954), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12591_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n29225), .I3(GND_net), .O(n16978));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12592_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n29225), .I3(GND_net), .O(n16979));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4128));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4129));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4131));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4122));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4124));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4126));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4120));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i29034_4_lut (.I0(n31_adj_4126), .I1(n29_adj_4124), .I2(n27_adj_4122), 
            .I3(n25_adj_4120), .O(n34671));
    defparam i29034_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29030_4_lut (.I0(n37_adj_4131), .I1(n35_adj_4129), .I2(n33_adj_4128), 
            .I3(n34671), .O(n34667));
    defparam i29030_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4119));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_43_LessThan_1210_i32_3_lut (.I0(n30_adj_4125), .I1(n93), 
            .I2(n35_adj_4129), .I3(GND_net), .O(n32_adj_4127));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1210_i36_3_lut (.I0(n28_adj_4123), .I1(n91), 
            .I2(n39_adj_4132), .I3(GND_net), .O(n36_adj_4130));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30412_4_lut (.I0(n36_adj_4130), .I1(n26_adj_4121), .I2(n39_adj_4132), 
            .I3(n34643), .O(n36051));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30412_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30413_3_lut (.I0(n36051), .I1(n90), .I2(n41_adj_4133), .I3(GND_net), 
            .O(n36052));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30413_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30366_3_lut (.I0(n36052), .I1(n89), .I2(n43_adj_4134), .I3(GND_net), 
            .O(n36005));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30366_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30053_4_lut (.I0(n43_adj_4134), .I1(n41_adj_4133), .I2(n39_adj_4132), 
            .I3(n34667), .O(n35692));
    defparam i30053_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30081_4_lut (.I0(n32_adj_4127), .I1(n24_adj_4119), .I2(n35_adj_4129), 
            .I3(n34669), .O(n35720));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30081_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12593_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n29225), .I3(GND_net), .O(n16980));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30297_3_lut (.I0(n36005), .I1(n88), .I2(n45_adj_4136), .I3(GND_net), 
            .O(n44_adj_4135));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30297_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30083_4_lut (.I0(n44_adj_4135), .I1(n35720), .I2(n45_adj_4136), 
            .I3(n35692), .O(n35722));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30083_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12594_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n29225), .I3(GND_net), .O(n16981));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12594_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(n35722), .I1(n15466), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'hceef;
    SB_LUT4 i12595_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n29225), .I3(GND_net), .O(n16982));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12595_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12596_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n29225), .I3(GND_net), .O(n16983));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12597_3_lut (.I0(color[17]), .I1(blue[1]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n16984));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12598_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n29225), .I3(GND_net), .O(n16985));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4115));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1756_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6800), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12599_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n29225), .I3(GND_net), .O(n16986));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12599_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4114));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12600_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n29225), .I3(GND_net), .O(n16987));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12600_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12601_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n29225), .I3(GND_net), .O(n16988));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12602_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n29225), .I3(GND_net), .O(n16989));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_3955), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12603_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n29225), .I3(GND_net), .O(n16990));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12603_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1757_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6801), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1758_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6802), .I2(n2622_adj_3998), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4118));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12604_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n29225), .I3(GND_net), .O(n16991));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12604_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12605_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n29225), .I3(GND_net), .O(n16992));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12605_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4117));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12606_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n29225), .I3(GND_net), .O(n16993));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12606_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12607_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n29225), .I3(GND_net), .O(n16994));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4110));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12608_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n29225), .I3(GND_net), .O(n16995));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4112));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12609_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n29225), .I3(GND_net), .O(n16996));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12609_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4113));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12610_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n29225), .I3(GND_net), .O(n16997));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12610_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12611_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n29225), .I3(GND_net), .O(n16998));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12611_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29048_4_lut (.I0(n33_adj_4113), .I1(n31_adj_4112), .I2(n29_adj_4110), 
            .I3(n27), .O(n34685));
    defparam i29048_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i12612_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n29225), .I3(GND_net), .O(n16999));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12612_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12613_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n29225), .I3(GND_net), .O(n17000));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12613_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12614_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n29225), .I3(GND_net), .O(n17001));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12614_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1137_i38_3_lut (.I0(n30_adj_4111), .I1(n91), 
            .I2(n41_adj_4118), .I3(GND_net), .O(n38_adj_4116));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30226_3_lut (.I0(n26), .I1(n95), .I2(n33_adj_4113), .I3(GND_net), 
            .O(n35865));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30226_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12615_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n29225), .I3(GND_net), .O(n17002));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30227_3_lut (.I0(n35865), .I1(n94), .I2(n35_adj_4114), .I3(GND_net), 
            .O(n35866));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30227_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29044_4_lut (.I0(n39_adj_4117), .I1(n37_adj_4115), .I2(n35_adj_4114), 
            .I3(n34685), .O(n34681));
    defparam i29044_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i12616_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n29225), .I3(GND_net), .O(n17003));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30410_4_lut (.I0(n38_adj_4116), .I1(n28_adj_4109), .I2(n41_adj_4118), 
            .I3(n34679), .O(n36049));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30410_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30076_3_lut (.I0(n35866), .I1(n93), .I2(n37_adj_4115), .I3(GND_net), 
            .O(n35715));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30076_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30502_4_lut (.I0(n35715), .I1(n36049), .I2(n41_adj_4118), 
            .I3(n34681), .O(n36141));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30502_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12617_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n29225), .I3(GND_net), .O(n17004));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12617_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30503_3_lut (.I0(n36141), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n36142));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30503_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30484_3_lut (.I0(n36142), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n36123));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30484_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(n36123), .I1(n15463), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'hceef;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_3937));   // verilog/TinyFPGA_B.v(206[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4105));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4104));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_3956), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4108));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4107));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4100));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4102));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4103));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12618_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n29225), .I3(GND_net), .O(n17005));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12618_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29066_4_lut (.I0(n35_adj_4103), .I1(n33_adj_4102), .I2(n31_adj_4100), 
            .I3(n29), .O(n34703));
    defparam i29066_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_i1775_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6819), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12619_3_lut (.I0(color[16]), .I1(blue[0]), .I2(send_to_neopixels), 
            .I3(GND_net), .O(n17006));   // verilog/TinyFPGA_B.v(46[8] 53[4])
    defparam i12619_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .GND_net(GND_net), .rx_data({rx_data}), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .n37085(n37085), .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), 
         .PWMLimit({PWMLimit}), .control_mode({control_mode}), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n17214(n17214), .n17213(n17213), .n17212(n17212), .n17211(n17211), 
         .n17210(n17210), .n17209(n17209), .n17208(n17208), .n17207(n17207), 
         .n17206(n17206), .n17205(n17205), .n17204(n17204), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n63(n63_adj_4017), .n31(n31_adj_4358), .n2421(n2421), .n13117(n13117), 
         .n17203(n17203), .n17202(n17202), .rx_data_ready(rx_data_ready), 
         .n17201(n17201), .n17200(n17200), .n17199(n17199), .n17198(n17198), 
         .n30199(n30199), .n17197(n17197), .n17196(n17196), .n17195(n17195), 
         .n17194(n17194), .n17193(n17193), .n17192(n17192), .n17191(n17191), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .n3915(n3915), 
         .n12917(n12917), .n17190(n17190), .n17189(n17189), .n17188(n17188), 
         .n17187(n17187), .n17186(n17186), .n17185(n17185), .n17184(n17184), 
         .\r_SM_Main_2__N_3259[0] (r_SM_Main_2__N_3259[0]), .n17183(n17183), 
         .n17182(n17182), .n17181(n17181), .n17180(n17180), .n17179(n17179), 
         .n17178(n17178), .n17177(n17177), .n17176(n17176), .n17175(n17175), 
         .n17174(n17174), .n17173(n17173), .n17172(n17172), .n17171(n17171), 
         .n17170(n17170), .n17169(n17169), .n17168(n17168), .n17167(n17167), 
         .n17166(n17166), .n17165(n17165), .n17164(n17164), .n17163(n17163), 
         .n17162(n17162), .n17161(n17161), .n17160(n17160), .n17159(n17159), 
         .n17158(n17158), .n17157(n17157), .n17156(n17156), .n17155(n17155), 
         .n17154(n17154), .n17153(n17153), .n17152(n17152), .n17151(n17151), 
         .n17150(n17150), .n17149(n17149), .n17148(n17148), .n17147(n17147), 
         .\data_in[3] ({\data_in[3] }), .\data_in[0] ({\data_in[0] }), .\data_in[2] ({\data_in[2] }), 
         .\data_in[1] ({\data_in[1] }), .n3761(n3761), .n22044(n22044), 
         .n740(n740), .n17146(n17146), .n17145(n17145), .n17144(n17144), 
         .n17143(n17143), .n17142(n17142), .n17141(n17141), .n17140(n17140), 
         .n17139(n17139), .n17138(n17138), .n17137(n17137), .n17136(n17136), 
         .n17135(n17135), .n17134(n17134), .n17133(n17133), .n15494(n15494), 
         .n15502(n15502), .n17132(n17132), .n15493(n15493), .n18493(n18493), 
         .n5(n5_adj_4018), .n37539(n37539), .n17131(n17131), .n17130(n17130), 
         .n17129(n17129), .n17128(n17128), .n17127(n17127), .n17126(n17126), 
         .n17125(n17125), .n17124(n17124), .n17123(n17123), .n17122(n17122), 
         .n17121(n17121), .n17120(n17120), .n17119(n17119), .n17118(n17118), 
         .n17117(n17117), .n17116(n17116), .n17115(n17115), .n17114(n17114), 
         .n17113(n17113), .n17112(n17112), .n17111(n17111), .n17110(n17110), 
         .n17109(n17109), .n17108(n17108), .n17107(n17107), .n17106(n17106), 
         .n17105(n17105), .n17104(n17104), .n17103(n17103), .n17102(n17102), 
         .n17101(n17101), .n17100(n17100), .n17099(n17099), .n17098(n17098), 
         .n17097(n17097), .n17096(n17096), .n17095(n17095), .n17094(n17094), 
         .n17093(n17093), .n17092(n17092), .n17091(n17091), .n17090(n17090), 
         .n17089(n17089), .n17088(n17088), .n17087(n17087), .n17086(n17086), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n17085(n17085), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n17084(n17084), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .\Kp[7] (Kp[7]), 
         .\Kp[6] (Kp[6]), .\Kp[5] (Kp[5]), .\Kp[4] (Kp[4]), .\Kp[3] (Kp[3]), 
         .\Kp[2] (Kp[2]), .\Kp[1] (Kp[1]), .n17076(n17076), .n17075(n17075), 
         .n17074(n17074), .n17073(n17073), .n17072(n17072), .n17071(n17071), 
         .n17070(n17070), .n17069(n17069), .n17068(n17068), .n17067(n17067), 
         .n15501(n15501), .n17066(n17066), .n17065(n17065), .n17064(n17064), 
         .n17063(n17063), .n17062(n17062), .n17061(n17061), .n17060(n17060), 
         .n17059(n17059), .n17058(n17058), .n17057(n17057), .n17056(n17056), 
         .n17055(n17055), .n17054(n17054), .n17053(n17053), .n17052(n17052), 
         .n17051(n17051), .n17050(n17050), .n17049(n17049), .n17048(n17048), 
         .n17047(n17047), .n17046(n17046), .n17040(n17040), .setpoint({setpoint}), 
         .n17039(n17039), .n17038(n17038), .n17037(n17037), .n17036(n17036), 
         .n17035(n17035), .n17034(n17034), .n17033(n17033), .n17032(n17032), 
         .n17031(n17031), .n17030(n17030), .n17029(n17029), .n17028(n17028), 
         .n17027(n17027), .n17026(n17026), .n17025(n17025), .n17024(n17024), 
         .n17023(n17023), .n17022(n17022), .n17021(n17021), .n17020(n17020), 
         .n17019(n17019), .gearBoxRatio({gearBoxRatio}), .n16770(n16770), 
         .n17018(n17018), .LED_c(LED_c), .n29611(n29611), .\Kp[0] (Kp[0]), 
         .n16899(n16899), .n4335(n4335), .n4312(n4312), .n4334(n4334), 
         .n4333(n4333), .n4332(n4332), .n4331(n4331), .n4330(n4330), 
         .n4329(n4329), .n4328(n4328), .n4327(n4327), .n4326(n4326), 
         .n4325(n4325), .n4324(n4324), .n4323(n4323), .n4322(n4322), 
         .n4321(n4321), .n4320(n4320), .n4319(n4319), .n4318(n4318), 
         .n4317(n4317), .n4316(n4316), .n4315(n4315), .n4314(n4314), 
         .n31259(n31259), .n4313(n4313), .n15495(n15495), .n5_adj_3(n5_adj_4359), 
         .tx_active(tx_active), .n16549(n16549), .VCC_net(VCC_net), .tx_o(tx_o), 
         .tx_enable(tx_enable), .n16816(n16816), .r_Bit_Index({r_Bit_Index}), 
         .n16819(n16819), .n29853(n29853), .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3185[2] (r_SM_Main_2__N_3185[2]), 
         .r_Rx_Data(r_Rx_Data), .PIN_13_N_65(PIN_13_N_65), .n16600(n16600), 
         .n16687(n16687), .n4573(n4573), .n17013(n17013), .n16841(n16841), 
         .n16840(n16840), .n16839(n16839), .n16835(n16835), .n16825(n16825), 
         .n16824(n16824), .n16823(n16823), .n21347(n21347), .n4(n4_adj_3976), 
         .n4_adj_4(n4_adj_3977), .n15244(n15244), .n15373(n15373), .n4_adj_5(n4_adj_3978)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(159[8] 179[4])
    SB_LUT4 div_43_i1761_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6805), .I2(n2625_adj_4001), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12626_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_3978), 
            .I3(n15373), .O(n17013));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12626_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i22_3_lut_adj_1603 (.I0(bit_ctr[29]), .I1(n34294), .I2(n4404), 
            .I3(GND_net), .O(n29081));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1603.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_1062_i40_3_lut (.I0(n32_adj_4101), .I1(n91), 
            .I2(n43_adj_4108), .I3(GND_net), .O(n40_adj_4106));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_i1762_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6806), .I2(n2626_adj_4002), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i12631_3_lut (.I0(setpoint[23]), .I1(n4335), .I2(n31259), 
            .I3(GND_net), .O(n17018));   // verilog/coms.v(126[12] 289[6])
    defparam i12631_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30230_3_lut (.I0(n28), .I1(n95), .I2(n35_adj_4103), .I3(GND_net), 
            .O(n35869));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30230_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12383_3_lut (.I0(setpoint[0]), .I1(n4312), .I2(n31259), .I3(GND_net), 
            .O(n16770));   // verilog/coms.v(126[12] 289[6])
    defparam i12383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30231_3_lut (.I0(n35869), .I1(n94), .I2(n37_adj_4104), .I3(GND_net), 
            .O(n35870));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30231_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29061_4_lut (.I0(n41_adj_4107), .I1(n39_adj_4105), .I2(n37_adj_4104), 
            .I3(n34703), .O(n34698));
    defparam i29061_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_i1764_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6808), .I2(n2628_adj_4004), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30228_4_lut (.I0(n40_adj_4106), .I1(n30_adj_4099), .I2(n43_adj_4108), 
            .I3(n34695), .O(n35867));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30228_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30072_3_lut (.I0(n35870), .I1(n93), .I2(n39_adj_4105), .I3(GND_net), 
            .O(n35711));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30072_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12384_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n29225), .I3(GND_net), .O(n16771));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30458_4_lut (.I0(n35711), .I1(n35867), .I2(n43_adj_4108), 
            .I3(n34698), .O(n36097));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30459_3_lut (.I0(n36097), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n36098));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30459_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_43_i1765_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6809), .I2(n2629_adj_4005), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n36098), .I1(n15460), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'hceef;
    SB_LUT4 i12632_3_lut (.I0(setpoint[22]), .I1(n4334), .I2(n31259), 
            .I3(GND_net), .O(n17019));   // verilog/coms.v(126[12] 289[6])
    defparam i12632_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12633_3_lut (.I0(setpoint[21]), .I1(n4333), .I2(n31259), 
            .I3(GND_net), .O(n17020));   // verilog/coms.v(126[12] 289[6])
    defparam i12633_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4095));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12634_3_lut (.I0(setpoint[20]), .I1(n4332), .I2(n31259), 
            .I3(GND_net), .O(n17021));   // verilog/coms.v(126[12] 289[6])
    defparam i12634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12635_3_lut (.I0(setpoint[19]), .I1(n4331), .I2(n31259), 
            .I3(GND_net), .O(n17022));   // verilog/coms.v(126[12] 289[6])
    defparam i12635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4094));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_3957), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4098));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4097));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4093));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i29081_4_lut (.I0(n37_adj_4093), .I1(n35), .I2(n33), .I3(n31), 
            .O(n34718));
    defparam i29081_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_43_LessThan_985_i42_3_lut (.I0(n34_adj_4092), .I1(n91), 
            .I2(n45_adj_4098), .I3(GND_net), .O(n42_adj_4096));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_43_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30290_3_lut (.I0(n30), .I1(n95), .I2(n37_adj_4093), .I3(GND_net), 
            .O(n35929));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30290_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12636_3_lut (.I0(setpoint[18]), .I1(n4330), .I2(n31259), 
            .I3(GND_net), .O(n17023));   // verilog/coms.v(126[12] 289[6])
    defparam i12636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1766_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6810), .I2(n2630_adj_4006), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30291_3_lut (.I0(n35929), .I1(n94), .I2(n39_adj_4094), .I3(GND_net), 
            .O(n35930));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30291_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29076_4_lut (.I0(n43_adj_4097), .I1(n41_adj_4095), .I2(n39_adj_4094), 
            .I3(n34718), .O(n34713));
    defparam i29076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29930_4_lut (.I0(n42_adj_4096), .I1(n32_adj_4091), .I2(n45_adj_4098), 
            .I3(n34711), .O(n35569));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29930_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30070_3_lut (.I0(n35930), .I1(n93), .I2(n41_adj_4095), .I3(GND_net), 
            .O(n35709));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30070_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30292_4_lut (.I0(n35709), .I1(n35569), .I2(n45_adj_4098), 
            .I3(n34713), .O(n35931));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30292_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1605 (.I0(n35931), .I1(n15457), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1605.LUT_INIT = 16'hceef;
    SB_LUT4 i12637_3_lut (.I0(setpoint[17]), .I1(n4329), .I2(n31259), 
            .I3(GND_net), .O(n17024));   // verilog/coms.v(126[12] 289[6])
    defparam i12637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4090));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4089));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4088));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_3958), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1767_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6811), .I2(n2631_adj_4007), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1773_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6817), .I2(n2637_adj_4013), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12638_3_lut (.I0(setpoint[16]), .I1(n4328), .I2(n31259), 
            .I3(GND_net), .O(n17025));   // verilog/coms.v(126[12] 289[6])
    defparam i12638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12639_3_lut (.I0(setpoint[15]), .I1(n4327), .I2(n31259), 
            .I3(GND_net), .O(n17026));   // verilog/coms.v(126[12] 289[6])
    defparam i12639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1774_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6818), .I2(n2638_adj_4014), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1759_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6803), .I2(n2623_adj_3999), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_43_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30067_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4088), .I3(GND_net), 
            .O(n35706));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30067_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12640_3_lut (.I0(setpoint[14]), .I1(n4326), .I2(n31259), 
            .I3(GND_net), .O(n17027));   // verilog/coms.v(126[12] 289[6])
    defparam i12640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30068_3_lut (.I0(n35706), .I1(n94), .I2(n41_adj_4089), .I3(GND_net), 
            .O(n35707));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30068_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29693_4_lut (.I0(n41_adj_4089), .I1(n39_adj_4088), .I2(n37), 
            .I3(n34742), .O(n35331));
    defparam i29693_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29926_3_lut (.I0(n34_adj_4087), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n35565));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29926_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29687_3_lut (.I0(n35707), .I1(n93), .I2(n43_adj_4090), .I3(GND_net), 
            .O(n35325));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29687_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12641_3_lut (.I0(setpoint[13]), .I1(n4325), .I2(n31259), 
            .I3(GND_net), .O(n17028));   // verilog/coms.v(126[12] 289[6])
    defparam i12641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29979_4_lut (.I0(n35325), .I1(n35565), .I2(n43_adj_4090), 
            .I3(n35331), .O(n35618));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29979_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12642_3_lut (.I0(setpoint[12]), .I1(n4324), .I2(n31259), 
            .I3(GND_net), .O(n17029));   // verilog/coms.v(126[12] 289[6])
    defparam i12642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29980_3_lut (.I0(n35618), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n35619));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29980_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1606 (.I0(n35619), .I1(n15454), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1606.LUT_INIT = 16'hceef;
    SB_LUT4 div_43_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4083));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12643_3_lut (.I0(setpoint[11]), .I1(n4323), .I2(n31259), 
            .I3(GND_net), .O(n17030));   // verilog/coms.v(126[12] 289[6])
    defparam i12643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4086));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12644_3_lut (.I0(setpoint[10]), .I1(n4322), .I2(n31259), 
            .I3(GND_net), .O(n17031));   // verilog/coms.v(126[12] 289[6])
    defparam i12644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1768_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6812), .I2(n2632_adj_4008), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_3959), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12645_3_lut (.I0(setpoint[9]), .I1(n4321), .I2(n31259), .I3(GND_net), 
            .O(n17032));   // verilog/coms.v(126[12] 289[6])
    defparam i12645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4085));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12646_3_lut (.I0(setpoint[8]), .I1(n4320), .I2(n31259), .I3(GND_net), 
            .O(n17033));   // verilog/coms.v(126[12] 289[6])
    defparam i12646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4084));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_43_i1763_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6807), .I2(n2627_adj_4003), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12647_3_lut (.I0(setpoint[7]), .I1(n4319), .I2(n31259), .I3(GND_net), 
            .O(n17034));   // verilog/coms.v(126[12] 289[6])
    defparam i12647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i1771_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6815), .I2(n2635_adj_4011), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i1760_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6804), .I2(n2624_adj_4000), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12648_3_lut (.I0(setpoint[6]), .I1(n4318), .I2(n31259), .I3(GND_net), 
            .O(n17035));   // verilog/coms.v(126[12] 289[6])
    defparam i12648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12649_3_lut (.I0(setpoint[5]), .I1(n4317), .I2(n31259), .I3(GND_net), 
            .O(n17036));   // verilog/coms.v(126[12] 289[6])
    defparam i12649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12650_3_lut (.I0(setpoint[4]), .I1(n4316), .I2(n31259), .I3(GND_net), 
            .O(n17037));   // verilog/coms.v(126[12] 289[6])
    defparam i12650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i29981_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4084), .I3(GND_net), 
            .O(n35620));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29981_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12651_3_lut (.I0(setpoint[3]), .I1(n4315), .I2(n31259), .I3(GND_net), 
            .O(n17038));   // verilog/coms.v(126[12] 289[6])
    defparam i12651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29982_3_lut (.I0(n35620), .I1(n94), .I2(n43_adj_4085), .I3(GND_net), 
            .O(n35621));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29982_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29699_4_lut (.I0(n43_adj_4085), .I1(n41_adj_4084), .I2(n39_adj_4083), 
            .I3(n34761), .O(n35337));
    defparam i29699_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i12652_3_lut (.I0(setpoint[2]), .I1(n4314), .I2(n31259), .I3(GND_net), 
            .O(n17039));   // verilog/coms.v(126[12] 289[6])
    defparam i12652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_43_LessThan_825_i38_3_lut (.I0(n36_adj_4081), .I1(n96), 
            .I2(n39_adj_4083), .I3(GND_net), .O(n38_adj_4082));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29685_3_lut (.I0(n35621), .I1(n93), .I2(n45_adj_4086), .I3(GND_net), 
            .O(n35323));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29685_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12653_3_lut (.I0(setpoint[1]), .I1(n4313), .I2(n31259), .I3(GND_net), 
            .O(n17040));   // verilog/coms.v(126[12] 289[6])
    defparam i12653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30065_4_lut (.I0(n35323), .I1(n38_adj_4082), .I2(n45_adj_4086), 
            .I3(n35337), .O(n35704));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30065_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n35704), .I1(n15451), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'hceef;
    SB_LUT4 i29254_4_lut (.I0(state[0]), .I1(start), .I2(n22016), .I3(\neo_pixel_transmitter.done ), 
            .O(n34298));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29254_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i29300_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34300));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29300_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_43_i1772_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6816), .I2(n2636_adj_4012), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i18_4_lut (.I0(n34300), .I1(n34298), .I2(state[1]), .I3(n22030), 
            .O(n29087));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i12659_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17046));   // verilog/coms.v(126[12] 289[6])
    defparam i12659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12660_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17047));   // verilog/coms.v(126[12] 289[6])
    defparam i12660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_3960), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12661_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17048));   // verilog/coms.v(126[12] 289[6])
    defparam i12661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12662_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17049));   // verilog/coms.v(126[12] 289[6])
    defparam i12662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12663_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17050));   // verilog/coms.v(126[12] 289[6])
    defparam i12663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12664_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17051));   // verilog/coms.v(126[12] 289[6])
    defparam i12664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4080));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12665_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17052));   // verilog/coms.v(126[12] 289[6])
    defparam i12665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12666_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17053));   // verilog/coms.v(126[12] 289[6])
    defparam i12666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12667_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17054));   // verilog/coms.v(126[12] 289[6])
    defparam i12667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12668_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17055));   // verilog/coms.v(126[12] 289[6])
    defparam i12668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12669_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17056));   // verilog/coms.v(126[12] 289[6])
    defparam i12669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12670_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17057));   // verilog/coms.v(126[12] 289[6])
    defparam i12670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12671_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17058));   // verilog/coms.v(126[12] 289[6])
    defparam i12671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i12672_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17059));   // verilog/coms.v(126[12] 289[6])
    defparam i12672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_742_i40_3_lut (.I0(n38_adj_4078), .I1(n96), 
            .I2(n41_adj_4080), .I3(GND_net), .O(n40_adj_4079));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30373_4_lut (.I0(n40_adj_4079), .I1(n36), .I2(n41_adj_4080), 
            .I3(n34768), .O(n36012));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30373_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12673_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17060));   // verilog/coms.v(126[12] 289[6])
    defparam i12673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30374_3_lut (.I0(n36012), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n36013));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30374_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30233_3_lut (.I0(n36013), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n35872));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i30233_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i12674_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17061));   // verilog/coms.v(126[12] 289[6])
    defparam i12674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n35872), .I1(n15448), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'hceef;
    SB_LUT4 i12699_3_lut_4_lut (.I0(\data_out_frame[0] [4]), .I1(n3915), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n16549), .O(n17086));   // verilog/coms.v(126[12] 289[6])
    defparam i12699_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i12698_3_lut_4_lut (.I0(\data_out_frame[0] [3]), .I1(n3915), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n16549), .O(n17085));   // verilog/coms.v(126[12] 289[6])
    defparam i12698_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i12675_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17062));   // verilog/coms.v(126[12] 289[6])
    defparam i12675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12697_3_lut_4_lut (.I0(\data_out_frame[0] [2]), .I1(n3915), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n16549), .O(n17084));   // verilog/coms.v(126[12] 289[6])
    defparam i12697_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i12676_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17063));   // verilog/coms.v(126[12] 289[6])
    defparam i12676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12677_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17064));   // verilog/coms.v(126[12] 289[6])
    defparam i12677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12678_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17065));   // verilog/coms.v(126[12] 289[6])
    defparam i12678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i1770_3_lut_3_lut (.I0(n2642_adj_4015), .I1(n6814), .I2(n2634_adj_4010), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4071));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12679_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17066));   // verilog/coms.v(126[12] 289[6])
    defparam i12679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4091));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29074_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n34711));
    defparam i29074_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4092));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4099));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29058_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n34695));
    defparam i29058_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i29141_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n34778));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29141_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4101));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4109));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29042_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n34679));
    defparam i29042_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4111));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29137_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n34774));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29137_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12680_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17067));   // verilog/coms.v(126[12] 289[6])
    defparam i12680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12681_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17068));   // verilog/coms.v(126[12] 289[6])
    defparam i12681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4121));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29006_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n34643));
    defparam i29006_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4123));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29032_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n34669));
    defparam i29032_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4125));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4139));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28989_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n34626));
    defparam i28989_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4141));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28994_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n34631));
    defparam i28994_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4143));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n17466(n17466), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n17465(n17465), .n17464(n17464), .n17463(n17463), 
            .n17462(n17462), .n17461(n17461), .n17460(n17460), .n17459(n17459), 
            .n17458(n17458), .n17457(n17457), .n17456(n17456), .n17455(n17455), 
            .n17454(n17454), .n17453(n17453), .n17452(n17452), .n17451(n17451), 
            .n17450(n17450), .n17449(n17449), .n17448(n17448), .n17447(n17447), 
            .n17446(n17446), .n17445(n17445), .n17444(n17444), .data_o({quadA_debounced_adj_3970, 
            quadB_debounced_adj_3971}), .GND_net(GND_net), .n2571({n2572, 
            n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
            n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
            n2589, n2590, n2591, n2592, n2593, n2594, n2595}), 
            .count_enable(count_enable_adj_3972), .n16906(n16906), .n17479(n17479), 
            .reg_B({reg_B_adj_4409}), .n31841(n31841), .PIN_7_c_1(PIN_7_c_1), 
            .PIN_6_c_0(PIN_6_c_0), .n16918(n16918)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(218[15] 223[4])
    SB_LUT4 div_43_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4157));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_i723_3_lut_3_lut (.I0(n1067), .I1(n6562), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i26837_3_lut_4_lut (.I0(n15495), .I1(n15501), .I2(n3761), 
            .I3(n740), .O(n32471));
    defparam i26837_3_lut_4_lut.LUT_INIT = 16'hfca8;
    SB_LUT4 i28965_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n34602));
    defparam i28965_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4159));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28971_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n34608));
    defparam i28971_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12682_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17069));   // verilog/coms.v(126[12] 289[6])
    defparam i12682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4161));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12683_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17070));   // verilog/coms.v(126[12] 289[6])
    defparam i12683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4174));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28945_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n34582));
    defparam i28945_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4176));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4178));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28949_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n34586));
    defparam i28949_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12684_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17071));   // verilog/coms.v(126[12] 289[6])
    defparam i12684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i722_3_lut_3_lut (.I0(n1067), .I1(n6561), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12685_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17072));   // verilog/coms.v(126[12] 289[6])
    defparam i12685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12686_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17073));   // verilog/coms.v(126[12] 289[6])
    defparam i12686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4195));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12687_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17074));   // verilog/coms.v(126[12] 289[6])
    defparam i12687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28923_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n34560));
    defparam i28923_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12688_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17075));   // verilog/coms.v(126[12] 289[6])
    defparam i12688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4197));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4199));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12689_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17076));   // verilog/coms.v(126[12] 289[6])
    defparam i12689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28927_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n34564));
    defparam i28927_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4213));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28888_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n34525));
    defparam i28888_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4215));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4217));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28867_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n34504));
    defparam i28867_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4219));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_i724_3_lut_3_lut (.I0(n1067), .I1(n6563), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4235));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28852_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n34489));
    defparam i28852_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12700_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n12917), .I3(GND_net), .O(n17087));   // verilog/coms.v(126[12] 289[6])
    defparam i12700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12701_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n12917), .I3(GND_net), .O(n17088));   // verilog/coms.v(126[12] 289[6])
    defparam i12701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12702_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n12917), .I3(GND_net), .O(n17089));   // verilog/coms.v(126[12] 289[6])
    defparam i12702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12703_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n12917), .I3(GND_net), .O(n17090));   // verilog/coms.v(126[12] 289[6])
    defparam i12703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12704_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n12917), .I3(GND_net), .O(n17091));   // verilog/coms.v(126[12] 289[6])
    defparam i12704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12705_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n12917), .I3(GND_net), .O(n17092));   // verilog/coms.v(126[12] 289[6])
    defparam i12705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12706_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n12917), .I3(GND_net), .O(n17093));   // verilog/coms.v(126[12] 289[6])
    defparam i12706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12707_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n12917), .I3(GND_net), .O(n17094));   // verilog/coms.v(126[12] 289[6])
    defparam i12707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12708_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n12917), .I3(GND_net), .O(n17095));   // verilog/coms.v(126[12] 289[6])
    defparam i12708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12709_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n12917), .I3(GND_net), .O(n17096));   // verilog/coms.v(126[12] 289[6])
    defparam i12709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12710_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n12917), .I3(GND_net), .O(n17097));   // verilog/coms.v(126[12] 289[6])
    defparam i12710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12711_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n12917), .I3(GND_net), .O(n17098));   // verilog/coms.v(126[12] 289[6])
    defparam i12711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12712_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n12917), .I3(GND_net), .O(n17099));   // verilog/coms.v(126[12] 289[6])
    defparam i12712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12713_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n12917), .I3(GND_net), .O(n17100));   // verilog/coms.v(126[12] 289[6])
    defparam i12713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12714_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n12917), .I3(GND_net), .O(n17101));   // verilog/coms.v(126[12] 289[6])
    defparam i12714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12715_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n12917), .I3(GND_net), .O(n17102));   // verilog/coms.v(126[12] 289[6])
    defparam i12715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12716_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n12917), .I3(GND_net), .O(n17103));   // verilog/coms.v(126[12] 289[6])
    defparam i12716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12717_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n12917), .I3(GND_net), .O(n17104));   // verilog/coms.v(126[12] 289[6])
    defparam i12717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12718_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n12917), .I3(GND_net), .O(n17105));   // verilog/coms.v(126[12] 289[6])
    defparam i12718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12719_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n12917), .I3(GND_net), .O(n17106));   // verilog/coms.v(126[12] 289[6])
    defparam i12719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12720_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n12917), .I3(GND_net), .O(n17107));   // verilog/coms.v(126[12] 289[6])
    defparam i12720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12721_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n12917), .I3(GND_net), .O(n17108));   // verilog/coms.v(126[12] 289[6])
    defparam i12721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12722_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n12917), .I3(GND_net), .O(n17109));   // verilog/coms.v(126[12] 289[6])
    defparam i12722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12723_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n12917), .I3(GND_net), .O(n17110));   // verilog/coms.v(126[12] 289[6])
    defparam i12723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12724_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n12917), .I3(GND_net), .O(n17111));   // verilog/coms.v(126[12] 289[6])
    defparam i12724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12725_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n12917), .I3(GND_net), .O(n17112));   // verilog/coms.v(126[12] 289[6])
    defparam i12725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12726_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n12917), .I3(GND_net), .O(n17113));   // verilog/coms.v(126[12] 289[6])
    defparam i12726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12727_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n12917), .I3(GND_net), .O(n17114));   // verilog/coms.v(126[12] 289[6])
    defparam i12727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12728_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n12917), .I3(GND_net), .O(n17115));   // verilog/coms.v(126[12] 289[6])
    defparam i12728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12729_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n12917), .I3(GND_net), .O(n17116));   // verilog/coms.v(126[12] 289[6])
    defparam i12729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12730_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n12917), .I3(GND_net), .O(n17117));   // verilog/coms.v(126[12] 289[6])
    defparam i12730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12731_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n12917), .I3(GND_net), .O(n17118));   // verilog/coms.v(126[12] 289[6])
    defparam i12731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12732_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n12917), .I3(GND_net), .O(n17119));   // verilog/coms.v(126[12] 289[6])
    defparam i12732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4237));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4239));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28838_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n34475));
    defparam i28838_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4241));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4257));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28821_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n34458));
    defparam i28821_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4259));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4261));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28804_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n34441));
    defparam i28804_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4263));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636_adj_4012), 
            .I3(GND_net), .O(n10_adj_4279));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633_adj_4009), 
            .I3(GND_net), .O(n14_adj_4283));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28752_2_lut_4_lut (.I0(n2623_adj_3999), .I1(n84), .I2(n2632_adj_4008), 
            .I3(n93), .O(n34389));
    defparam i28752_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623_adj_3999), 
            .I3(GND_net), .O(n16_adj_4285));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631_adj_4007), 
            .I3(GND_net), .O(n12_adj_4281));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28784_2_lut_4_lut (.I0(n2631_adj_4007), .I1(n92), .I2(n2635_adj_4011), 
            .I3(n96), .O(n34421));
    defparam i28784_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15502), .I1(r_SM_Main_2__N_3259[0]), .I2(tx_active), 
            .I3(n22044), .O(n31_adj_4358));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 div_43_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4303));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4301));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_43_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4305));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28788_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n34425));
    defparam i28788_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4307));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28723_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n34360));
    defparam i28723_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_43_i720_3_lut_3_lut (.I0(n1067), .I1(n6559), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i725_3_lut_3_lut (.I0(n1067), .I1(n6564), .I2(n374), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_25_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3934));   // verilog/TinyFPGA_B.v(128[23:28])
    defparam unary_minus_25_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29123_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29123_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_43_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2), .I3(n5_adj_4356), 
            .O(n30813));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_43_i721_3_lut_3_lut (.I0(n1067), .I1(n6560), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i29099_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n370), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29099_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_43_i719_3_lut_3_lut (.I0(n1067), .I1(n6558), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_43_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_3938), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_43_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_3967), 
            .I3(n30813), .O(n30817));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i29090_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n371), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29090_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_43_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_3940), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_43_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15430), 
            .O(n249));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_43_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_3939), 
            .I3(n30817), .O(n30819));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n17442(n17442), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n17441(n17441), .n17440(n17440), .n17439(n17439), 
            .n17438(n17438), .n17437(n17437), .n17436(n17436), .n17435(n17435), 
            .n17434(n17434), .n17433(n17433), .n17432(n17432), .n17431(n17431), 
            .n17430(n17430), .n17429(n17429), .n17428(n17428), .n17427(n17427), 
            .n17426(n17426), .n17425(n17425), .n17424(n17424), .n17423(n17423), 
            .n17422(n17422), .n17421(n17421), .n17420(n17420), .data_o({quadA_debounced, 
            quadB_debounced}), .n2621({n2622, n2623, n2624, n2625, 
            n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
            n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
            n2642, n2643, n2644, n2645}), .GND_net(GND_net), .count_enable(count_enable), 
            .n16904(n16904), .n17467(n17467), .reg_B({reg_B}), .n31114(n31114), 
            .PIN_2_c_1(PIN_2_c_1), .PIN_1_c_0(PIN_1_c_0), .n16907(n16907)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(210[15] 215[4])
    SB_LUT4 i1_2_lut_4_lut_adj_1609 (.I0(n98), .I1(n97), .I2(n96), .I3(n15439), 
            .O(n15430));
    defparam i1_2_lut_4_lut_adj_1609.LUT_INIT = 16'hff7f;
    SB_LUT4 div_43_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2_adj_3941), 
            .I3(n649), .O(n784));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i1_2_lut_3_lut_adj_1610 (.I0(n97), .I1(n96), .I2(n15439), 
            .I3(GND_net), .O(n15433));
    defparam i1_2_lut_3_lut_adj_1610.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1611 (.I0(n95), .I1(n94), .I2(n93), .I3(n15448), 
            .O(n15439));
    defparam i1_2_lut_4_lut_adj_1611.LUT_INIT = 16'hff7f;
    SB_LUT4 i29078_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n372), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i29078_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i1_2_lut_3_lut_adj_1612 (.I0(n94), .I1(n93), .I2(n15448), 
            .I3(GND_net), .O(n15442));
    defparam i1_2_lut_3_lut_adj_1612.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1613 (.I0(n92), .I1(n91), .I2(n90), .I3(n15457), 
            .O(n15448));
    defparam i1_2_lut_4_lut_adj_1613.LUT_INIT = 16'hff7f;
    SB_LUT4 div_43_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4355), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_43_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_3936), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i1_2_lut_3_lut_adj_1614 (.I0(n91), .I1(n90), .I2(n15457), 
            .I3(GND_net), .O(n15451));
    defparam i1_2_lut_3_lut_adj_1614.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1615 (.I0(n89), .I1(n88), .I2(n87), .I3(n15466), 
            .O(n15457));
    defparam i1_2_lut_4_lut_adj_1615.LUT_INIT = 16'hff7f;
    SB_LUT4 div_43_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_3973), 
            .I3(n30819), .O(n914));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 i1_2_lut_3_lut_adj_1616 (.I0(n88), .I1(n87), .I2(n15466), 
            .I3(GND_net), .O(n15460));
    defparam i1_2_lut_3_lut_adj_1616.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1617 (.I0(n86), .I1(n85), .I2(n84), .I3(n15475), 
            .O(n15466));
    defparam i1_2_lut_4_lut_adj_1617.LUT_INIT = 16'hff7f;
    SB_LUT4 i12733_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n12917), .I3(GND_net), .O(n17120));   // verilog/coms.v(126[12] 289[6])
    defparam i12733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12734_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n12917), .I3(GND_net), .O(n17121));   // verilog/coms.v(126[12] 289[6])
    defparam i12734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12735_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n12917), .I3(GND_net), .O(n17122));   // verilog/coms.v(126[12] 289[6])
    defparam i12735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12736_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n12917), .I3(GND_net), .O(n17123));   // verilog/coms.v(126[12] 289[6])
    defparam i12736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4019), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_43_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4075));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1618 (.I0(n85), .I1(n84), .I2(n15475), 
            .I3(GND_net), .O(n15469));
    defparam i1_2_lut_3_lut_adj_1618.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1619 (.I0(n83), .I1(n82), .I2(n81), .I3(n15484), 
            .O(n15475));
    defparam i1_2_lut_4_lut_adj_1619.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1620 (.I0(n82), .I1(n81), .I2(n15484), 
            .I3(GND_net), .O(n15478));
    defparam i1_2_lut_3_lut_adj_1620.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1621 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n15484));
    defparam i1_2_lut_4_lut_adj_1621.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1622 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n15487));
    defparam i1_2_lut_3_lut_adj_1622.LUT_INIT = 16'hf7f7;
    SB_LUT4 i20015_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_3967));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20015_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i20039_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4_adj_3940));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20039_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i20071_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4355));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam i20071_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i12737_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n12917), .I3(GND_net), .O(n17124));   // verilog/coms.v(126[12] 289[6])
    defparam i12737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12738_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n12917), .I3(GND_net), .O(n17125));   // verilog/coms.v(126[12] 289[6])
    defparam i12738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12739_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n12917), .I3(GND_net), .O(n17126));   // verilog/coms.v(126[12] 289[6])
    defparam i12739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_43_i636_3_lut_3_lut (.I0(n938), .I1(n6552), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(206[21:53])
    defparam div_43_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    \pwm(32000000,20000,32000000,23,1)  PWM (.pwm_setpoint({pwm_setpoint}), 
            .\half_duty_new[0] (half_duty_new[0]), .CLK_c(CLK_c), .PIN_19_c_0(PIN_19_c_0), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n925(n925), .\half_duty[0][1] (\half_duty[0] [1]), 
            .n17487(n17487), .\half_duty[0][7] (\half_duty[0] [7]), .n17486(n17486), 
            .\half_duty[0][6] (\half_duty[0] [6]), .n17485(n17485), .\half_duty[0][5] (\half_duty[0] [5]), 
            .n17484(n17484), .\half_duty[0][4] (\half_duty[0] [4]), .n17483(n17483), 
            .\half_duty[0][3] (\half_duty[0] [3]), .n17482(n17482), .\half_duty[0][2] (\half_duty[0] [2]), 
            .n17481(n17481), .\half_duty_new[7] (half_duty_new[7]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[5] (half_duty_new[5]), .\half_duty_new[4] (half_duty_new[4]), 
            .\half_duty_new[3] (half_duty_new[3]), .\half_duty_new[2] (half_duty_new[2]), 
            .\half_duty_new[1] (half_duty_new[1]), .\half_duty[0][0] (\half_duty[0] [0]), 
            .n16936(n16936)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(110[43] 116[3])
    motorControl control (.\Kp[1] (Kp[1]), .GND_net(GND_net), .\Kp[0] (Kp[0]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .PWMLimit({PWMLimit}), .setpoint({setpoint}), 
            .duty({duty}), .clk32MHz(clk32MHz), .motor_state({motor_state}), 
            .VCC_net(VCC_net), .n36858(n36858)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(190[16] 203[4])
    SB_LUT4 i12740_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n12917), .I3(GND_net), .O(n17127));   // verilog/coms.v(126[12] 289[6])
    defparam i12740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12741_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n12917), .I3(GND_net), .O(n17128));   // verilog/coms.v(126[12] 289[6])
    defparam i12741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12742_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n12917), .I3(GND_net), .O(n17129));   // verilog/coms.v(126[12] 289[6])
    defparam i12742_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (timer, GND_net, \neo_pixel_transmitter.done , clk32MHz, 
            n29069, VCC_net, bit_ctr, \neo_pixel_transmitter.t0 , n29137, 
            n29135, n29133, n29131, n29129, n29127, n29125, n29123, 
            n29121, n29119, n29117, n29115, n29113, n29111, n29109, 
            n29107, n29105, n29103, n29097, n29095, n29093, n29091, 
            n29089, n29085, n29083, n29071, n29073, n29075, n34308, 
            n19, n34303, \state[0] , \state[1] , start, n34301, 
            n34295, n34294, n34293, n34307, n34292, n34302, n34288, 
            n34323, n34322, n34320, n34296, n34319, n34291, n34318, 
            n34290, n34317, \state_3__N_298[1] , n15387, n919, n4404, 
            \color[18] , \color[19] , n34321, \color[17] , \color[16] , 
            n34289, n34316, n34305, n34306, n34315, n34314, n34313, 
            n34304, n34312, n16527, n30957, n34311, PIN_8_c, n29087, 
            n16771, n29081, n17005, n17004, n17003, n17002, n17001, 
            n17000, n16999, n16998, n16997, n16996, n16995, n16994, 
            n16993, n16992, n16991, n16990, n16989, n16988, n16987, 
            n16986, n16985, n16983, n16982, n16981, n16980, n16979, 
            n16978, n16977, n16976, n16975, n16974, n29079, n16923, 
            n34310, n29077, n34309, n22030, n29225, \color[22] , 
            \color[23] , \color[21] , \color[20] , n22016) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [31:0]timer;
    input GND_net;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    input n29069;
    input VCC_net;
    output [31:0]bit_ctr;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n29137;
    input n29135;
    input n29133;
    input n29131;
    input n29129;
    input n29127;
    input n29125;
    input n29123;
    input n29121;
    input n29119;
    input n29117;
    input n29115;
    input n29113;
    input n29111;
    input n29109;
    input n29107;
    input n29105;
    input n29103;
    input n29097;
    input n29095;
    input n29093;
    input n29091;
    input n29089;
    input n29085;
    input n29083;
    input n29071;
    input n29073;
    input n29075;
    output n34308;
    input n19;
    output n34303;
    output \state[0] ;
    output \state[1] ;
    output start;
    output n34301;
    output n34295;
    output n34294;
    output n34293;
    output n34307;
    output n34292;
    output n34302;
    output n34288;
    output n34323;
    output n34322;
    output n34320;
    output n34296;
    output n34319;
    output n34291;
    output n34318;
    output n34290;
    output n34317;
    output \state_3__N_298[1] ;
    output n15387;
    output n919;
    output n4404;
    input \color[18] ;
    input \color[19] ;
    output n34321;
    input \color[17] ;
    input \color[16] ;
    output n34289;
    output n34316;
    output n34305;
    output n34306;
    output n34315;
    output n34314;
    output n34313;
    output n34304;
    output n34312;
    output n16527;
    output n30957;
    output n34311;
    output PIN_8_c;
    input n29087;
    input n16771;
    input n29081;
    input n17005;
    input n17004;
    input n17003;
    input n17002;
    input n17001;
    input n17000;
    input n16999;
    input n16998;
    input n16997;
    input n16996;
    input n16995;
    input n16994;
    input n16993;
    input n16992;
    input n16991;
    input n16990;
    input n16989;
    input n16988;
    input n16987;
    input n16986;
    input n16985;
    input n16983;
    input n16982;
    input n16981;
    input n16980;
    input n16979;
    input n16978;
    input n16977;
    input n16976;
    input n16975;
    input n16974;
    input n29079;
    input n16923;
    output n34310;
    input n29077;
    output n34309;
    output n22030;
    output n29225;
    input \color[22] ;
    input \color[23] ;
    input \color[21] ;
    input \color[20] ;
    output n22016;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n24815;
    wire [31:0]n1;
    
    wire n24816, n25436, n1999, n2027, n25437, n28, n24814;
    wire [31:0]one_wire_N_449;
    
    wire n2099, n2000, n25435, n21, n24813, n2100, n2001, n25434;
    wire [31:0]n133;
    
    wire n25493, n27, n24812, \neo_pixel_transmitter.done_N_506 , n37051, 
        n2101, n2002, n25433, n2102, n2003, n25432, n2103, n2004, 
        n25431, n25494, n30, n24811, n29, n24810, n2104, n2005, 
        n25430, n25492, n25491, n25, n24809, n2105, n2006, n25429, 
        n2106, n2007, n25428, n25490, n2107, n2008, n25427, n24, 
        n24808, n2108, n2009, n36857, n25426, n2109, n2192, n2093, 
        n2126, n25425, n2193, n2094, n25424, n2194, n2095, n25423, 
        n25489, n2195, n2096, n25422, n2196, n2097, n25421, n24807, 
        n2197, n2098, n25420, n25488, n25487, n2198, n25419, n25486, 
        n2199, n25418, n2200, n25417, n2201, n25416, n2202, n25415, 
        n2203, n25414, n2204, n25413, n2205, n25412, n2206, n25411, 
        n2207, n25410, n24806, n2208, n36859, n25409, n2209, n2291, 
        n2225, n25408, n2292, n25407, n2293, n25406, n2294, n25405, 
        n2295, n25404, n2296, n25403, n25485, n24618, n2297, n25402, 
        n25484, n2298, n25401, n24610, n25483, n2299, n25400, 
        n2300, n25399, n2301, n25398, n25482, n2324, n36861, n24805, 
        n1806, n1803, n1798, n1805, n24_adj_3804, n1808, n1804, 
        n1802, n1807, n22_adj_3805, n1800, n1799, n1797, n1801, 
        n23_adj_3806, n1796, n1809, n21_adj_3807, n1829, n24619, 
        n2302, n25397, n22_adj_3810, n2309, n30_adj_3811, n2306, 
        n34, n2307, n2305, n32, n2304, n33, n2308, n2303, n31_adj_3812, 
        n25396, n24804, n25395, n25394, n25481, n25393, n24803, 
        n25392, n36860, n25391, n25480, n24611, n2390, n25390, 
        n2391, n25389, n2392, n25388, n25479, n2393, n25387, n24802, 
        n23_adj_3815, n22_adj_3816, n36, n26_adj_3817, n37, n15393, 
        n30197, n24801, n25478, n2394, n25386, n24800, n2395, 
        n25385, n26076, n111, n116, n1895, n25477, n2396, n25384, 
        n24799, n2397, n25383, n1896, n25476, n2398, n25382, n1897, 
        n25475, n2399, n25381, n1898, n25474, n2400, n25380, n2401, 
        n25379, n2402, n25378, n2403, n25377, n2404, n25376, n2405, 
        n25375, n1899, n25473, n24798, n1900, n25472, n2406, n25374, 
        n1901, n25471, n2407, n25373, n18_adj_3818, n2408, n25372, 
        n1902, n25470, n807, n14115, n30829, n838, n1903, n25469, 
        n2409, n1904, n25468, n1905, n25467, n24797, n30953, n24796, 
        n4, n1906, n25466, n20_adj_3821, n1907, n25465, n24638, 
        n1908, n36862, n25464, n1909, n24637, n7, n24636, n1928, 
        n36865, n24635, n24617, n24634, n24609, n2489, n2423, 
        n25304, n2490, n25303, n2491, n25302, n2492, n25301, n2493, 
        n25300, n1994, n25456, n2494, n25299, n2495, n25298, n1995, 
        n25455, n2496, n25297, n36864, n2497, n25296, n2498, n25295, 
        n2499, n25294, n2500, n25293, n24633, n1996, n25454, n2501, 
        n25292, n2502, n25291, n2503, n25290, n1997, n25453, n26_adj_3822, 
        n19_adj_3823, n16_adj_3824, n24_adj_3825, n28_adj_3826, n2504, 
        n25289, n2505, n25288, n27_adj_3827, n33_adj_3828, n32_adj_3829, 
        n31_adj_3830, n35, n37_adj_3831, n2506, n25287, n2507, n25286, 
        n1998, n25452, n28_adj_3832, n31_adj_3833, n22_adj_3834, n30_adj_3835, 
        n34_adj_3836, n21_adj_3837, n2508, n25285, n2509, n25451, 
        n24632, n24631, n24630, n24616, n25450, n25449, n25448, 
        n25447, n25446, n24629, n25445, n25444, n25443, n25442, 
        n24615, n24628, n24614, n24627, n18_adj_3838, n21839, n30_adj_3839, 
        n28_adj_3840, n29_adj_3841, n27_adj_3842, n25921, n30886, 
        n15386, n10, n14_adj_3843, n15289, n30_adj_3844, n48, n46, 
        n47, n45, n44, n43, n54, n49, n4377, n36990, n24608, 
        n36993, n24613, n2588, n2522, n25179, n2589, n25178, n2590, 
        n25177, n2591, n25176, n2592, n25175, n2593, n25174, n2594, 
        n25173, n2595, n25172, n2596, n25171, n2597, n25170, n2598, 
        n25169, n2599, n25168, n2600, n25167, n24626, n2601, n25166, 
        n2602, n25165, n2603, n25164, n2604, n25163, n2605, n25162, 
        n2606, n25161, n24612, n2607, n25160, n2608, n36866, n25159, 
        n24625, n2609, n24624, n24623, n24622, n24826, n24825;
    wire [3:0]state_3__N_298;
    
    wire n24621, n24824, n2687, n2621, n25119, n2688, n25118, 
        n2689, n25117, n2690, n25116, n2691, n25115, n2692, n25114, 
        n2693, n25113, n2694, n25112, n2695, n25111, n2696, n25110, 
        n2697, n25109, n2698, n25108, n2699, n25107, n2700, n25106, 
        n2701, n25105, n2702, n25104, n2703, n25103, n2704, n25102, 
        n2705, n25101, n2706, n25100, n2707, n25099, n2708, n36867, 
        n25098, n2709, n2786, n2720, n25067, n2787, n25066, n2788, 
        n25065, n2789, n25064, n2790, n25063, n2791, n25062, n2792, 
        n25061, n2793, n25060, n2794, n25059, n2795, n25058, n2796, 
        n25057, n2797, n25056, n2798, n25055, n2799, n25054, n2800, 
        n25053, n2801, n25052, n2802, n25051, n2803, n25050, n2804, 
        n25049, n2805, n25048, n2806, n25047, n2807, n25046, n2808, 
        n36868, n25045, n2809, n2885, n2819, n25029, n2886, n25028, 
        n2887, n25027, n2888, n25026, n2889, n25025, n2890, n25024, 
        n2891, n25023, n2892, n25022, n2893, n25021, n2894, n25020, 
        n2895, n25019, n2896, n25018, n2897, n25017, n2898, n25016, 
        n2899, n25015, n2900, n25014, n2901, n25013, n2902, n25012, 
        n2903, n25011, n2904, n25010, n2905, n25009, n2906, n25008, 
        n2907, n25007, n2908, n36869, n25006, n2909, \neo_pixel_transmitter.done_N_512 , 
        n31011, n32288, n2984, n2918, n24994, n2985, n24993, n2986, 
        n24992, n2987, n24991, n2988, n24990, n2989, n24989, n2990, 
        n24988, n2991, n24987, n2992, n24986, n2993, n24985, n2994, 
        n24984, n24823, n2995, n24983, n2996, n24982, n2997, n24981, 
        n2998, n24980, n2999, n24979, n3000, n24978, n3001, n24977, 
        n3002, n24976, n3003, n24975, n3004, n24974, n3005, n24973, 
        n3006, n24972;
    wire [31:0]n971;
    
    wire n905, n25645, n906, n25644, n25643, n16628, n25642, n3007, 
        n24971, n14113, n25641, n1103, n4_adj_3846, n1037, n25640, 
        n1104, n1005, n25639, n3008, n36870, n24970, n1105, n1006, 
        n25638, n3009, n1106, n1007, n25637, n3083, n3017, n24969, 
        n1107, n1008, n25636, n3084, n24968, n1108, n1009, n36871, 
        n25635, n3085, n24967, n25441, n1109, n3086, n24966, n24822, 
        n1202, n1136, n25634, n1203, n25633, n1204, n25632, n3087, 
        n24965, n1205, n25631, n1206, n25630, n1207, n25629, n1208, 
        n36873, n25628, n1209, n1301, n1235, n25627, n1302, n25626, 
        n1303, n25625, n1304, n25624, n1305, n25623, n1306, n25622, 
        n1307, n25621, n3088, n24964, n25440, n1308, n36874, n25620, 
        n3089, n24963, n1309, n1400, n1334, n25619, n3090, n24962, 
        n1401, n25618, n3091, n24961, n3092, n24960, n3093, n24959, 
        n25439, n24821, n1402, n25617, n1403, n25616, n3094, n24958, 
        n25438, n3095, n24957, n3096, n24956, n24820, n3097, n24955, 
        n3098, n24954, n3099, n24953, n1404, n25615, n3100, n24952, 
        n1405, n25614, n3101, n24951, n1406, n25613, n1407, n25612, 
        n1408, n36875, n25611, n3102, n24950, n1409, n1499, n1433, 
        n25610, n1500, n25609, n1501, n25608, n1502, n25607, n3103, 
        n24949, n1503, n25606, n3104, n24948, n1504, n25605, n1505, 
        n25604, n1506, n25603, n1507, n25602, n1508, n36876, n25601, 
        n1509, n1598, n1532, n25600, n1599, n25599, n3105, n24947, 
        n1600, n25598, n1601, n25597, n1602, n25596, n1603, n25595, 
        n1604, n25594, n1605, n25593, n1606, n25592, n1607, n25591, 
        n1608, n36877, n25590, n1609, n3106, n24946, n3107, n24945, 
        n3108, n36872, n24944, n3109, n24620, n3182, n3116, n24943, 
        n3183, n24942, n3184, n24941, n3185, n24940, n3186, n24939, 
        n24819, n3187, n24938, n3188, n24937, n3189, n24936, n1697, 
        n1631, n25543, n3190, n24935, n1698, n25542, n24818, n1699, 
        n25541, n3191, n24934, n1700, n25540, n3192, n24933, n1701, 
        n25539, n1702, n25538, n3193, n24932, n1703, n25537, n1704, 
        n25536, n1705, n25535, n1706, n25534, n3194, n24931, n1707, 
        n25533, n1708, n36879, n25532, n1709, n1730, n25531, n25530, 
        n25529, n25528, n25527, n25526, n3195, n24930, n25525, 
        n25524, n25523, n3196, n24929, n3197, n24928, n25522, 
        n25521, n25520, n3198, n24927, n36880, n25519, n3199, 
        n24926, n3200, n24925, n24817, n3201, n24924, n3202, n24923, 
        n3203, n24922, n3204, n24921, n3205, n24920, n3206, n24919, 
        n3207, n24918, n3208, n36878, n24917, n3209, n25508, n25507, 
        n25506, n25505, n25504, n25503, n25502, n25501, n25500, 
        n25499, n25498, n25497, n25496, n25495, n18_adj_3849, n28_adj_3850, 
        n26_adj_3851, n17_adj_3852, n21_adj_3853, n20_adj_3854, n24_adj_3855, 
        n27_adj_3856, n20_adj_3857, n13_adj_3858, n18_adj_3859, n22_adj_3860, 
        n36_adj_3861, n46_adj_3862, n42, n44_adj_3863, n31_adj_3864, 
        n50, n48_adj_3865, n49_adj_3866, n47_adj_3867, n18_adj_3868, 
        n16_adj_3869, n20_adj_3870, n31001, n7_adj_3871, n21950, n16_adj_3872, 
        n17_adj_3873, n36894, n36897, n708, n26372, n10_adj_3874, 
        n12_adj_3875, n16_adj_3876, n14_adj_3877, n9_adj_3878, n30800, 
        n34325, n21964, n12_adj_3879, n35417, n35418, n40, n44_adj_3880, 
        n42_adj_3881, n43_adj_3882, n41, n38, n46_adj_3883, n50_adj_3884, 
        n37_adj_3885, n27151, n739, n8_adj_3886, n32529, n6_adj_3887, 
        n60, n30837, n33_adj_3888, n41_adj_3889, n38_adj_3890, n43_adj_3891, 
        n40_adj_3892, n46_adj_3893, n39, n47_adj_3894, n30888, n30997, 
        n40_adj_3895, n38_adj_3896, n39_adj_3897, n37_adj_3898, n34_adj_3899, 
        n42_adj_3900, n46_adj_3901, n33_adj_3902, n28_adj_3903, n38_adj_3904, 
        n21876, n36_adj_3905, n42_adj_3906, n40_adj_3907, n41_adj_3908, 
        n39_adj_3909, n36_adj_3910, n25_adj_3911, n34_adj_3912, n40_adj_3913, 
        n38_adj_3914, n39_adj_3915, n37_adj_3916, n21940, n48_adj_3917, 
        n46_adj_3918, n47_adj_3919, n45_adj_3920, n44_adj_3921, n43_adj_3922, 
        n54_adj_3923, n49_adj_3924, n21992, n922, n5_adj_3925, n25_adj_3926, 
        n24_adj_3927, n34_adj_3928, n22_adj_3929, n38_adj_3930, n36_adj_3931, 
        n37_adj_3932, n35_adj_3933;
    
    SB_CARRY sub_14_add_2_22 (.CI(n24815), .I0(timer[20]), .I1(n1[20]), 
            .CO(n24816));
    SB_CARRY mod_5_add_1406_13 (.CI(n25436), .I0(n1999), .I1(n2027), .CO(n25437));
    SB_LUT4 sub_14_add_2_21_lut (.I0(one_wire_N_449[29]), .I1(timer[19]), 
            .I2(n1[19]), .I3(n24814), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n25435), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n25435), .I0(n2000), .I1(n2027), .CO(n25436));
    SB_CARRY sub_14_add_2_21 (.CI(n24814), .I0(timer[19]), .I1(n1[19]), 
            .CO(n24815));
    SB_LUT4 sub_14_add_2_20_lut (.I0(one_wire_N_449[27]), .I1(timer[18]), 
            .I2(n1[18]), .I3(n24813), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n25434), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n25493), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n24813), .I0(timer[18]), .I1(n1[18]), 
            .CO(n24814));
    SB_CARRY mod_5_add_1406_11 (.CI(n25434), .I0(n2001), .I1(n2027), .CO(n25435));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_449[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n24812), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n37051), .D(\neo_pixel_transmitter.done_N_506 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_19 (.CI(n24812), .I0(timer[17]), .I1(n1[17]), 
            .CO(n24813));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n25433), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(VCC_net), 
            .D(n29069));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_10 (.CI(n25433), .I0(n2002), .I1(n2027), .CO(n25434));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n25432), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n25432), .I0(n2003), .I1(n2027), .CO(n25433));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n25431), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n25431), .I0(n2004), .I1(n2027), .CO(n25432));
    SB_CARRY timer_1129_add_4_18 (.CI(n25493), .I0(GND_net), .I1(timer[16]), 
            .CO(n25494));
    SB_LUT4 sub_14_add_2_18_lut (.I0(one_wire_N_449[23]), .I1(timer[16]), 
            .I2(n1[16]), .I3(n24811), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n24811), .I0(timer[16]), .I1(n1[16]), 
            .CO(n24812));
    SB_LUT4 sub_14_add_2_17_lut (.I0(one_wire_N_449[20]), .I1(timer[15]), 
            .I2(n1[15]), .I3(n24810), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n25430), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n25492), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n24810), .I0(timer[15]), .I1(n1[15]), 
            .CO(n24811));
    SB_CARRY timer_1129_add_4_17 (.CI(n25492), .I0(GND_net), .I1(timer[15]), 
            .CO(n25493));
    SB_CARRY mod_5_add_1406_7 (.CI(n25430), .I0(n2005), .I1(n2027), .CO(n25431));
    SB_LUT4 timer_1129_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n25491), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_16 (.CI(n25491), .I0(GND_net), .I1(timer[14]), 
            .CO(n25492));
    SB_LUT4 sub_14_add_2_16_lut (.I0(one_wire_N_449[21]), .I1(timer[14]), 
            .I2(n1[14]), .I3(n24809), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n25429), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n25429), .I0(n2006), .I1(n2027), .CO(n25430));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n25428), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n25490), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_15 (.CI(n25490), .I0(GND_net), .I1(timer[13]), 
            .CO(n25491));
    SB_CARRY mod_5_add_1406_5 (.CI(n25428), .I0(n2007), .I1(n2027), .CO(n25429));
    SB_CARRY sub_14_add_2_16 (.CI(n24809), .I0(timer[14]), .I1(n1[14]), 
            .CO(n24810));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n25427), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_15_lut (.I0(one_wire_N_449[22]), .I1(timer[13]), 
            .I2(n1[13]), .I3(n24808), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1406_4 (.CI(n25427), .I0(n2008), .I1(n2027), .CO(n25428));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n36857), 
            .I3(n25426), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_3 (.CI(n25426), .I0(n2009), .I1(n36857), .CO(n25427));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n36857), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n36857), 
            .CO(n25426));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n25425), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_15 (.CI(n24808), .I0(timer[13]), .I1(n1[13]), 
            .CO(n24809));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n25424), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n25424), .I0(n2094), .I1(n2126), .CO(n25425));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n25423), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n25423), .I0(n2095), .I1(n2126), .CO(n25424));
    SB_LUT4 timer_1129_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n25489), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n25422), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n25422), .I0(n2096), .I1(n2126), .CO(n25423));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n25421), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1129_add_4_14 (.CI(n25489), .I0(GND_net), .I1(timer[12]), 
            .CO(n25490));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n24807), .O(one_wire_N_449[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n25421), .I0(n2097), .I1(n2126), .CO(n25422));
    SB_CARRY sub_14_add_2_14 (.CI(n24807), .I0(timer[12]), .I1(n1[12]), 
            .CO(n24808));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n25420), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n25488), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n25420), .I0(n2098), .I1(n2126), .CO(n25421));
    SB_CARRY timer_1129_add_4_13 (.CI(n25488), .I0(GND_net), .I1(timer[11]), 
            .CO(n25489));
    SB_LUT4 timer_1129_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n25487), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_12 (.CI(n25487), .I0(GND_net), .I1(timer[10]), 
            .CO(n25488));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n25419), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n25419), .I0(n2099), .I1(n2126), .CO(n25420));
    SB_LUT4 timer_1129_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n25486), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n25418), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n25418), .I0(n2100), .I1(n2126), .CO(n25419));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n25417), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_11 (.CI(n25417), .I0(n2101), .I1(n2126), .CO(n25418));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n25416), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n25416), .I0(n2102), .I1(n2126), .CO(n25417));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n25415), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n25415), .I0(n2103), .I1(n2126), .CO(n25416));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n25414), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n25414), .I0(n2104), .I1(n2126), .CO(n25415));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n25413), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n25413), .I0(n2105), .I1(n2126), .CO(n25414));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n25412), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n25412), .I0(n2106), .I1(n2126), .CO(n25413));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n25411), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n25411), .I0(n2107), .I1(n2126), .CO(n25412));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n25410), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n29137));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n29135));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n29133));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n29131));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n29129));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n29127));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n29125));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n29123));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n24806), .O(one_wire_N_449[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n29121));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n29119));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n29117));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n29115));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n29113));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n29111));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n29109));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n29107));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n29105));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n29103));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n29097));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n29095));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n29093));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n29091));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n29089));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n29085));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n29083));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(VCC_net), 
            .D(n29071));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(VCC_net), 
            .D(n29073));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(VCC_net), 
            .D(n29075));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_4 (.CI(n25410), .I0(n2108), .I1(n2126), .CO(n25411));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n36859), 
            .I3(n25409), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n25409), .I0(n2109), .I1(n36859), .CO(n25410));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n36859), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n36859), 
            .CO(n25409));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n25408), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n25407), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1129_add_4_11 (.CI(n25486), .I0(GND_net), .I1(timer[9]), 
            .CO(n25487));
    SB_CARRY mod_5_add_1540_19 (.CI(n25407), .I0(n2193), .I1(n2225), .CO(n25408));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n25406), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n25406), .I0(n2194), .I1(n2225), .CO(n25407));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n25405), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n25405), .I0(n2195), .I1(n2225), .CO(n25406));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n25404), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n25404), .I0(n2196), .I1(n2225), .CO(n25405));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n25403), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n25485), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_13_lut (.I0(n19), .I1(bit_ctr[11]), .I2(GND_net), .I3(n24618), 
            .O(n34308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_13 (.CI(n24806), .I0(timer[11]), .I1(n1[11]), 
            .CO(n24807));
    SB_CARRY mod_5_add_1540_15 (.CI(n25403), .I0(n2197), .I1(n2225), .CO(n25404));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n25402), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1129_add_4_10 (.CI(n25485), .I0(GND_net), .I1(timer[8]), 
            .CO(n25486));
    SB_CARRY mod_5_add_1540_14 (.CI(n25402), .I0(n2198), .I1(n2225), .CO(n25403));
    SB_LUT4 timer_1129_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n25484), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n25401), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n25401), .I0(n2199), .I1(n2225), .CO(n25402));
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n24610), 
            .O(n34303)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1129_add_4_9 (.CI(n25484), .I0(GND_net), .I1(timer[7]), 
            .CO(n25485));
    SB_LUT4 timer_1129_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n25483), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_8 (.CI(n25483), .I0(GND_net), .I1(timer[6]), 
            .CO(n25484));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n25400), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n25400), .I0(n2200), .I1(n2225), .CO(n25401));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n25399), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n25399), .I0(n2201), .I1(n2225), .CO(n25400));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n25398), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1129_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n25482), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n25398), .I0(n2202), .I1(n2225), .CO(n25399));
    SB_LUT4 i31224_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36861));
    defparam i31224_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n24805), .O(one_wire_N_449[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_3804));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_3805));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_3806));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21_adj_3807));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut (.I0(n21_adj_3807), .I1(n23_adj_3806), .I2(n22_adj_3805), 
            .I3(n24_adj_3804), .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_12 (.CI(n24805), .I0(timer[10]), .I1(n1[10]), 
            .CO(n24806));
    SB_CARRY add_21_13 (.CI(n24618), .I0(bit_ctr[11]), .I1(GND_net), .CO(n24619));
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n25397), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_3810));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1540_9 (.CI(n25397), .I0(n2203), .I1(n2225), .CO(n25398));
    SB_LUT4 i11_4_lut (.I0(bit_ctr[12]), .I1(n22_adj_3810), .I2(n2299), 
            .I3(n2309), .O(n30_adj_3811));
    defparam i11_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut (.I0(n2294), .I1(n30_adj_3811), .I2(n2306), .I3(n2297), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1413 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32));
    defparam i13_4_lut_adj_1413.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_3812));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31_adj_3812), .I1(n33), .I2(n32), .I3(n34), 
            .O(n2324));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n25396), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_8 (.CI(n25396), .I0(n2204), .I1(n2225), .CO(n25397));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n24804), .O(one_wire_N_449[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n25395), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1129_add_4_7 (.CI(n25482), .I0(GND_net), .I1(timer[5]), 
            .CO(n25483));
    SB_CARRY mod_5_add_1540_7 (.CI(n25395), .I0(n2205), .I1(n2225), .CO(n25396));
    SB_CARRY sub_14_add_2_11 (.CI(n24804), .I0(timer[9]), .I1(n1[9]), 
            .CO(n24805));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n25394), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n25394), .I0(n2206), .I1(n2225), .CO(n25395));
    SB_LUT4 timer_1129_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n25481), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n25393), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n25393), .I0(n2207), .I1(n2225), .CO(n25394));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n24803), .O(one_wire_N_449[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n25392), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n25392), .I0(n2208), .I1(n2225), .CO(n25393));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n36860), 
            .I3(n25391), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n25391), .I0(n2209), .I1(n36860), .CO(n25392));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n36860), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1129_add_4_6 (.CI(n25481), .I0(GND_net), .I1(timer[4]), 
            .CO(n25482));
    SB_LUT4 timer_1129_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n25480), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_5 (.CI(n25480), .I0(GND_net), .I1(timer[3]), 
            .CO(n25481));
    SB_CARRY add_21_5 (.CI(n24610), .I0(bit_ctr[3]), .I1(GND_net), .CO(n24611));
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n36860), 
            .CO(n25391));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n25390), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n24803), .I0(timer[8]), .I1(n1[8]), 
            .CO(n24804));
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n25389), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n25389), .I0(n2292), .I1(n2324), .CO(n25390));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n25388), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n25388), .I0(n2293), .I1(n2324), .CO(n25389));
    SB_LUT4 timer_1129_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n25479), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n25387), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n24802), .O(one_wire_N_449[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_4 (.CI(n25479), .I0(GND_net), .I1(timer[2]), 
            .CO(n25480));
    SB_CARRY mod_5_add_1607_18 (.CI(n25387), .I0(n2294), .I1(n2324), .CO(n25388));
    SB_LUT4 i16_4_lut (.I0(n21), .I1(n23_adj_3815), .I2(n22_adj_3816), 
            .I3(n24), .O(n36));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_9 (.CI(n24802), .I0(timer[7]), .I1(n1[7]), .CO(n24803));
    SB_LUT4 i17_4_lut (.I0(n25), .I1(n27), .I2(n26_adj_3817), .I3(n28), 
            .O(n37));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n29), .I2(n36), .I3(n30), .O(n15393));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30522_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n30197));
    defparam i30522_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n24801), .O(one_wire_N_449[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1129_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n25478), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n25386), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_8 (.CI(n24801), .I0(timer[6]), .I1(n1[6]), .CO(n24802));
    SB_CARRY timer_1129_add_4_3 (.CI(n25478), .I0(GND_net), .I1(timer[1]), 
            .CO(n25479));
    SB_LUT4 timer_1129_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n24800), .O(one_wire_N_449[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n25386), .I0(n2295), .I1(n2324), .CO(n25387));
    SB_CARRY timer_1129_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n25478));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n25385), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_7 (.CI(n24800), .I0(timer[5]), .I1(n1[5]), .CO(n24801));
    SB_LUT4 i1_4_lut (.I0(one_wire_N_449[4]), .I1(one_wire_N_449[3]), .I2(n30197), 
            .I3(n26076), .O(n111));
    defparam i1_4_lut.LUT_INIT = 16'h5155;
    SB_LUT4 i1_4_lut_adj_1414 (.I0(n111), .I1(n30197), .I2(one_wire_N_449[2]), 
            .I3(one_wire_N_449[3]), .O(n116));
    defparam i1_4_lut_adj_1414.LUT_INIT = 16'haeee;
    SB_CARRY mod_5_add_1607_16 (.CI(n25385), .I0(n2296), .I1(n2324), .CO(n25386));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n25477), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n25384), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n24799), .O(one_wire_N_449[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n25384), .I0(n2297), .I1(n2324), .CO(n25385));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n25383), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n25476), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n25383), .I0(n2298), .I1(n2324), .CO(n25384));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n25382), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n25476), .I0(n1797), .I1(n1829), .CO(n25477));
    SB_CARRY mod_5_add_1607_13 (.CI(n25382), .I0(n2299), .I1(n2324), .CO(n25383));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n25475), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n25475), .I0(n1798), .I1(n1829), .CO(n25476));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n25381), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n25381), .I0(n2300), .I1(n2324), .CO(n25382));
    SB_CARRY sub_14_add_2_6 (.CI(n24799), .I0(timer[4]), .I1(n1[4]), .CO(n24800));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n25474), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n25380), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n25380), .I0(n2301), .I1(n2324), .CO(n25381));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n25379), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n25379), .I0(n2302), .I1(n2324), .CO(n25380));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n25378), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n25378), .I0(n2303), .I1(n2324), .CO(n25379));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n25377), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n25474), .I0(n1799), .I1(n1829), .CO(n25475));
    SB_CARRY mod_5_add_1607_8 (.CI(n25377), .I0(n2304), .I1(n2324), .CO(n25378));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n25376), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n25376), .I0(n2305), .I1(n2324), .CO(n25377));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n25375), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n25473), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n24798), .O(one_wire_N_449[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n24798), .I0(timer[3]), .I1(n1[3]), .CO(n24799));
    SB_CARRY mod_5_add_1607_6 (.CI(n25375), .I0(n2306), .I1(n2324), .CO(n25376));
    SB_CARRY mod_5_add_1272_12 (.CI(n25473), .I0(n1800), .I1(n1829), .CO(n25474));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n25472), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n25374), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n25374), .I0(n2307), .I1(n2324), .CO(n25375));
    SB_CARRY mod_5_add_1272_11 (.CI(n25472), .I0(n1801), .I1(n1829), .CO(n25473));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n25471), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n25373), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n25471), .I0(n1802), .I1(n1829), .CO(n25472));
    SB_CARRY mod_5_add_1607_4 (.CI(n25373), .I0(n2308), .I1(n2324), .CO(n25374));
    SB_LUT4 i7_4_lut (.I0(one_wire_N_449[10]), .I1(one_wire_N_449[9]), .I2(n116), 
            .I3(\state[1] ), .O(n18_adj_3818));
    defparam i7_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n36861), 
            .I3(n25372), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n25372), .I0(n2309), .I1(n36861), .CO(n25373));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n25470), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_4_lut (.I0(n807), .I1(n14115), .I2(n30829), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_CARRY mod_5_add_1272_9 (.CI(n25470), .I0(n1803), .I1(n1829), .CO(n25471));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n25469), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n36861), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_8 (.CI(n25469), .I0(n1804), .I1(n1829), .CO(n25470));
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n36861), 
            .CO(n25372));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n25468), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n25468), .I0(n1805), .I1(n1829), .CO(n25469));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n25467), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n24797), .O(one_wire_N_449[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30523_3_lut_4_lut (.I0(n14115), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n30829), .O(n30953));   // verilog/neopixel.v(22[26:36])
    defparam i30523_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_CARRY mod_5_add_1272_6 (.CI(n25467), .I0(n1806), .I1(n1829), .CO(n25468));
    SB_CARRY sub_14_add_2_4 (.CI(n24797), .I0(timer[2]), .I1(n1[2]), .CO(n24798));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4), .I1(timer[1]), .I2(n1[1]), .I3(n24796), 
            .O(n26076)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n25466), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n24796), .I0(timer[1]), .I1(n1[1]), .CO(n24797));
    SB_CARRY mod_5_add_1272_5 (.CI(n25466), .I0(n1807), .I1(n1829), .CO(n25467));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_449[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i9_4_lut_adj_1415 (.I0(one_wire_N_449[5]), .I1(n18_adj_3818), 
            .I2(one_wire_N_449[8]), .I3(start), .O(n20_adj_3821));
    defparam i9_4_lut_adj_1415.LUT_INIT = 16'h0004;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n25465), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n24638), 
            .O(n34301)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1272_4 (.CI(n25465), .I0(n1808), .I1(n1829), .CO(n25466));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n36862), 
            .I3(n25464), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n25464), .I0(n1809), .I1(n36862), .CO(n25465));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n36862), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n36862), 
            .CO(n25464));
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n24637), 
            .O(n34295)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i31223_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36860));
    defparam i31223_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_449[11]), .I1(one_wire_N_449[6]), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_21_32 (.CI(n24637), .I0(bit_ctr[30]), .I1(GND_net), .CO(n24638));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n24796));
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_31_lut (.I0(n19), .I1(bit_ctr[29]), .I2(GND_net), .I3(n24636), 
            .O(n34294)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31228_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36865));
    defparam i31228_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_31 (.CI(n24636), .I0(bit_ctr[29]), .I1(GND_net), .CO(n24637));
    SB_LUT4 add_21_30_lut (.I0(n19), .I1(bit_ctr[28]), .I2(GND_net), .I3(n24635), 
            .O(n34293)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_12_lut (.I0(n19), .I1(bit_ctr[10]), .I2(GND_net), .I3(n24617), 
            .O(n34307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_30 (.CI(n24635), .I0(bit_ctr[28]), .I1(GND_net), .CO(n24636));
    SB_LUT4 add_21_29_lut (.I0(n19), .I1(bit_ctr[27]), .I2(GND_net), .I3(n24634), 
            .O(n34292)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n24609), 
            .O(n34302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n25304), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n25303), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_29 (.CI(n24634), .I0(bit_ctr[27]), .I1(GND_net), .CO(n24635));
    SB_CARRY mod_5_add_1674_21 (.CI(n25303), .I0(n2391), .I1(n2423), .CO(n25304));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n25302), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n25302), .I0(n2392), .I1(n2423), .CO(n25303));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n25301), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n25301), .I0(n2393), .I1(n2423), .CO(n25302));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n25300), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n25456), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n25300), .I0(n2394), .I1(n2423), .CO(n25301));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n25299), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n25299), .I0(n2395), .I1(n2423), .CO(n25300));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n25298), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n25298), .I0(n2396), .I1(n2423), .CO(n25299));
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n25455), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n25297), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31227_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36864));
    defparam i31227_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1674_15 (.CI(n25297), .I0(n2397), .I1(n2423), .CO(n25298));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n25296), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n25296), .I0(n2398), .I1(n2423), .CO(n25297));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n25295), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_12 (.CI(n24617), .I0(bit_ctr[10]), .I1(GND_net), .CO(n24618));
    SB_CARRY mod_5_add_1674_13 (.CI(n25295), .I0(n2399), .I1(n2423), .CO(n25296));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n25294), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n25294), .I0(n2400), .I1(n2423), .CO(n25295));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n25293), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_28_lut (.I0(n19), .I1(bit_ctr[26]), .I2(GND_net), .I3(n24633), 
            .O(n34288)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1339_16 (.CI(n25455), .I0(n1896), .I1(n1928), .CO(n25456));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n25454), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n25293), .I0(n2401), .I1(n2423), .CO(n25294));
    SB_CARRY mod_5_add_1339_15 (.CI(n25454), .I0(n1897), .I1(n1928), .CO(n25455));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n25292), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n25292), .I0(n2402), .I1(n2423), .CO(n25293));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n25291), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n25291), .I0(n2403), .I1(n2423), .CO(n25292));
    SB_CARRY add_21_28 (.CI(n24633), .I0(bit_ctr[26]), .I1(GND_net), .CO(n24634));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n25290), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n25453), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1416 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_3822));
    defparam i11_4_lut_adj_1416.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_3823));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_3824));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1417 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_3825));
    defparam i9_4_lut_adj_1417.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1418 (.I0(n19_adj_3823), .I1(n26_adj_3822), .I2(n1905), 
            .I3(n1903), .O(n28_adj_3826));
    defparam i13_4_lut_adj_1418.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1419 (.I0(n1896), .I1(n28_adj_3826), .I2(n24_adj_3825), 
            .I3(n16_adj_3824), .O(n1928));
    defparam i14_4_lut_adj_1419.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_8 (.CI(n25290), .I0(n2404), .I1(n2423), .CO(n25291));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n25289), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n25289), .I0(n2405), .I1(n2423), .CO(n25290));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n25288), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(one_wire_N_449[7]), .I2(n15393), .I3(n20_adj_3821), 
            .O(n37051));
    defparam i4_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_3_lut_adj_1420 (.I0(bit_ctr[11]), .I1(n2405), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_3827));
    defparam i7_3_lut_adj_1420.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1421 (.I0(n2392), .I1(n2390), .I2(n2394), .I3(n2396), 
            .O(n33_adj_3828));
    defparam i13_4_lut_adj_1421.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1422 (.I0(n2399), .I1(n2402), .I2(n2407), .I3(n2406), 
            .O(n32_adj_3829));
    defparam i12_4_lut_adj_1422.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1423 (.I0(n2408), .I1(n2395), .I2(n2391), .I3(n2398), 
            .O(n31_adj_3830));
    defparam i11_4_lut_adj_1423.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1424 (.I0(n2393), .I1(n2397), .I2(n2401), .I3(n2403), 
            .O(n35));
    defparam i15_4_lut_adj_1424.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1425 (.I0(n33_adj_3828), .I1(n27_adj_3827), .I2(n2404), 
            .I3(n2400), .O(n37_adj_3831));
    defparam i17_4_lut_adj_1425.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1426 (.I0(n37_adj_3831), .I1(n35), .I2(n31_adj_3830), 
            .I3(n32_adj_3829), .O(n2423));
    defparam i19_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_6 (.CI(n25288), .I0(n2406), .I1(n2423), .CO(n25289));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n25287), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n25453), .I0(n1898), .I1(n1928), .CO(n25454));
    SB_CARRY mod_5_add_1674_5 (.CI(n25287), .I0(n2407), .I1(n2423), .CO(n25288));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n25286), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n25452), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1427 (.I0(n2205), .I1(n2199), .I2(n2198), .I3(n2203), 
            .O(n28_adj_3832));
    defparam i10_4_lut_adj_1427.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1428 (.I0(n2194), .I1(n2200), .I2(n2192), .I3(n2201), 
            .O(n31_adj_3833));
    defparam i13_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1429 (.I0(n2204), .I1(bit_ctr[13]), .I2(n2209), 
            .I3(GND_net), .O(n22_adj_3834));
    defparam i4_3_lut_adj_1429.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1430 (.I0(n2197), .I1(n2208), .I2(n2207), .I3(n2193), 
            .O(n30_adj_3835));
    defparam i12_4_lut_adj_1430.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1431 (.I0(n31_adj_3833), .I1(n2202), .I2(n28_adj_3832), 
            .I3(n2206), .O(n34_adj_3836));
    defparam i16_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1432 (.I0(n2196), .I1(n2195), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_3837));
    defparam i3_2_lut_adj_1432.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1433 (.I0(n21_adj_3837), .I1(n34_adj_3836), .I2(n30_adj_3835), 
            .I3(n22_adj_3834), .O(n2225));
    defparam i17_4_lut_adj_1433.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1339_13 (.CI(n25452), .I0(n1899), .I1(n1928), .CO(n25453));
    SB_CARRY mod_5_add_1674_4 (.CI(n25286), .I0(n2408), .I1(n2423), .CO(n25287));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n36864), 
            .I3(n25285), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n25285), .I0(n2409), .I1(n36864), .CO(n25286));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n36864), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n36864), 
            .CO(n25285));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n25451), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_27_lut (.I0(n19), .I1(bit_ctr[25]), .I2(GND_net), .I3(n24632), 
            .O(n34323)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_27 (.CI(n24632), .I0(bit_ctr[25]), .I1(GND_net), .CO(n24633));
    SB_LUT4 add_21_26_lut (.I0(n19), .I1(bit_ctr[24]), .I2(GND_net), .I3(n24631), 
            .O(n34322)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_26 (.CI(n24631), .I0(bit_ctr[24]), .I1(GND_net), .CO(n24632));
    SB_LUT4 add_21_25_lut (.I0(n19), .I1(bit_ctr[23]), .I2(GND_net), .I3(n24630), 
            .O(n34320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_11_lut (.I0(n19), .I1(bit_ctr[9]), .I2(GND_net), .I3(n24616), 
            .O(n34296)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1339_12 (.CI(n25451), .I0(n1900), .I1(n1928), .CO(n25452));
    SB_CARRY add_21_25 (.CI(n24630), .I0(bit_ctr[23]), .I1(GND_net), .CO(n24631));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n25450), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n25450), .I0(n1901), .I1(n1928), .CO(n25451));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n25449), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n25449), .I0(n1902), .I1(n1928), .CO(n25450));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n25448), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n25448), .I0(n1903), .I1(n1928), .CO(n25449));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n25447), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n25447), .I0(n1904), .I1(n1928), .CO(n25448));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n25446), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n24616), .I0(bit_ctr[9]), .I1(GND_net), .CO(n24617));
    SB_CARRY mod_5_add_1339_7 (.CI(n25446), .I0(n1905), .I1(n1928), .CO(n25447));
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n24629), 
            .O(n34319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n25445), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n25445), .I0(n1906), .I1(n1928), .CO(n25446));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n25444), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n25444), .I0(n1907), .I1(n1928), .CO(n25445));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n25443), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n25443), .I0(n1908), .I1(n1928), .CO(n25444));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n36865), 
            .I3(n25442), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n25437), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_24 (.CI(n24629), .I0(bit_ctr[22]), .I1(GND_net), .CO(n24630));
    SB_LUT4 add_21_10_lut (.I0(n19), .I1(bit_ctr[8]), .I2(GND_net), .I3(n24615), 
            .O(n34291)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_10 (.CI(n24615), .I0(bit_ctr[8]), .I1(GND_net), .CO(n24616));
    SB_DFF timer_1129__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1339_3 (.CI(n25442), .I0(n1909), .I1(n36865), .CO(n25443));
    SB_LUT4 add_21_23_lut (.I0(n19), .I1(bit_ctr[21]), .I2(GND_net), .I3(n24628), 
            .O(n34318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_23 (.CI(n24628), .I0(bit_ctr[21]), .I1(GND_net), .CO(n24629));
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n24614), 
            .O(n34290)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i31222_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36859));
    defparam i31222_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_4 (.CI(n24609), .I0(bit_ctr[2]), .I1(GND_net), .CO(n24610));
    SB_CARRY add_21_9 (.CI(n24614), .I0(bit_ctr[7]), .I1(GND_net), .CO(n24615));
    SB_LUT4 add_21_22_lut (.I0(n19), .I1(bit_ctr[20]), .I2(GND_net), .I3(n24627), 
            .O(n34317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3838));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'heeee;
    SB_LUT4 i17469_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n21839));
    defparam i17469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1435 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_3838), 
            .O(n30_adj_3839));
    defparam i13_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1436 (.I0(n2098), .I1(n21839), .I2(n2094), .I3(n2099), 
            .O(n28_adj_3840));
    defparam i11_4_lut_adj_1436.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1437 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_3841));
    defparam i12_4_lut_adj_1437.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1438 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_3842));
    defparam i10_4_lut_adj_1438.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1439 (.I0(n27_adj_3842), .I1(n29_adj_3841), .I2(n28_adj_3840), 
            .I3(n30_adj_3839), .O(n2126));
    defparam i16_4_lut_adj_1439.LUT_INIT = 16'hfffe;
    SB_LUT4 i31220_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36857));
    defparam i31220_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_449[3]), .I1(one_wire_N_449[4]), .I2(one_wire_N_449[2]), 
            .I3(GND_net), .O(n25921));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut (.I0(n26076), .I1(one_wire_N_449[4]), .I2(one_wire_N_449[3]), 
            .I3(GND_net), .O(n30886));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 equal_322_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n15386));
    defparam equal_322_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut_adj_1440 (.I0(one_wire_N_449[10]), .I1(one_wire_N_449[8]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/neopixel.v(104[14:39])
    defparam i2_2_lut_adj_1440.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_449[5]), .I1(one_wire_N_449[11]), .I2(one_wire_N_449[7]), 
            .I3(n15393), .O(n14_adj_3843));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1441 (.I0(one_wire_N_449[9]), .I1(n14_adj_3843), 
            .I2(n10), .I3(one_wire_N_449[6]), .O(n15289));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1441.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1442 (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_3844));
    defparam i2_2_lut_adj_1442.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1443 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut_adj_1443.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1444 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut_adj_1444.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1445 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut_adj_1445.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1446 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut_adj_1446.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1447 (.I0(bit_ctr[3]), .I1(n30_adj_3844), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut_adj_1447.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_298[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2017_3_lut (.I0(n15387), .I1(\state_3__N_298[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4377));
    defparam i2017_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n919), .I2(n4377), .I3(\state[0] ), 
            .O(n4404));
    defparam i2_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 mux_645_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_506 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_645_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(\color[18] ), .I2(\color[19] ), 
            .I3(bit_ctr[1]), .O(n36990));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 add_21_3_lut (.I0(n19), .I1(bit_ctr[1]), .I2(GND_net), .I3(n24608), 
            .O(n34321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n36990_bdd_4_lut (.I0(n36990), .I1(\color[17] ), .I2(\color[16] ), 
            .I3(bit_ctr[1]), .O(n36993));
    defparam n36990_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_21_22 (.CI(n24627), .I0(bit_ctr[20]), .I1(GND_net), .CO(n24628));
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n24613), 
            .O(n34289)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n25179), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n25178), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n25178), .I0(n2490), .I1(n2522), .CO(n25179));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n25177), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n25177), .I0(n2491), .I1(n2522), .CO(n25178));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n25176), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n25176), .I0(n2492), .I1(n2522), .CO(n25177));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n25175), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n25175), .I0(n2493), .I1(n2522), .CO(n25176));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n25174), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n25174), .I0(n2494), .I1(n2522), .CO(n25175));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n25173), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n25173), .I0(n2495), .I1(n2522), .CO(n25174));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n25172), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n25172), .I0(n2496), .I1(n2522), .CO(n25173));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n25171), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n25171), .I0(n2497), .I1(n2522), .CO(n25172));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n25170), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n25170), .I0(n2498), .I1(n2522), .CO(n25171));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n25169), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n25169), .I0(n2499), .I1(n2522), .CO(n25170));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n25168), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n25168), .I0(n2500), .I1(n2522), .CO(n25169));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n25167), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n25167), .I0(n2501), .I1(n2522), .CO(n25168));
    SB_LUT4 add_21_21_lut (.I0(n19), .I1(bit_ctr[19]), .I2(GND_net), .I3(n24626), 
            .O(n34316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n25166), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n25166), .I0(n2502), .I1(n2522), .CO(n25167));
    SB_CARRY add_21_21 (.CI(n24626), .I0(bit_ctr[19]), .I1(GND_net), .CO(n24627));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n25165), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n24608), .I0(bit_ctr[1]), .I1(GND_net), .CO(n24609));
    SB_CARRY mod_5_add_1741_9 (.CI(n25165), .I0(n2503), .I1(n2522), .CO(n25166));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n25164), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n25164), .I0(n2504), .I1(n2522), .CO(n25165));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n25163), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n25163), .I0(n2505), .I1(n2522), .CO(n25164));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n25162), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n25162), .I0(n2506), .I1(n2522), .CO(n25163));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n25161), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n24613), .I0(bit_ctr[6]), .I1(GND_net), .CO(n24614));
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n34305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_5 (.CI(n25161), .I0(n2507), .I1(n2522), .CO(n25162));
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n24612), 
            .O(n34306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n25160), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n25160), .I0(n2508), .I1(n2522), .CO(n25161));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n36866), 
            .I3(n25159), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n24625), 
            .O(n34315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_3 (.CI(n25159), .I0(n2509), .I1(n36866), .CO(n25160));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n36866), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n36866), 
            .CO(n25159));
    SB_CARRY add_21_20 (.CI(n24625), .I0(bit_ctr[18]), .I1(GND_net), .CO(n24626));
    SB_LUT4 add_21_19_lut (.I0(n19), .I1(bit_ctr[17]), .I2(GND_net), .I3(n24624), 
            .O(n34314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_7 (.CI(n24612), .I0(bit_ctr[5]), .I1(GND_net), .CO(n24613));
    SB_CARRY add_21_19 (.CI(n24624), .I0(bit_ctr[17]), .I1(GND_net), .CO(n24625));
    SB_LUT4 add_21_18_lut (.I0(n19), .I1(bit_ctr[16]), .I2(GND_net), .I3(n24623), 
            .O(n34313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n24611), 
            .O(n34304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_18 (.CI(n24623), .I0(bit_ctr[16]), .I1(GND_net), .CO(n24624));
    SB_LUT4 add_21_17_lut (.I0(n19), .I1(bit_ctr[15]), .I2(GND_net), .I3(n24622), 
            .O(n34312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_17 (.CI(n24622), .I0(bit_ctr[15]), .I1(GND_net), .CO(n24623));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_449[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n24826), .O(n22_adj_3816)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_449[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n24825), .O(n23_adj_3815)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n24825), .I0(timer[30]), .I1(n1[30]), 
            .CO(n24826));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n16527), .D(state_3__N_298[0]), 
            .S(n30957));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n24621), 
            .O(n34311)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n24608));
    SB_LUT4 sub_14_add_2_31_lut (.I0(GND_net), .I1(timer[29]), .I2(n1[29]), 
            .I3(n24824), .O(one_wire_N_449[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n24611), .I0(bit_ctr[4]), .I1(GND_net), .CO(n24612));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n25119), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n25118), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n25118), .I0(n2589), .I1(n2621), .CO(n25119));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n25117), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n25117), .I0(n2590), .I1(n2621), .CO(n25118));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n25116), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n25116), .I0(n2591), .I1(n2621), .CO(n25117));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n25115), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n25115), .I0(n2592), .I1(n2621), .CO(n25116));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n25114), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n25114), .I0(n2593), .I1(n2621), .CO(n25115));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n25113), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n25113), .I0(n2594), .I1(n2621), .CO(n25114));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n25112), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n25112), .I0(n2595), .I1(n2621), .CO(n25113));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n25111), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n25111), .I0(n2596), .I1(n2621), .CO(n25112));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n25110), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n25110), .I0(n2597), .I1(n2621), .CO(n25111));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n25109), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n25109), .I0(n2598), .I1(n2621), .CO(n25110));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n25108), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n25108), .I0(n2599), .I1(n2621), .CO(n25109));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n25107), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n25107), .I0(n2600), .I1(n2621), .CO(n25108));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n25106), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n25106), .I0(n2601), .I1(n2621), .CO(n25107));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n25105), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n25105), .I0(n2602), .I1(n2621), .CO(n25106));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n25104), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n25104), .I0(n2603), .I1(n2621), .CO(n25105));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n25103), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n25103), .I0(n2604), .I1(n2621), .CO(n25104));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n25102), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n25102), .I0(n2605), .I1(n2621), .CO(n25103));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n25101), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n25101), .I0(n2606), .I1(n2621), .CO(n25102));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n25100), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n25100), .I0(n2607), .I1(n2621), .CO(n25101));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n25099), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n25099), .I0(n2608), .I1(n2621), .CO(n25100));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n36867), 
            .I3(n25098), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n25098), .I0(n2609), .I1(n36867), .CO(n25099));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n36867), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n36867), 
            .CO(n25098));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n25067), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n25066), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n25066), .I0(n2688), .I1(n2720), .CO(n25067));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n25065), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n25065), .I0(n2689), .I1(n2720), .CO(n25066));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n25064), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n25064), .I0(n2690), .I1(n2720), .CO(n25065));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n25063), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n25063), .I0(n2691), .I1(n2720), .CO(n25064));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n25062), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n25062), .I0(n2692), .I1(n2720), .CO(n25063));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n25061), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n25061), .I0(n2693), .I1(n2720), .CO(n25062));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n25060), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n25060), .I0(n2694), .I1(n2720), .CO(n25061));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n25059), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n25059), .I0(n2695), .I1(n2720), .CO(n25060));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n25058), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n25058), .I0(n2696), .I1(n2720), .CO(n25059));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n25057), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n25057), .I0(n2697), .I1(n2720), .CO(n25058));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n25056), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n25056), .I0(n2698), .I1(n2720), .CO(n25057));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n25055), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n25055), .I0(n2699), .I1(n2720), .CO(n25056));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n25054), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n25054), .I0(n2700), .I1(n2720), .CO(n25055));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n25053), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n25053), .I0(n2701), .I1(n2720), .CO(n25054));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n25052), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n25052), .I0(n2702), .I1(n2720), .CO(n25053));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n25051), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n25051), .I0(n2703), .I1(n2720), .CO(n25052));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n25050), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n25050), .I0(n2704), .I1(n2720), .CO(n25051));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n25049), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n25049), .I0(n2705), .I1(n2720), .CO(n25050));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n25048), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n25048), .I0(n2706), .I1(n2720), .CO(n25049));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n25047), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n25047), .I0(n2707), .I1(n2720), .CO(n25048));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n25046), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n25046), .I0(n2708), .I1(n2720), .CO(n25047));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n36868), 
            .I3(n25045), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n25045), .I0(n2709), .I1(n36868), .CO(n25046));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n36868), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n36868), 
            .CO(n25045));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n25029), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n25028), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n25028), .I0(n2787), .I1(n2819), .CO(n25029));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n25027), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n25027), .I0(n2788), .I1(n2819), .CO(n25028));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n25026), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n25026), .I0(n2789), .I1(n2819), .CO(n25027));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n25025), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n25025), .I0(n2790), .I1(n2819), .CO(n25026));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n25024), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n25024), .I0(n2791), .I1(n2819), .CO(n25025));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n25023), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n25023), .I0(n2792), .I1(n2819), .CO(n25024));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n25022), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n25022), .I0(n2793), .I1(n2819), .CO(n25023));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n25021), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n25021), .I0(n2794), .I1(n2819), .CO(n25022));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n25020), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n25020), .I0(n2795), .I1(n2819), .CO(n25021));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n25019), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n25019), .I0(n2796), .I1(n2819), .CO(n25020));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n25018), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n25018), .I0(n2797), .I1(n2819), .CO(n25019));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n25017), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n25017), .I0(n2798), .I1(n2819), .CO(n25018));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n25016), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n25016), .I0(n2799), .I1(n2819), .CO(n25017));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n25015), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n25015), .I0(n2800), .I1(n2819), .CO(n25016));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n25014), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n25014), .I0(n2801), .I1(n2819), .CO(n25015));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n25013), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n25013), .I0(n2802), .I1(n2819), .CO(n25014));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n25012), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n25012), .I0(n2803), .I1(n2819), .CO(n25013));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n25011), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n25011), .I0(n2804), .I1(n2819), .CO(n25012));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n25010), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n25010), .I0(n2805), .I1(n2819), .CO(n25011));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n25009), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n25009), .I0(n2806), .I1(n2819), .CO(n25010));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n25008), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n25008), .I0(n2807), .I1(n2819), .CO(n25009));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n25007), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n25007), .I0(n2808), .I1(n2819), .CO(n25008));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n36869), 
            .I3(n25006), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n25006), .I0(n2809), .I1(n36869), .CO(n25007));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n36869), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n36869), 
            .CO(n25006));
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n31011), .D(\neo_pixel_transmitter.done_N_512 ), 
            .R(n32288));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_31 (.CI(n24824), .I0(timer[29]), .I1(n1[29]), 
            .CO(n24825));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n24994), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n24993), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n24993), .I0(n2886), .I1(n2918), .CO(n24994));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n24992), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n24992), .I0(n2887), .I1(n2918), .CO(n24993));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n24991), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n24991), .I0(n2888), .I1(n2918), .CO(n24992));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n24990), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n24990), .I0(n2889), .I1(n2918), .CO(n24991));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n24989), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n24989), .I0(n2890), .I1(n2918), .CO(n24990));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n24988), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n24988), .I0(n2891), .I1(n2918), .CO(n24989));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n24987), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n24987), .I0(n2892), .I1(n2918), .CO(n24988));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n24986), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n24986), .I0(n2893), .I1(n2918), .CO(n24987));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n24985), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n24985), .I0(n2894), .I1(n2918), .CO(n24986));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n24984), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_449[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n24823), .O(n26_adj_3817)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_17 (.CI(n24984), .I0(n2895), .I1(n2918), .CO(n24985));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n24983), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n24983), .I0(n2896), .I1(n2918), .CO(n24984));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n24982), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n24982), .I0(n2897), .I1(n2918), .CO(n24983));
    SB_CARRY sub_14_add_2_30 (.CI(n24823), .I0(timer[28]), .I1(n1[28]), 
            .CO(n24824));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n24981), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_14 (.CI(n24981), .I0(n2898), .I1(n2918), .CO(n24982));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n24980), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n24980), .I0(n2899), .I1(n2918), .CO(n24981));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n24979), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n24979), .I0(n2900), .I1(n2918), .CO(n24980));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n24978), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n24978), .I0(n2901), .I1(n2918), .CO(n24979));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n24977), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n24977), .I0(n2902), .I1(n2918), .CO(n24978));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n24976), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n24976), .I0(n2903), .I1(n2918), .CO(n24977));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n24975), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n24975), .I0(n2904), .I1(n2918), .CO(n24976));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n24974), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n24974), .I0(n2905), .I1(n2918), .CO(n24975));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n24973), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n24973), .I0(n2906), .I1(n2918), .CO(n24974));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n24972), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n25645), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n25644), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n25644), .I0(n906), .I1(VCC_net), .CO(n25645));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n30953), .I2(VCC_net), 
            .I3(n25643), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n25643), .I0(n30953), .I1(VCC_net), 
            .CO(n25644));
    SB_CARRY mod_5_add_2009_5 (.CI(n24972), .I0(n2907), .I1(n2918), .CO(n24973));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n16628), .I2(VCC_net), 
            .I3(n25642), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n24971), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_4 (.CI(n25642), .I0(n16628), .I1(VCC_net), 
            .CO(n25643));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14113), .I2(GND_net), 
            .I3(n25641), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n25641), .I0(n14113), .I1(GND_net), 
            .CO(n25642));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n25641));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_3846), .I1(n4_adj_3846), .I2(n1037), 
            .I3(n25640), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n25639), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n25639), .I0(n1005), .I1(n1037), .CO(n25640));
    SB_CARRY mod_5_add_2009_4 (.CI(n24971), .I0(n2908), .I1(n2918), .CO(n24972));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n36870), 
            .I3(n24970), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n24970), .I0(n2909), .I1(n36870), .CO(n24971));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n25638), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n36870), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_6 (.CI(n25638), .I0(n1006), .I1(n1037), .CO(n25639));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n36870), 
            .CO(n24970));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n25637), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n24969), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n25637), .I0(n1007), .I1(n1037), .CO(n25638));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n25636), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n24621), .I0(bit_ctr[14]), .I1(GND_net), .CO(n24622));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n24968), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n36865), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_27 (.CI(n24968), .I0(n2985), .I1(n3017), .CO(n24969));
    SB_CARRY mod_5_add_736_4 (.CI(n25636), .I0(n1008), .I1(n1037), .CO(n25637));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n36871), 
            .I3(n25635), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n36865), 
            .CO(n25442));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n24967), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n25441), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n24967), .I0(n2986), .I1(n3017), .CO(n24968));
    SB_CARRY mod_5_add_736_3 (.CI(n25635), .I0(n1009), .I1(n36871), .CO(n25636));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n36871), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n24966), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n36871), 
            .CO(n25635));
    SB_LUT4 sub_14_add_2_29_lut (.I0(GND_net), .I1(timer[27]), .I2(n1[27]), 
            .I3(n24822), .O(one_wire_N_449[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n25634), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n25633), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n25633), .I0(n1104), .I1(n1136), .CO(n25634));
    SB_CARRY mod_5_add_2076_25 (.CI(n24966), .I0(n2987), .I1(n3017), .CO(n24967));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n25632), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n25632), .I0(n1105), .I1(n1136), .CO(n25633));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n24965), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n25631), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n25631), .I0(n1106), .I1(n1136), .CO(n25632));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n25630), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n25630), .I0(n1107), .I1(n1136), .CO(n25631));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n25629), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n25629), .I0(n1108), .I1(n1136), .CO(n25630));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n36873), 
            .I3(n25628), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n25628), .I0(n1109), .I1(n36873), .CO(n25629));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n36873), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_24 (.CI(n24965), .I0(n2988), .I1(n3017), .CO(n24966));
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n36873), 
            .CO(n25628));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n25627), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n25626), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n25626), .I0(n1203), .I1(n1235), .CO(n25627));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n25625), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n25625), .I0(n1204), .I1(n1235), .CO(n25626));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n25624), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n25624), .I0(n1205), .I1(n1235), .CO(n25625));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n25623), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n25623), .I0(n1206), .I1(n1235), .CO(n25624));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n25622), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n25622), .I0(n1207), .I1(n1235), .CO(n25623));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n25621), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n24964), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n25621), .I0(n1208), .I1(n1235), .CO(n25622));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n25440), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n36874), 
            .I3(n25620), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_17 (.CI(n25440), .I0(n1995), .I1(n2027), .CO(n25441));
    SB_CARRY mod_5_add_870_3 (.CI(n25620), .I0(n1209), .I1(n36874), .CO(n25621));
    SB_CARRY mod_5_add_2076_23 (.CI(n24964), .I0(n2989), .I1(n3017), .CO(n24965));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n24963), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n36874), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_22 (.CI(n24963), .I0(n2990), .I1(n3017), .CO(n24964));
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n36874), 
            .CO(n25620));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n25619), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n24962), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n25618), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n24962), .I0(n2991), .I1(n3017), .CO(n24963));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n24961), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n24961), .I0(n2992), .I1(n3017), .CO(n24962));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n24960), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_29 (.CI(n24822), .I0(timer[27]), .I1(n1[27]), 
            .CO(n24823));
    SB_CARRY mod_5_add_2076_19 (.CI(n24960), .I0(n2993), .I1(n3017), .CO(n24961));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n24959), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n25439), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n24821), .O(one_wire_N_449[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n25618), .I0(n1302), .I1(n1334), .CO(n25619));
    SB_CARRY mod_5_add_2076_18 (.CI(n24959), .I0(n2994), .I1(n3017), .CO(n24960));
    SB_CARRY mod_5_add_1406_16 (.CI(n25439), .I0(n1996), .I1(n2027), .CO(n25440));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n25617), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n25617), .I0(n1303), .I1(n1334), .CO(n25618));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n25616), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n24958), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_28 (.CI(n24821), .I0(timer[26]), .I1(n1[26]), 
            .CO(n24822));
    SB_CARRY mod_5_add_2076_17 (.CI(n24958), .I0(n2995), .I1(n3017), .CO(n24959));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n25438), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n25616), .I0(n1304), .I1(n1334), .CO(n25617));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n24957), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n25438), .I0(n1997), .I1(n2027), .CO(n25439));
    SB_CARRY mod_5_add_2076_16 (.CI(n24957), .I0(n2996), .I1(n3017), .CO(n24958));
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n29087));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n24956), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n24820), .O(one_wire_N_449[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n25436), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n24956), .I0(n2997), .I1(n3017), .CO(n24957));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n24955), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n24955), .I0(n2998), .I1(n3017), .CO(n24956));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n24954), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n24954), .I0(n2999), .I1(n3017), .CO(n24955));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n24953), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n25615), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n24953), .I0(n3000), .I1(n3017), .CO(n24954));
    SB_CARRY mod_5_add_937_7 (.CI(n25615), .I0(n1305), .I1(n1334), .CO(n25616));
    SB_DFF timer_1129__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n24952), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n25614), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n24952), .I0(n3001), .I1(n3017), .CO(n24953));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n24951), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n24951), .I0(n3002), .I1(n3017), .CO(n24952));
    SB_CARRY mod_5_add_937_6 (.CI(n25614), .I0(n1306), .I1(n1334), .CO(n25615));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n25613), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n25613), .I0(n1307), .I1(n1334), .CO(n25614));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n25612), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n25612), .I0(n1308), .I1(n1334), .CO(n25613));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n36875), 
            .I3(n25611), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n24950), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_3 (.CI(n25611), .I0(n1309), .I1(n36875), .CO(n25612));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n36875), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_9 (.CI(n24950), .I0(n3003), .I1(n3017), .CO(n24951));
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n36875), 
            .CO(n25611));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n25610), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n25609), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n25609), .I0(n1401), .I1(n1433), .CO(n25610));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n25608), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n25608), .I0(n1402), .I1(n1433), .CO(n25609));
    SB_DFF timer_1129__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1129__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n25607), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n16771));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n29081));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n24949), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n24949), .I0(n3004), .I1(n3017), .CO(n24950));
    SB_CARRY mod_5_add_1004_9 (.CI(n25607), .I0(n1403), .I1(n1433), .CO(n25608));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n25606), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n24948), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17004));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_8 (.CI(n25606), .I0(n1404), .I1(n1433), .CO(n25607));
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17003));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n25605), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17002));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_7 (.CI(n25605), .I0(n1405), .I1(n1433), .CO(n25606));
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17001));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n25604), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17000));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_6 (.CI(n25604), .I0(n1406), .I1(n1433), .CO(n25605));
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n16999));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n25603), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n16998));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_5 (.CI(n25603), .I0(n1407), .I1(n1433), .CO(n25604));
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n16997));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n25602), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n16996));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_4 (.CI(n25602), .I0(n1408), .I1(n1433), .CO(n25603));
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n16995));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n36876), 
            .I3(n25601), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n16994));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_3 (.CI(n25601), .I0(n1409), .I1(n36876), .CO(n25602));
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n16993));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n36876), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n16992));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n36876), 
            .CO(n25601));
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n16991));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n25600), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n16990));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_7 (.CI(n24948), .I0(n3005), .I1(n3017), .CO(n24949));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n25599), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n16989));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n24947), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n25599), .I0(n1500), .I1(n1532), .CO(n25600));
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n16988));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n25598), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n16987));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_11 (.CI(n25598), .I0(n1501), .I1(n1532), .CO(n25599));
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n16986));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n25597), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n16985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_10 (.CI(n25597), .I0(n1502), .I1(n1532), .CO(n25598));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n25596), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n16983));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_9 (.CI(n25596), .I0(n1503), .I1(n1532), .CO(n25597));
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n16982));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n25595), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n16981));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_8 (.CI(n25595), .I0(n1504), .I1(n1532), .CO(n25596));
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n16980));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n25594), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n16979));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_7 (.CI(n25594), .I0(n1505), .I1(n1532), .CO(n25595));
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n16978));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n25593), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n16977));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_6 (.CI(n25593), .I0(n1506), .I1(n1532), .CO(n25594));
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n16976));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n25592), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n16975));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_5 (.CI(n25592), .I0(n1507), .I1(n1532), .CO(n25593));
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n16974));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n25591), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n25591), .I0(n1508), .I1(n1532), .CO(n25592));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n36877), 
            .I3(n25590), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n25590), .I0(n1509), .I1(n36877), .CO(n25591));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n36877), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n36877), 
            .CO(n25590));
    SB_CARRY mod_5_add_2076_6 (.CI(n24947), .I0(n3006), .I1(n3017), .CO(n24948));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n24946), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n24946), .I0(n3007), .I1(n3017), .CO(n24947));
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n29079));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n24945), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n24945), .I0(n3008), .I1(n3017), .CO(n24946));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n36872), 
            .I3(n24944), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n24944), .I0(n3009), .I1(n36872), .CO(n24945));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n36872), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n16923));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n24620), 
            .O(n34310)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n36872), 
            .CO(n24944));
    SB_CARRY sub_14_add_2_27 (.CI(n24820), .I0(timer[25]), .I1(n1[25]), 
            .CO(n24821));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n24943), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n24942), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n24942), .I0(n3084), .I1(n3116), .CO(n24943));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n24941), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n24941), .I0(n3085), .I1(n3116), .CO(n24942));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n24940), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n24940), .I0(n3086), .I1(n3116), .CO(n24941));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n24939), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n24939), .I0(n3087), .I1(n3116), .CO(n24940));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n24819), .O(one_wire_N_449[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n24938), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n24938), .I0(n3088), .I1(n3116), .CO(n24939));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n24937), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_26 (.CI(n24819), .I0(timer[24]), .I1(n1[24]), 
            .CO(n24820));
    SB_CARRY mod_5_add_2143_23 (.CI(n24937), .I0(n3089), .I1(n3116), .CO(n24938));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n24936), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n24936), .I0(n3090), .I1(n3116), .CO(n24937));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n25543), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n24935), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n25542), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n24935), .I0(n3091), .I1(n3116), .CO(n24936));
    SB_CARRY mod_5_add_1138_13 (.CI(n25542), .I0(n1599), .I1(n1631), .CO(n25543));
    SB_LUT4 sub_14_add_2_25_lut (.I0(GND_net), .I1(timer[23]), .I2(n1[23]), 
            .I3(n24818), .O(one_wire_N_449[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n25541), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n24934), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n25541), .I0(n1600), .I1(n1631), .CO(n25542));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n25540), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n24934), .I0(n3092), .I1(n3116), .CO(n24935));
    SB_CARRY mod_5_add_1138_11 (.CI(n25540), .I0(n1601), .I1(n1631), .CO(n25541));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n24933), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n25539), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n25539), .I0(n1602), .I1(n1631), .CO(n25540));
    SB_CARRY mod_5_add_2143_19 (.CI(n24933), .I0(n3093), .I1(n3116), .CO(n24934));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n25538), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n24932), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n25538), .I0(n1603), .I1(n1631), .CO(n25539));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n25537), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n24932), .I0(n3094), .I1(n3116), .CO(n24933));
    SB_CARRY mod_5_add_1138_8 (.CI(n25537), .I0(n1604), .I1(n1631), .CO(n25538));
    SB_CARRY sub_14_add_2_25 (.CI(n24818), .I0(timer[23]), .I1(n1[23]), 
            .CO(n24819));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n25536), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n25536), .I0(n1605), .I1(n1631), .CO(n25537));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n25535), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n25535), .I0(n1606), .I1(n1631), .CO(n25536));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n25534), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n25534), .I0(n1607), .I1(n1631), .CO(n25535));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n24931), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n25533), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n25533), .I0(n1608), .I1(n1631), .CO(n25534));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n36879), 
            .I3(n25532), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n25532), .I0(n1609), .I1(n36879), .CO(n25533));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n36879), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n36879), 
            .CO(n25532));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n25531), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n25530), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n25530), .I0(n1698), .I1(n1730), .CO(n25531));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n25529), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n25529), .I0(n1699), .I1(n1730), .CO(n25530));
    SB_CARRY mod_5_add_1406_14 (.CI(n25437), .I0(n1998), .I1(n2027), .CO(n25438));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n25528), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n25528), .I0(n1700), .I1(n1730), .CO(n25529));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n25527), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n25527), .I0(n1701), .I1(n1730), .CO(n25528));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n25526), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n24931), .I0(n3095), .I1(n3116), .CO(n24932));
    SB_CARRY mod_5_add_1205_10 (.CI(n25526), .I0(n1702), .I1(n1730), .CO(n25527));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n24930), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n25525), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n25525), .I0(n1703), .I1(n1730), .CO(n25526));
    SB_CARRY mod_5_add_2143_16 (.CI(n24930), .I0(n3096), .I1(n3116), .CO(n24931));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n25524), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n25524), .I0(n1704), .I1(n1730), .CO(n25525));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n25523), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n24929), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n25523), .I0(n1705), .I1(n1730), .CO(n25524));
    SB_CARRY mod_5_add_2143_15 (.CI(n24929), .I0(n3097), .I1(n3116), .CO(n24930));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n24928), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n25522), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n25522), .I0(n1706), .I1(n1730), .CO(n25523));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n25521), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n25521), .I0(n1707), .I1(n1730), .CO(n25522));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n25520), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n24928), .I0(n3098), .I1(n3116), .CO(n24929));
    SB_CARRY mod_5_add_1205_4 (.CI(n25520), .I0(n1708), .I1(n1730), .CO(n25521));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n24927), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n24927), .I0(n3099), .I1(n3116), .CO(n24928));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n36880), 
            .I3(n25519), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n25519), .I0(n1709), .I1(n36880), .CO(n25520));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n24926), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n24926), .I0(n3100), .I1(n3116), .CO(n24927));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n24925), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n24925), .I0(n3101), .I1(n3116), .CO(n24926));
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n24817), .O(one_wire_N_449[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n24924), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n24924), .I0(n3102), .I1(n3116), .CO(n24925));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n36880), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n36880), 
            .CO(n25519));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n24923), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n24923), .I0(n3103), .I1(n3116), .CO(n24924));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n24922), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n24922), .I0(n3104), .I1(n3116), .CO(n24923));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n24921), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n24921), .I0(n3105), .I1(n3116), .CO(n24922));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n24920), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n24920), .I0(n3106), .I1(n3116), .CO(n24921));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n24919), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n29077));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2143_5 (.CI(n24919), .I0(n3107), .I1(n3116), .CO(n24920));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n24918), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_24 (.CI(n24817), .I0(timer[22]), .I1(n1[22]), 
            .CO(n24818));
    SB_CARRY mod_5_add_2143_4 (.CI(n24918), .I0(n3108), .I1(n3116), .CO(n24919));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n36878), 
            .I3(n24917), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n24917), .I0(n3109), .I1(n36878), .CO(n24918));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n36878), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1129_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n25508), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1129_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n25507), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_32 (.CI(n25507), .I0(GND_net), .I1(timer[30]), 
            .CO(n25508));
    SB_LUT4 timer_1129_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n25506), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_31 (.CI(n25506), .I0(GND_net), .I1(timer[29]), 
            .CO(n25507));
    SB_LUT4 timer_1129_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n25505), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_30 (.CI(n25505), .I0(GND_net), .I1(timer[28]), 
            .CO(n25506));
    SB_LUT4 timer_1129_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n25504), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_29 (.CI(n25504), .I0(GND_net), .I1(timer[27]), 
            .CO(n25505));
    SB_LUT4 timer_1129_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n25503), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n36878), 
            .CO(n24917));
    SB_CARRY timer_1129_add_4_28 (.CI(n25503), .I0(GND_net), .I1(timer[26]), 
            .CO(n25504));
    SB_LUT4 sub_14_add_2_23_lut (.I0(GND_net), .I1(timer[21]), .I2(n1[21]), 
            .I3(n24816), .O(one_wire_N_449[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1129_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n25502), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_27 (.CI(n25502), .I0(GND_net), .I1(timer[25]), 
            .CO(n25503));
    SB_LUT4 timer_1129_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n25501), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_26 (.CI(n25501), .I0(GND_net), .I1(timer[24]), 
            .CO(n25502));
    SB_LUT4 timer_1129_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n25500), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_25 (.CI(n25500), .I0(GND_net), .I1(timer[23]), 
            .CO(n25501));
    SB_CARRY sub_14_add_2_23 (.CI(n24816), .I0(timer[21]), .I1(n1[21]), 
            .CO(n24817));
    SB_CARRY add_21_15 (.CI(n24620), .I0(bit_ctr[13]), .I1(GND_net), .CO(n24621));
    SB_LUT4 timer_1129_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n25499), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_24 (.CI(n25499), .I0(GND_net), .I1(timer[22]), 
            .CO(n25500));
    SB_LUT4 sub_14_add_2_22_lut (.I0(GND_net), .I1(timer[20]), .I2(n1[20]), 
            .I3(n24815), .O(one_wire_N_449[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1129_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n25498), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_23 (.CI(n25498), .I0(GND_net), .I1(timer[21]), 
            .CO(n25499));
    SB_LUT4 timer_1129_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n25497), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_22 (.CI(n25497), .I0(GND_net), .I1(timer[20]), 
            .CO(n25498));
    SB_LUT4 timer_1129_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n25496), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_21 (.CI(n25496), .I0(GND_net), .I1(timer[19]), 
            .CO(n25497));
    SB_LUT4 timer_1129_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n25495), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_20 (.CI(n25495), .I0(GND_net), .I1(timer[18]), 
            .CO(n25496));
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n24619), 
            .O(n34309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1129_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n25494), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1129_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1129_add_4_19 (.CI(n25494), .I0(GND_net), .I1(timer[17]), 
            .CO(n25495));
    SB_CARRY add_21_14 (.CI(n24619), .I0(bit_ctr[12]), .I1(GND_net), .CO(n24620));
    SB_LUT4 i2_2_lut_adj_1448 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3849));
    defparam i2_2_lut_adj_1448.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1449 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_3850));
    defparam i12_4_lut_adj_1449.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1450 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_3851));
    defparam i10_4_lut_adj_1450.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31241_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36878));
    defparam i31241_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31243_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36880));
    defparam i31243_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1451 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_3852));
    defparam i4_3_lut_adj_1451.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1452 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_3853));
    defparam i8_4_lut_adj_1452.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1453 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_3854));
    defparam i7_3_lut_adj_1453.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1454 (.I0(n21_adj_3853), .I1(n17_adj_3852), .I2(n1702), 
            .I3(n1697), .O(n24_adj_3855));
    defparam i11_4_lut_adj_1454.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1455 (.I0(n1700), .I1(n24_adj_3855), .I2(n20_adj_3854), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1455.LUT_INIT = 16'hfffe;
    SB_LUT4 i31242_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36879));
    defparam i31242_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1456 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_3856));
    defparam i11_4_lut_adj_1456.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1457 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_3857));
    defparam i8_4_lut_adj_1457.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1458 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_3858));
    defparam i1_3_lut_adj_1458.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3859));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1459 (.I0(n13_adj_3858), .I1(n20_adj_3857), .I2(n1605), 
            .I3(n1599), .O(n22_adj_3860));
    defparam i10_4_lut_adj_1459.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1460 (.I0(n1601), .I1(n22_adj_3860), .I2(n18_adj_3859), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1460.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_2_lut (.I0(n3106), .I1(n3103), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_3861));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1461 (.I0(n3085), .I1(n3094), .I2(n3093), .I3(n3108), 
            .O(n46_adj_3862));
    defparam i19_4_lut_adj_1461.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1462 (.I0(n3098), .I1(n3090), .I2(n3087), .I3(n3092), 
            .O(n42));
    defparam i15_4_lut_adj_1462.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1463 (.I0(n3099), .I1(n3100), .I2(n3107), .I3(n3095), 
            .O(n44_adj_3863));
    defparam i17_4_lut_adj_1463.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1464 (.I0(n3102), .I1(bit_ctr[4]), .I2(n3109), 
            .I3(GND_net), .O(n31_adj_3864));
    defparam i4_3_lut_adj_1464.LUT_INIT = 16'heaea;
    SB_LUT4 i23_4_lut (.I0(n3091), .I1(n46_adj_3862), .I2(n36_adj_3861), 
            .I3(n3096), .O(n50));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1465 (.I0(n3088), .I1(n42), .I2(n3105), .I3(n3086), 
            .O(n48_adj_3865));
    defparam i21_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n31_adj_3864), .I1(n44_adj_3863), .I2(n3104), 
            .I3(n3101), .O(n49_adj_3866));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1466 (.I0(n3084), .I1(n3089), .I2(n3083), .I3(n3097), 
            .O(n47_adj_3867));
    defparam i20_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1467 (.I0(n47_adj_3867), .I1(n49_adj_3866), .I2(n48_adj_3865), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1467.LUT_INIT = 16'hfffe;
    SB_LUT4 i31235_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36872));
    defparam i31235_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31225_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36862));
    defparam i31225_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31240_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36877));
    defparam i31240_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1468 (.I0(n1502), .I1(n1508), .I2(n1503), .I3(n1506), 
            .O(n18_adj_3868));
    defparam i7_4_lut_adj_1468.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(n1499), .I1(bit_ctr[20]), .I2(n1509), .I3(GND_net), 
            .O(n16_adj_3869));
    defparam i5_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i9_4_lut_adj_1469 (.I0(n1501), .I1(n18_adj_3868), .I2(n1505), 
            .I3(n1500), .O(n20_adj_3870));
    defparam i9_4_lut_adj_1469.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1470 (.I0(n1504), .I1(n20_adj_3870), .I2(n16_adj_3869), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1470.LUT_INIT = 16'hfffe;
    SB_LUT4 i31239_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36876));
    defparam i31239_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25369_4_lut (.I0(n15289), .I1(n30886), .I2(n25921), .I3(\state[0] ), 
            .O(n31001));
    defparam i25369_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut_adj_1471 (.I0(n31001), .I1(\state[1] ), .I2(start), 
            .I3(\neo_pixel_transmitter.done ), .O(n7_adj_3871));
    defparam i20_4_lut_adj_1471.LUT_INIT = 16'hcfcd;
    SB_LUT4 i1_4_lut_adj_1472 (.I0(n22030), .I1(n7_adj_3871), .I2(n15386), 
            .I3(\state[1] ), .O(n29225));
    defparam i1_4_lut_adj_1472.LUT_INIT = 16'hccc4;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17580_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n21950));
    defparam i17580_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1473 (.I0(n1405), .I1(n21950), .I2(n1403), .I3(n1406), 
            .O(n16_adj_3872));
    defparam i6_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1474 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_3873));
    defparam i7_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1475 (.I0(n17_adj_3873), .I1(n1408), .I2(n16_adj_3872), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31238_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36875));
    defparam i31238_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31334 (.I0(bit_ctr[0]), .I1(\color[22] ), 
            .I2(\color[23] ), .I3(bit_ctr[1]), .O(n36894));
    defparam bit_ctr_0__bdd_4_lut_31334.LUT_INIT = 16'he4aa;
    SB_LUT4 n36894_bdd_4_lut (.I0(n36894), .I1(\color[21] ), .I2(\color[20] ), 
            .I3(bit_ctr[1]), .O(n36897));
    defparam n36894_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i471_3_lut_4_lut_4_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(bit_ctr[29]), .I3(GND_net), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_4_lut_4_lut_4_lut_3_lut.LUT_INIT = 16'h4242;
    SB_LUT4 i1_2_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(GND_net), .O(n26372));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h9292;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1476 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_3874));
    defparam i1_2_lut_adj_1476.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_3875));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1477 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_3874), 
            .O(n16_adj_3876));
    defparam i7_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1478 (.I0(n1307), .I1(n16_adj_3876), .I2(n12_adj_3875), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1478.LUT_INIT = 16'hfffe;
    SB_LUT4 i31237_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36874));
    defparam i31237_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1479 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_3877));
    defparam i6_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1480 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_3878));
    defparam i1_3_lut_adj_1480.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1481 (.I0(n9_adj_3878), .I1(n14_adj_3877), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(n22030), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n30800));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i31236_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36873));
    defparam i31236_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29296_2_lut_3_lut (.I0(n22016), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n34325));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29296_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i17594_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n21964));
    defparam i17594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n21964), .I3(n1108), 
            .O(n12_adj_3879));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1482 (.I0(n1107), .I1(n12_adj_3879), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29779_3_lut_4_lut (.I0(\state[1] ), .I1(n35417), .I2(start), 
            .I3(n15289), .O(n35418));
    defparam i29779_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31234_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36871));
    defparam i31234_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut_adj_1483 (.I0(n22016), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n32288));
    defparam i3_4_lut_4_lut_adj_1483.LUT_INIT = 16'h0004;
    SB_LUT4 i14_4_lut_adj_1484 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40));
    defparam i14_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1485 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_3880));
    defparam i18_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1486 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_3881));
    defparam i16_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1487 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_3882));
    defparam i17_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1488 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41));
    defparam i15_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_3883));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43_adj_3882), .I2(n42_adj_3881), 
            .I3(n44_adj_3880), .O(n50_adj_3884));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_3885));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_3885), .I1(n50_adj_3884), .I2(n46_adj_3883), 
            .I3(n38), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31211_2_lut (.I0(n27151), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i31211_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31213_2_lut (.I0(n27151), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i31213_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31233_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36870));
    defparam i31233_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29570_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n16628));
    defparam i29570_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n27151), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut_adj_1489 (.I0(n30953), .I1(n905), .I2(n16628), .I3(GND_net), 
            .O(n8_adj_3886));
    defparam i3_3_lut_adj_1489.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut_adj_1490 (.I0(bit_ctr[26]), .I1(n8_adj_3886), .I2(n906), 
            .I3(n14113), .O(n27151));
    defparam i4_4_lut_adj_1490.LUT_INIT = 16'h040c;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n27151), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14113), .I1(n971[27]), .I2(n27151), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26893_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n32529));
    defparam i26893_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1491 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_3887));
    defparam i2_3_lut_adj_1491.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n27151), .I1(n6_adj_3887), .I2(n1005), .I3(n32529), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i31207_2_lut (.I0(n27151), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_3846));   // verilog/neopixel.v(22[26:36])
    defparam i31207_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14113));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_2_lut_adj_1493 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n14115));
    defparam i1_2_lut_adj_1493.LUT_INIT = 16'h6666;
    SB_LUT4 i29564_3_lut (.I0(n26372), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n30829));
    defparam i29564_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n30837), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_3888));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1494 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_3889));
    defparam i16_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_3890));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1495 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_3891));
    defparam i18_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1496 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_3892));
    defparam i15_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1497 (.I0(n41_adj_3889), .I1(n33_adj_3888), .I2(n2889), 
            .I3(n2901), .O(n46_adj_3893));
    defparam i21_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1498 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39));
    defparam i14_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1499 (.I0(n43_adj_3891), .I1(n2904), .I2(n38_adj_3890), 
            .I3(n2893), .O(n47_adj_3894));
    defparam i22_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1500 (.I0(n47_adj_3894), .I1(n39), .I2(n46_adj_3893), 
            .I3(n40_adj_3892), .O(n2918));
    defparam i24_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i25265_2_lut (.I0(start), .I1(n15289), .I2(GND_net), .I3(GND_net), 
            .O(n30888));
    defparam i25265_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29978_4_lut (.I0(n25921), .I1(n30886), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n35417));
    defparam i29978_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n30888), .I1(n22016), .I2(\state[1] ), .I3(n30886), 
            .O(n30997));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n30997), .I1(n35418), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n31011));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_512 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31232_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36869));
    defparam i31232_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1501 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_3895));
    defparam i16_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1502 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_3896));
    defparam i14_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1503 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_3897));
    defparam i15_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1504 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_3898));
    defparam i13_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_3899));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1505 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_3900));
    defparam i18_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1506 (.I0(n37_adj_3898), .I1(n39_adj_3897), .I2(n38_adj_3896), 
            .I3(n40_adj_3895), .O(n46_adj_3901));
    defparam i22_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_3902));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1507 (.I0(n33_adj_3902), .I1(n46_adj_3901), .I2(n42_adj_3900), 
            .I3(n34_adj_3899), .O(n2819));
    defparam i23_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i31231_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36868));
    defparam i31231_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_3903));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1508 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_3904));
    defparam i15_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i17506_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n21876));
    defparam i17506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1509 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n21876), 
            .O(n36_adj_3905));
    defparam i13_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1510 (.I0(n2700), .I1(n38_adj_3904), .I2(n28_adj_3903), 
            .I3(n2705), .O(n42_adj_3906));
    defparam i19_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1511 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_3907));
    defparam i17_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1512 (.I0(n2687), .I1(n36_adj_3905), .I2(n2703), 
            .I3(n2695), .O(n41_adj_3908));
    defparam i18_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1513 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_3909));
    defparam i16_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1514 (.I0(n39_adj_3909), .I1(n41_adj_3908), .I2(n40_adj_3907), 
            .I3(n42_adj_3906), .O(n2720));
    defparam i22_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 i31230_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36867));
    defparam i31230_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1515 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_3910));
    defparam i14_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1516 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_3911));
    defparam i3_3_lut_adj_1516.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1517 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_3912));
    defparam i12_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1518 (.I0(n25_adj_3911), .I1(n36_adj_3910), .I2(n2594), 
            .I3(n2589), .O(n40_adj_3913));
    defparam i18_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1519 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_3914));
    defparam i16_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_3912), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_3915));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1520 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_3916));
    defparam i15_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1521 (.I0(n37_adj_3916), .I1(n39_adj_3915), .I2(n38_adj_3914), 
            .I3(n40_adj_3913), .O(n2621));
    defparam i21_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17570_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n21940));
    defparam i17570_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1522 (.I0(n3196), .I1(n3208), .I2(n3199), .I3(n3188), 
            .O(n48_adj_3917));
    defparam i20_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1523 (.I0(n3195), .I1(n3202), .I2(n3187), .I3(n3194), 
            .O(n46_adj_3918));
    defparam i18_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1524 (.I0(n3200), .I1(n3185), .I2(n3182), .I3(n3192), 
            .O(n47_adj_3919));
    defparam i19_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1525 (.I0(n3201), .I1(n3197), .I2(n3190), .I3(n3183), 
            .O(n45_adj_3920));
    defparam i17_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1526 (.I0(n3184), .I1(n3205), .I2(n3206), .I3(n3186), 
            .O(n44_adj_3921));
    defparam i16_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1527 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n21940), 
            .O(n43_adj_3922));
    defparam i15_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1528 (.I0(n45_adj_3920), .I1(n47_adj_3919), .I2(n46_adj_3918), 
            .I3(n48_adj_3917), .O(n54_adj_3923));
    defparam i26_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1529 (.I0(n3191), .I1(n3207), .I2(n3204), .I3(n3203), 
            .O(n49_adj_3924));
    defparam i21_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1530 (.I0(n49_adj_3924), .I1(n54_adj_3923), .I2(n43_adj_3922), 
            .I3(n44_adj_3921), .O(n21992));
    defparam i27_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i17646_4_lut (.I0(one_wire_N_449[9]), .I1(n15393), .I2(one_wire_N_449[11]), 
            .I3(one_wire_N_449[10]), .O(n22016));
    defparam i17646_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i229_2_lut (.I0(n22016), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n922));   // verilog/neopixel.v(103[9] 111[12])
    defparam i229_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i25216_4_lut (.I0(n15289), .I1(n25921), .I2(n30886), .I3(\state[0] ), 
            .O(n22030));   // verilog/neopixel.v(36[4] 116[11])
    defparam i25216_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i15_4_lut_adj_1531 (.I0(n22030), .I1(n34325), .I2(\state[1] ), 
            .I3(n15386), .O(n30957));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1531.LUT_INIT = 16'h303a;
    SB_LUT4 i1_4_lut_adj_1532 (.I0(\state[0] ), .I1(n30800), .I2(n922), 
            .I3(\state[1] ), .O(n16527));
    defparam i1_4_lut_adj_1532.LUT_INIT = 16'hafcc;
    SB_LUT4 i1_4_lut_adj_1533 (.I0(\state_3__N_298[1] ), .I1(n36993), .I2(n36897), 
            .I3(bit_ctr[2]), .O(n5_adj_3925));
    defparam i1_4_lut_adj_1533.LUT_INIT = 16'h5044;
    SB_LUT4 i3_4_lut_adj_1534 (.I0(n5_adj_3925), .I1(n3209), .I2(bit_ctr[3]), 
            .I3(n21992), .O(state_3__N_298[0]));
    defparam i3_4_lut_adj_1534.LUT_INIT = 16'h2008;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut_adj_1535 (.I0(bit_ctr[15]), .I1(n18_adj_3849), .I2(n2006), 
            .I3(n2009), .O(n25_adj_3926));
    defparam i9_4_lut_adj_1535.LUT_INIT = 16'hfefc;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut (.I0(n15289), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n30886), .O(n15387));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i1_3_lut_4_lut_adj_1536 (.I0(n25921), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n15289), .O(n919));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_3_lut_4_lut_adj_1536.LUT_INIT = 16'hf3f7;
    SB_LUT4 i15_4_lut_adj_1537 (.I0(n25_adj_3926), .I1(n27_adj_3856), .I2(n26_adj_3851), 
            .I3(n28_adj_3850), .O(n2027));
    defparam i15_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i3557_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n30829), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3557_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[28]), .O(n739));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h29bd;
    SB_LUT4 i25217_2_lut_4_lut (.I0(bit_ctr[28]), .I1(bit_ctr[29]), .I2(bit_ctr[30]), 
            .I3(bit_ctr[31]), .O(n30837));
    defparam i25217_2_lut_4_lut.LUT_INIT = 16'h8208;
    SB_LUT4 i31229_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36866));
    defparam i31229_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1538 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_3927));
    defparam i3_2_lut_adj_1538.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1539 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_3928));
    defparam i13_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1540 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_3929));
    defparam i1_3_lut_adj_1540.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1541 (.I0(n2490), .I1(n34_adj_3928), .I2(n24_adj_3927), 
            .I3(n2494), .O(n38_adj_3930));
    defparam i17_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1542 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_3931));
    defparam i15_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1543 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_3929), 
            .O(n37_adj_3932));
    defparam i16_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1544 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_3933));
    defparam i14_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1545 (.I0(n35_adj_3933), .I1(n37_adj_3932), .I2(n36_adj_3931), 
            .I3(n38_adj_3930), .O(n2522));
    defparam i20_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, GND_net, rx_data, \data_out_frame[20] , \data_out_frame[16] , 
            \data_out_frame[17] , \data_out_frame[18] , \data_out_frame[19] , 
            \data_out_frame[14] , \data_out_frame[5] , \data_out_frame[7] , 
            \data_out_frame[9] , \data_out_frame[11] , \data_out_frame[6] , 
            n37085, \FRAME_MATCHER.state[2] , PWMLimit, control_mode, 
            \FRAME_MATCHER.state[0] , n17214, n17213, n17212, n17211, 
            n17210, n17209, n17208, n17207, n17206, n17205, n17204, 
            \data_out_frame[8] , \data_out_frame[10] , \data_out_frame[15] , 
            \data_out_frame[12] , \data_out_frame[13] , n63, n31, n2421, 
            n13117, n17203, n17202, rx_data_ready, n17201, n17200, 
            n17199, n17198, n30199, n17197, n17196, n17195, n17194, 
            n17193, n17192, n17191, \FRAME_MATCHER.state[3] , n3915, 
            n12917, n17190, n17189, n17188, n17187, n17186, n17185, 
            n17184, \r_SM_Main_2__N_3259[0] , n17183, n17182, n17181, 
            n17180, n17179, n17178, n17177, n17176, n17175, n17174, 
            n17173, n17172, n17171, n17170, n17169, n17168, n17167, 
            n17166, n17165, n17164, n17163, n17162, n17161, n17160, 
            n17159, n17158, n17157, n17156, n17155, n17154, n17153, 
            n17152, n17151, n17150, n17149, n17148, n17147, \data_in[3] , 
            \data_in[0] , \data_in[2] , \data_in[1] , n3761, n22044, 
            n740, n17146, n17145, n17144, n17143, n17142, n17141, 
            n17140, n17139, n17138, n17137, n17136, n17135, n17134, 
            n17133, n15494, n15502, n17132, n15493, n18493, n5, 
            n37539, n17131, n17130, n17129, n17128, n17127, n17126, 
            n17125, n17124, n17123, n17122, n17121, n17120, n17119, 
            n17118, n17117, n17116, n17115, n17114, n17113, n17112, 
            n17111, n17110, n17109, n17108, n17107, n17106, n17105, 
            n17104, n17103, n17102, n17101, n17100, n17099, n17098, 
            n17097, n17096, n17095, n17094, n17093, n17092, n17091, 
            n17090, n17089, n17088, n17087, n17086, \data_out_frame[0][4] , 
            n17085, \data_out_frame[0][3] , n17084, \data_out_frame[0][2] , 
            \Kp[7] , \Kp[6] , \Kp[5] , \Kp[4] , \Kp[3] , \Kp[2] , 
            \Kp[1] , n17076, n17075, n17074, n17073, n17072, n17071, 
            n17070, n17069, n17068, n17067, n15501, n17066, n17065, 
            n17064, n17063, n17062, n17061, n17060, n17059, n17058, 
            n17057, n17056, n17055, n17054, n17053, n17052, n17051, 
            n17050, n17049, n17048, n17047, n17046, n17040, setpoint, 
            n17039, n17038, n17037, n17036, n17035, n17034, n17033, 
            n17032, n17031, n17030, n17029, n17028, n17027, n17026, 
            n17025, n17024, n17023, n17022, n17021, n17020, n17019, 
            gearBoxRatio, n16770, n17018, LED_c, n29611, \Kp[0] , 
            n16899, n4335, n4312, n4334, n4333, n4332, n4331, 
            n4330, n4329, n4328, n4327, n4326, n4325, n4324, n4323, 
            n4322, n4321, n4320, n4319, n4318, n4317, n4316, n4315, 
            n4314, n31259, n4313, n15495, n5_adj_3, tx_active, n16549, 
            VCC_net, tx_o, tx_enable, n16816, r_Bit_Index, n16819, 
            n29853, r_SM_Main, \r_SM_Main_2__N_3185[2] , r_Rx_Data, 
            PIN_13_N_65, n16600, n16687, n4573, n17013, n16841, 
            n16840, n16839, n16835, n16825, n16824, n16823, n21347, 
            n4, n4_adj_4, n15244, n15373, n4_adj_5) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input GND_net;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[6] ;
    input n37085;
    output \FRAME_MATCHER.state[2] ;
    output [23:0]PWMLimit;
    output [7:0]control_mode;
    output \FRAME_MATCHER.state[0] ;
    input n17214;
    input n17213;
    input n17212;
    input n17211;
    input n17210;
    input n17209;
    input n17208;
    input n17207;
    input n17206;
    input n17205;
    input n17204;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    output n63;
    input n31;
    output n2421;
    output n13117;
    input n17203;
    input n17202;
    output rx_data_ready;
    input n17201;
    input n17200;
    input n17199;
    input n17198;
    output n30199;
    input n17197;
    input n17196;
    input n17195;
    input n17194;
    input n17193;
    input n17192;
    input n17191;
    output \FRAME_MATCHER.state[3] ;
    output n3915;
    output n12917;
    input n17190;
    input n17189;
    input n17188;
    input n17187;
    input n17186;
    input n17185;
    input n17184;
    output \r_SM_Main_2__N_3259[0] ;
    input n17183;
    input n17182;
    input n17181;
    input n17180;
    input n17179;
    input n17178;
    input n17177;
    input n17176;
    input n17175;
    input n17174;
    input n17173;
    input n17172;
    input n17171;
    input n17170;
    input n17169;
    input n17168;
    input n17167;
    input n17166;
    input n17165;
    input n17164;
    input n17163;
    input n17162;
    input n17161;
    input n17160;
    input n17159;
    input n17158;
    input n17157;
    input n17156;
    input n17155;
    input n17154;
    input n17153;
    input n17152;
    input n17151;
    input n17150;
    input n17149;
    input n17148;
    input n17147;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[1] ;
    output n3761;
    output n22044;
    output n740;
    input n17146;
    input n17145;
    input n17144;
    input n17143;
    input n17142;
    input n17141;
    input n17140;
    input n17139;
    input n17138;
    input n17137;
    input n17136;
    input n17135;
    input n17134;
    input n17133;
    output n15494;
    output n15502;
    input n17132;
    output n15493;
    output n18493;
    output n5;
    output n37539;
    input n17131;
    input n17130;
    input n17129;
    input n17128;
    input n17127;
    input n17126;
    input n17125;
    input n17124;
    input n17123;
    input n17122;
    input n17121;
    input n17120;
    input n17119;
    input n17118;
    input n17117;
    input n17116;
    input n17115;
    input n17114;
    input n17113;
    input n17112;
    input n17111;
    input n17110;
    input n17109;
    input n17108;
    input n17107;
    input n17106;
    input n17105;
    input n17104;
    input n17103;
    input n17102;
    input n17101;
    input n17100;
    input n17099;
    input n17098;
    input n17097;
    input n17096;
    input n17095;
    input n17094;
    input n17093;
    input n17092;
    input n17091;
    input n17090;
    input n17089;
    input n17088;
    input n17087;
    input n17086;
    output \data_out_frame[0][4] ;
    input n17085;
    output \data_out_frame[0][3] ;
    input n17084;
    output \data_out_frame[0][2] ;
    output \Kp[7] ;
    output \Kp[6] ;
    output \Kp[5] ;
    output \Kp[4] ;
    output \Kp[3] ;
    output \Kp[2] ;
    output \Kp[1] ;
    input n17076;
    input n17075;
    input n17074;
    input n17073;
    input n17072;
    input n17071;
    input n17070;
    input n17069;
    input n17068;
    input n17067;
    output n15501;
    input n17066;
    input n17065;
    input n17064;
    input n17063;
    input n17062;
    input n17061;
    input n17060;
    input n17059;
    input n17058;
    input n17057;
    input n17056;
    input n17055;
    input n17054;
    input n17053;
    input n17052;
    input n17051;
    input n17050;
    input n17049;
    input n17048;
    input n17047;
    input n17046;
    input n17040;
    output [23:0]setpoint;
    input n17039;
    input n17038;
    input n17037;
    input n17036;
    input n17035;
    input n17034;
    input n17033;
    input n17032;
    input n17031;
    input n17030;
    input n17029;
    input n17028;
    input n17027;
    input n17026;
    input n17025;
    input n17024;
    input n17023;
    input n17022;
    input n17021;
    input n17020;
    input n17019;
    output [23:0]gearBoxRatio;
    input n16770;
    input n17018;
    output LED_c;
    input n29611;
    output \Kp[0] ;
    input n16899;
    output n4335;
    output n4312;
    output n4334;
    output n4333;
    output n4332;
    output n4331;
    output n4330;
    output n4329;
    output n4328;
    output n4327;
    output n4326;
    output n4325;
    output n4324;
    output n4323;
    output n4322;
    output n4321;
    output n4320;
    output n4319;
    output n4318;
    output n4317;
    output n4316;
    output n4315;
    output n4314;
    output n31259;
    output n4313;
    output n15495;
    output n5_adj_3;
    output tx_active;
    output n16549;
    input VCC_net;
    output tx_o;
    output tx_enable;
    input n16816;
    output [2:0]r_Bit_Index;
    input n16819;
    input n29853;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3185[2] ;
    output r_Rx_Data;
    input PIN_13_N_65;
    output n16600;
    output n16687;
    output n4573;
    input n17013;
    input n16841;
    input n16840;
    input n16839;
    input n16835;
    input n16825;
    input n16824;
    input n16823;
    output n21347;
    output n4;
    output n4_adj_4;
    output n15244;
    output n15373;
    output n4_adj_5;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n17302;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    
    wire n30651, n30624;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    
    wire n6, n30326, n17301;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    
    wire n17346;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n17345, n17344, n17343, n17342, n24669;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n24670, n17341;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    
    wire n17257;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    
    wire n17340, n17339, n17338, n17337, n17336, n17335, n17334, 
        n2, n24668, n1731, n10, n31262;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    
    wire n17275, n17256, n17255, n17314;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n17313, n2_adj_3533, n3, n17254, n17312, n2_adj_3534, n24667, 
        n17276, n2_adj_3535, n24666, n17277, n17311, n17253;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n34170, n17260, n17259, n17252, n17251;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n19, n16, n17250, n2_adj_3536, n24665, n17, n34171, n19_adj_3537, 
        n16217, n30612, n30371, n31387, n16_adj_3538, n17_adj_3539, 
        n34172, n19_adj_3540, n30767, n30434, n17249, n30793, n30294, 
        n30579, n16_adj_3541, n17_adj_3542, n34175, n19_adj_3543, 
        n15054, n16246, n30392, n15781, n27248, n15636, n30734, 
        n11, n5_c, n34176, n16377, n17248, n17247, n27165, n30507;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    
    wire n27171, n17246, n17245;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    
    wire n17244, n17243, n30663, n15880, n30407, n6_adj_3544, n17242, 
        n17241, n17240, n17239, n17238, n17237;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    
    wire n31_c, n21283;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n4311, n17236, n17235, n16356, n30645, n27173, n18, n17234, 
        n17233, n17521, n17520, n17232, n17519, n17518, n17517, 
        n29349, n16862, n17231, n26497, n30513, n17230, n17229;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    
    wire n29343, n17228, n17419, n17418, n17417, n17416, n17415, 
        n17414, n17413, n2_adj_3545, n24664, n17412, n17411, n17410, 
        n17409, n17408, n17407, n17406, n17405, n17404, n17403, 
        n17402, n17401, n17400, n17399, n17398, n17397, n17396, 
        n17395, n17394, n17393, n17392, tx_transmit_N_3151, n22052, 
        n17391, n17390, n17389;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n17388, n17387, n17386, n17385, n17384, n17383, n17382, 
        n17381;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n17380, n17379, n17378, n17377, n17376, n17375, n17374, 
        n17373;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    
    wire n17372, n17371, n17370, n17369, n17368, n17367, n17366, 
        n17365;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    
    wire n17364, n17363, n17362, n17361, n17360, n17359, n17358, 
        n17357, n17356, n17355, n17354, n17353, n17352, n17351, 
        n17350, n17349, n17348, n30568, n30716, n17347, n17310, 
        n17300, n17299, n17298, n17297, n17296, n17295, n17294, 
        n17227, n17226, n17225, n17224, n17223, n17222, n17221;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n17220, n17219, n17218, n17217, n17216, n17215, n17309, 
        n30698, n27213, n14, n15541, n30764, n15624, n30441, n30302, 
        n17293;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    
    wire n16_adj_3546, n30657, n16491, n11438;
    wire [7:0]n2236;
    
    wire n17_adj_3547, n17292, n27271, n15085, n31193, n30450, n6_adj_3548, 
        n17291, n17290, n17289, n17288, n34278, n26563, n32127, 
        n31605, n30601, n19_adj_3549, n32547, n32548, n16214, n30582, 
        n32551, n30284, n30701, n32550, n32544, n32545, n32542, 
        n10_adj_3550, n30187;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n17326, n32541, n17327, n17328, n17329, n17330, n17331, 
        n17332, n17333;
    wire [31:0]n93;
    
    wire n29603, n10_adj_3552, n30172, n63_adj_3553, n63_adj_3554, 
        n61, n133, n1, n29637, n29639, n17287, n29641, n29643, 
        n29645, n6_adj_3555, n29667, n29623, n29597, n29647, n2_adj_3556, 
        n24663, n29621, n5_adj_3557, n17286, n32644, n32559, n37011, 
        n32561, n29649, n29651, n29653, n29619, n29617, n29655, 
        n54, n67, n7, n29797, n7_adj_3558, n29793, n7_adj_3559, 
        n7_adj_3560, n29789, n29785, n17285;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    
    wire n2430, n3_adj_3561, n7_adj_3562, n29781, n29777, n12, n26493, 
        n29801, n2_adj_3563, n24662, n29773, n7_adj_3564, \FRAME_MATCHER.rx_data_ready_prev , 
        n7_adj_3565, n2_adj_3566, n24661, n7_adj_3567, n7_adj_3568, 
        n21272, n10_adj_3569, Kp_23__N_832, n30784, Kp_23__N_794, 
        n30368, n30704, n15894, n56, n17308, n17303, n29769, n21813, 
        n29765, n30575, n29761, n30545, n29757, n29753, n30176, 
        n29749, n29745, n2_adj_3570, n24660, n29741, n29733, n21802, 
        n21274, n21790, n29565, n29545, n29543, n17307, n29541, 
        n29539, n30190, n17318, n17319, n17320, n17321, n17322, 
        n17323, n17324, n17325, n2_adj_3571, n24659, Kp_23__N_1289, 
        n2_adj_3572, n24658;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    
    wire n15671, n10_adj_3573, n30404, n15772, n30631, n30221, n15587, 
        n14_adj_3574, n16139, n10_adj_3575, n16302, Kp_23__N_1405, 
        n2_adj_3576, n24657, n15264, n15224, n10_adj_3577, n2_adj_3578, 
        n24656, n17306, Kp_23__N_962, n16_adj_3579, n2_adj_3580, n24655, 
        n2_adj_3581, n24654, n15824, n2_adj_3582, n24653, n2_adj_3583, 
        n24652, n34257, n24688, n24687, n34256, n24686, n22, n24651, 
        n34258, n24685, n21292, n22062, n50, n34460, n34462, n47, 
        n22054, n4_c, n32519, n38, n39, n37, n32515, n46, n32517;
    wire [31:0]\FRAME_MATCHER.state_31__N_2428 ;
    
    wire n5784, n34255, n24684, n30266, n30675, n6_adj_3584, n27227, 
        n27225, n30504, n26717, n16149, n26948, n30672, n30591, 
        n16255, n16360, n6_adj_3585, n30707, Kp_23__N_1280, n27261, 
        n30491, n26635, n30341, n22_adj_3586, n30510, n24, n23, 
        n25, n15982, n30660, n30483, n13, n15, n14_adj_3587, n30494, 
        n30678, n30235, n30542, n30539, n30420, n14_adj_3588, n30740, 
        n10_adj_3589, n16321, n164, n26401, n30648, n8, n16262, 
        n30469, n30600, n27234, n32089, Kp_23__N_829, n30498, n6_adj_3590, 
        Kp_23__N_1498, n30737, n30722, n30725, n16_adj_3591, n15_adj_3592, 
        n14_adj_3593, n30212, n14_adj_3594, n30263, n30554, n15_adj_3595, 
        n15790, n15573, n30480, n10_adj_3596, n26712, n14_adj_3597, 
        n15697, n15_adj_3598, n15604, n30606, n30397, n30790, n15746, 
        n10_adj_3599, n30232, Kp_23__N_1327, n30710, n30758, n30291, 
        n7_adj_3600, n16098, n16_adj_3601, n30356, n30628, n17_adj_3602, 
        n15525, n30393, n4_adj_3603, n8_adj_3604, Kp_23__N_1019, n12_adj_3605, 
        n30519, n16094, n10_adj_3606, n14_adj_3607, n15704, n30455, 
        n15557, n30205, n16067, n15753, n14_adj_3608, n15_adj_3609, 
        n30414, n16146, n30340, n27276, n26388, n30666, n30288, 
        n30452, n15844, n6_adj_3610, n30609, n16208, n15994, n15677, 
        n14_adj_3611, Kp_23__N_823, n30536, n15725, n30180, n16901, 
        n30429, n7_adj_3612, n30353, n27175, n16114, n14_adj_3613, 
        n15_adj_3614, n30336, n6_adj_3615, n30374, n6_adj_3616, n30426, 
        n4_adj_3617, n30807, n34331, n15_adj_3618, n28, n26, n27, 
        n25_adj_3619, n30093, n30201, n6_adj_3620, n234, n30203, 
        n63_adj_3621, n30254, n34, n58, n56_adj_3622, n57, n30458, 
        n55, n52, n30778, n54_adj_3623, n30359, n53, n64, n30528, 
        n59, n14_adj_3624, n14_adj_3625, n24683, n13_adj_3626, n13_adj_3627, 
        n16_adj_3628, n17_adj_3629, n12_adj_3630, n31718, n31188, 
        n26767, n26452, n31425, n31345, n6_adj_3631, n14_adj_3632, 
        n26930, n5_adj_3633, n13_adj_3634, n10_adj_3635, n31451, n32479, 
        n14_adj_3636, n30603, n15_adj_3637, n31682, n30329, n26405, 
        n31191, n31442, n30595, n30474, n18_adj_3638, n31180, n32525, 
        n26_adj_3639, n27_adj_3640, n30516, n25_adj_3641, n31_adj_3642, 
        n24682, n18507, n12846, n34330, n2_adj_3643, n24681, n2_adj_3644, 
        n24680, n2_adj_3645, n24679, n2_adj_3646, n24678, n6_adj_3647, 
        n15369, n2_adj_3648, n5_adj_3649, n10_adj_3650, n14_adj_3651, 
        n15283, n16_adj_3652, n37044, n37047, n37038, n37041, n15355, 
        n17_adj_3653, n15427, n16_adj_3654, n17_adj_3655, n20, n10_adj_3656, 
        n15421, n37026, n2_adj_3657, n24677, n37029, n37020, n37023, 
        n37014, n37017, n37008, n21899, n15239, n4_adj_3658, n36996, 
        n36999, n36984, n36978, n36981, n15358, n6_adj_3659, n63_adj_3660, 
        n42, n40, n41, n39_adj_3661, n38_adj_3662, n37_adj_3663, 
        n36972, n36975, n36966, n36969, n36960, n48, n43, n10_adj_3664, 
        n15424, n7_adj_3665, n32465, n10_adj_3666, n14_adj_3667, n16_adj_3668, 
        n22_adj_3669, n20_adj_3670, n24_adj_3671, n2857, n15504, n2_adj_3673, 
        n24676, n17278, n21269, n17_adj_3674, n16_adj_3675, n36963, 
        n17279, n2_adj_3676, n24675, n17262, n17280, n17281, n2_adj_3677, 
        n24674, n2_adj_3678, n24673, n17284, n17283, n17282, n3_adj_3679, 
        n3_adj_3680, n3_adj_3681, n3_adj_3682, n3_adj_3683, n3_adj_3684, 
        n3_adj_3685, n3_adj_3686, n3_adj_3687, n3_adj_3688, n3_adj_3689, 
        n3_adj_3690, n3_adj_3691, n3_adj_3692, n3_adj_3693, n3_adj_3694, 
        n3_adj_3695, n2_adj_3696, n3_adj_3697, n2_adj_3698, n3_adj_3699, 
        n2_adj_3700, n3_adj_3701, n2_adj_3702, n3_adj_3703, n3_adj_3704, 
        n3_adj_3705, n3_adj_3706, n3_adj_3707, n3_adj_3708, n3_adj_3709, 
        n3_adj_3710, n3_adj_3711, n3_adj_3712, n16553, n31499, n31154, 
        n31813, n31828, n31232, n31697, n31402, n32201, n32039, 
        n31333, n31184, n30323, n30344, n31393, n37190, n29613, 
        n29609, n8_adj_3713, n8_adj_3714, n8_adj_3715, n8_adj_3716, 
        n24672, n10_adj_3717, n30362, n19_adj_3718, n34169, n36954, 
        n10_adj_3719, n17083, n17082, n17081, n17080, n17079, n17078, 
        n17077, n17274, n17305, n24_adj_3720, n17273, n17272, n17271, 
        n17270, n17304, n17_adj_3721, n16_adj_3722, n36957, n14_adj_3723, 
        n24671, n10_adj_3724, n6_adj_3725, n15361, n36948, n36951, 
        n17261, n17269, n17268, n17267, n17266, n17265, n17317, 
        n17258, n16772, n16318, n12_adj_3726, n16967, n16966, n16965, 
        n16964, n16963, n16962, n16961, n16960, n16959, n16958, 
        n16957, n16956, n16955, n16954, n16953, n16952, n16951, 
        n16950, n16949, n16948, n16947, n16946, n16944, n30948, 
        n30168, n16903, n16902, n16900, n30634, n17264, n17263, 
        n17316, n17315, n10_adj_3727, n30164, n36942, n36945, n36936, 
        n36939, n36930, n36933, n36924, n36927, n36918, n36921, 
        n36912, n30522, n1237, n36915, n36906, n36909, n15506, 
        n36900, n36903, n10_adj_3728, n36882, n30548, n30365, n36885, 
        n6_adj_3729, n15863, n30224, n27167, n30781, n30588, n6_adj_3730, 
        n30770, n30559, n30315, n30695, n21540, n18518, n15630, 
        n6_adj_3731, n16_adj_3732, n6_adj_3733, n10_adj_3734, n30565, 
        n30572, n30322, n26487;
    wire [31:0]\FRAME_MATCHER.state_31__N_2396 ;
    
    wire n961, n30417, n30594, n19_adj_3736, n34853, n5_adj_3737, 
        n32539, n32540, n32577, n32579, n32578, n19_adj_3738, n34849, 
        n5_adj_3739, n32536, n32537, n32574, n32576, n32575, n34844, 
        n5_adj_3740, n32571, n32573, n32572, n35797, n36987, n35801;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n34271, n6_adj_3741, n5_adj_3742, n32568, n32570, n32569, 
        n34268, n6_adj_3743, n5_adj_3744, n32565, n32567, n32566, 
        n34825, n5_adj_3745, n32562, n32564, n16_adj_3746, n5782, 
        n30761, n17_adj_3747, n32330, n13185, n7_adj_3748, n30890, 
        n5_adj_3749, n6_adj_3750, n30343, n16389, n10_adj_3751, n30691, 
        n30257, n16_adj_3752, n30447, n30752, n17_adj_3753, n30298, 
        n15760, n26362, n18_adj_3754, n26378, n30435, n20_adj_3755, 
        n15_adj_3756, n12_adj_3757, n15034, n27257, n13_adj_3758, 
        n32059, n16042, n2_adj_3759, n30787, n30208, n8_adj_3760, 
        n30728, n30438, n12_adj_3761, n6_adj_3762, n30731, n30350, 
        n6_adj_3763, n10_adj_3764, n27001, n30746, n30486, n12_adj_3765, 
        n30617, n1595, n30533, n30669, n6_adj_3766, n31361, n30501, 
        n15532, n15986, n1967, n18_adj_3767, n30743, n20_adj_3768, 
        n30681, n30377, n30597, n30333, n27179, n30585, n15_adj_3769, 
        n15766, n30281, n12_adj_3770, n30749, n30687, n30276, n30637, 
        n30562, n12_adj_3771, n30260, n30461, n7_adj_3772, n18_adj_3773, 
        n16_adj_3774, n20_adj_3775, n30525, n30218, n12_adj_3776, 
        n26562, n30384, n30684, n30318, n6_adj_3777, n30551, n15651, 
        n30719, n30465, n16226, n16426, n30444, n12_adj_3778, n30381, 
        n15886, n30305, n16335, n10_adj_3779, n30411, n30250, n14_adj_3780, 
        n1112, n1256, n13_adj_3781, n14_adj_3782, n13_adj_3783, n12_adj_3784, 
        n16_adj_3785, n17_adj_3786, n32150, n30, n28_adj_3787, n29, 
        n27_adj_3788, n32152, n54_adj_3789, n52_adj_3790, n53_adj_3791, 
        n51, n48_adj_3792, n50_adj_3793, n16048, n49, n60, n55_adj_3794, 
        n14_adj_3795, n31635, n12_adj_3796;
    
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n17302));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut (.I0(n30651), .I1(n30624), .I2(\data_in_frame[13] [5]), 
            .I3(n6), .O(n30326));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n17301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n17346));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n17345));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n17344));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n17343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n17342));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_21 (.CI(n24669), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n24670));
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n17341));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n17340));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n17339));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n17338));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n17337));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n17336));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n17335));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n17334));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_20_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n24668), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12888_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n17275));
    defparam i12888_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n17314));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n17313));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3533), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17254));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_20 (.CI(n24668), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n24669));
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n17312));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_19_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n24667), .O(n2_adj_3534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_19 (.CI(n24667), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n24668));
    SB_LUT4 i12889_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n17276));
    defparam i12889_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_44_18_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n24666), .O(n2_adj_3535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_18 (.CI(n24666), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n24667));
    SB_LUT4 i12890_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n17277));
    defparam i12890_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n17311));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17253));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i29206_2_lut (.I0(\data_out_frame[22] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34170));
    defparam i29206_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17252));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17251));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17250));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_17_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n24665), .O(n2_adj_3536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29201_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34171));
    defparam i29201_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3537));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(n16217), .I1(n30612), .I2(\data_out_frame[18] [6]), 
            .I3(n30371), .O(n31387));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3538));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3539));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29198_2_lut (.I0(\data_out_frame[22] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34172));
    defparam i29198_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3540));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[14] [4]), .I1(n30767), .I2(\data_out_frame[16] [5]), 
            .I3(GND_net), .O(n30434));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17249));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_861 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n30793));
    defparam i1_2_lut_3_lut_adj_861.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_862 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(n30294), .I3(\data_out_frame[11] [7]), .O(n30579));
    defparam i2_3_lut_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3541));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3542));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28882_2_lut (.I0(\data_out_frame[22] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34175));
    defparam i28882_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3543));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_863 (.I0(\data_out_frame[14] [7]), .I1(n15054), 
            .I2(n16246), .I3(GND_net), .O(n30392));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_863.LUT_INIT = 16'h9696;
    SB_LUT4 i4_3_lut_4_lut (.I0(n15781), .I1(n27248), .I2(n15636), .I3(n30734), 
            .O(n11));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29187_2_lut (.I0(\data_out_frame[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34176));
    defparam i29187_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_864 (.I0(\data_out_frame[14] [7]), .I1(n15054), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n16377));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_864.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17247));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_865 (.I0(n27165), .I1(n30507), .I2(\data_in_frame[17] [7]), 
            .I3(GND_net), .O(n27171));
    defparam i1_2_lut_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17246));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17245));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17243));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_866 (.I0(n27165), .I1(n30507), .I2(\data_in_frame[17] [6]), 
            .I3(GND_net), .O(n30663));
    defparam i1_2_lut_3_lut_adj_866.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n15880), .I1(n30407), .I2(n16246), 
            .I3(\data_out_frame[16] [7]), .O(n6_adj_3544));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17237));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_867 (.I0(n31_c), .I1(n21283), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n4311));
    defparam i1_2_lut_3_lut_adj_867.LUT_INIT = 16'h1010;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17236));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17235));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_868 (.I0(n16356), .I1(n30645), .I2(n27173), 
            .I3(GND_net), .O(n18));
    defparam i1_2_lut_3_lut_adj_868.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17233));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n17521));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n17520));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n17232));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n17519));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n17518));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n17517));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n29349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n16862));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n17231));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_869 (.I0(n16356), .I1(n30645), .I2(n26497), 
            .I3(GND_net), .O(n30513));
    defparam i1_2_lut_3_lut_adj_869.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n17230));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17229));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_17 (.CI(n24665), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n24666));
    SB_DFF byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
           .D(n29343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17228));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(clk32MHz), 
           .D(n37085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n17419));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n17418));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n17417));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n17416));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n17415));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n17414));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n17413));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_16_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n24664), .O(n2_adj_3545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n17412));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n17411));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n17410));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n17409));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n17408));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n17407));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n17406));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n17405));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n17404));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n17403));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n17402));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n17401));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n17400));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n17399));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n17398));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n17397));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n17396));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n17395));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n17394));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n17393));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n17392));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_657_i1_3_lut_4_lut (.I0(n31_c), .I1(n21283), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(tx_transmit_N_3151), .O(n22052));
    defparam mux_657_i1_3_lut_4_lut.LUT_INIT = 16'h0efe;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n17391));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n17390));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n17389));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n17388));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n17387));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n17386));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n17385));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n17384));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n17383));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n17382));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n17381));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n17380));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n17379));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n17378));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n17377));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n17376));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n17375));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n17374));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n17373));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n17372));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n17371));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n17370));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n17369));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n17368));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n17367));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n17366));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n17365));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n17364));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n17363));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n17362));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n17361));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n17360));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n17359));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n17358));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n17357));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n17356));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n17355));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n17354));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n17353));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n17352));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n17351));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n17350));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n17349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n17348));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_870 (.I0(n16356), .I1(n30645), .I2(n30612), 
            .I3(n30568), .O(n30716));
    defparam i2_3_lut_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n17347));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n17310));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n17300));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n17299));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n17298));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n17297));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n17296));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n17295));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n17294));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17227));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17226));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17225));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17224));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17223));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17222));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17221));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17220));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17219));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17218));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17217));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17216));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17215));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17214));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17213));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n17309));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17212));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17211));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[16] [7]), .I1(n16246), .I2(n30698), 
            .I3(n27213), .O(n14));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17210));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17209));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_871 (.I0(\data_out_frame[17] [0]), .I1(n15541), 
            .I2(\data_out_frame[18] [7]), .I3(n30407), .O(n30764));
    defparam i2_3_lut_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_872 (.I0(n15624), .I1(\data_out_frame[17] [4]), 
            .I2(n30441), .I3(GND_net), .O(n30302));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_3_lut_adj_872.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n17293));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3546));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_873 (.I0(n15624), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n30657));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_3_lut_adj_873.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut (.I0(n16491), .I1(n11438), .I2(n2236[1]), .I3(byte_transmit_counter[1]), 
            .O(n16862));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17208));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17207));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3547));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17206));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut_4_lut_adj_874 (.I0(n16491), .I1(n11438), .I2(n2236[6]), 
            .I3(byte_transmit_counter[6]), .O(n17520));
    defparam i1_4_lut_4_lut_adj_874.LUT_INIT = 16'hd580;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17205));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17204));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n17292));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_875 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [1]), 
            .I2(n27271), .I3(n15085), .O(n31193));
    defparam i2_3_lut_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_876 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [1]), 
            .I2(n30450), .I3(GND_net), .O(n6_adj_3548));
    defparam i1_2_lut_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n17291));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n17290));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n17289));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n17288));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i29243_2_lut (.I0(\data_out_frame[22] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34278));
    defparam i29243_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_877 (.I0(n26563), .I1(n32127), .I2(n31605), 
            .I3(n30601), .O(n30507));
    defparam i2_3_lut_4_lut_adj_877.LUT_INIT = 16'h9669;
    SB_CARRY add_44_16 (.CI(n24664), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n24665));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3549));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26910_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32547));
    defparam i26910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26911_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32548));
    defparam i26911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_878 (.I0(n15624), .I1(n16214), .I2(\data_out_frame[17] [5]), 
            .I3(GND_net), .O(n30582));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_878.LUT_INIT = 16'h9696;
    SB_LUT4 i26914_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32551));
    defparam i26914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_879 (.I0(n15624), .I1(n16214), .I2(n30284), 
            .I3(\data_out_frame[20] [0]), .O(n30701));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i26913_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32550));
    defparam i26913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26907_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32544));
    defparam i26907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26908_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32545));
    defparam i26908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26905_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32542));
    defparam i26905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12939_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n17326));
    defparam i12939_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i26904_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n32541));
    defparam i26904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12940_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n17327));
    defparam i12940_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12941_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n17328));
    defparam i12941_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12942_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n17329));
    defparam i12942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12943_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n17330));
    defparam i12943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12944_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n17331));
    defparam i12944_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12945_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n17332));
    defparam i12945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12946_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30187), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n17333));
    defparam i12946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut (.I0(n93[1]), .I1(n63), .I2(n31), .I3(n2421), 
            .O(n29603));   // verilog/coms.v(143[4] 146[7])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hbbb0;
    SB_LUT4 i12971_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n17358));
    defparam i12971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_880 (.I0(n63_adj_3553), .I1(n63_adj_3554), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n93[1]));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_880.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_881 (.I0(n63_adj_3553), .I1(n63_adj_3554), 
            .I2(n63), .I3(GND_net), .O(n13117));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_881.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [28]), 
            .O(n29637));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_882 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [25]), 
            .O(n29639));
    defparam i1_2_lut_4_lut_adj_882.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n17287));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_883 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [24]), 
            .O(n29641));
    defparam i1_2_lut_4_lut_adj_883.LUT_INIT = 16'hfe00;
    SB_LUT4 i12972_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n17359));
    defparam i12972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_884 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [22]), 
            .O(n29643));
    defparam i1_2_lut_4_lut_adj_884.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_885 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [21]), 
            .O(n29645));
    defparam i1_2_lut_4_lut_adj_885.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3555));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'ha300;
    SB_LUT4 i1_2_lut_4_lut_adj_886 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [20]), 
            .O(n29667));
    defparam i1_2_lut_4_lut_adj_886.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_887 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [19]), 
            .O(n29623));
    defparam i1_2_lut_4_lut_adj_887.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_888 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [13]), 
            .O(n29597));
    defparam i1_2_lut_4_lut_adj_888.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_889 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [12]), 
            .O(n29647));
    defparam i1_2_lut_4_lut_adj_889.LUT_INIT = 16'hfe00;
    SB_LUT4 add_44_15_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n24663), .O(n2_adj_3556)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_890 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [10]), 
            .O(n29621));
    defparam i1_2_lut_4_lut_adj_890.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3557));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n17286));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i26922_3_lut (.I0(n5_adj_3557), .I1(n6_adj_3555), .I2(n32644), 
            .I3(GND_net), .O(n32559));
    defparam i26922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26924_4_lut (.I0(n32559), .I1(n37011), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32561));
    defparam i26924_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_891 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [9]), 
            .O(n29649));
    defparam i1_2_lut_4_lut_adj_891.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_892 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [8]), 
            .O(n29651));
    defparam i1_2_lut_4_lut_adj_892.LUT_INIT = 16'hfe00;
    SB_LUT4 i12973_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n17360));
    defparam i12973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12974_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n17361));
    defparam i12974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17203));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_893 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [7]), 
            .O(n29653));
    defparam i1_2_lut_4_lut_adj_893.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_894 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [6]), 
            .O(n29619));
    defparam i1_2_lut_4_lut_adj_894.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_895 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [5]), 
            .O(n29617));
    defparam i1_2_lut_4_lut_adj_895.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_896 (.I0(n61), .I1(n133), .I2(n1), .I3(\FRAME_MATCHER.state [4]), 
            .O(n29655));
    defparam i1_2_lut_4_lut_adj_896.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_897 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_3_lut_adj_897.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_898 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n29797));
    defparam i1_2_lut_3_lut_adj_898.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_899 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n7_adj_3558));
    defparam i1_2_lut_3_lut_adj_899.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_900 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n29793));
    defparam i1_2_lut_3_lut_adj_900.LUT_INIT = 16'he0e0;
    SB_LUT4 i12975_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n17362));
    defparam i12975_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12976_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n17363));
    defparam i12976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_901 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n7_adj_3559));
    defparam i1_2_lut_3_lut_adj_901.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_902 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n7_adj_3560));
    defparam i1_2_lut_3_lut_adj_902.LUT_INIT = 16'he0e0;
    SB_LUT4 i12977_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n17364));
    defparam i12977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17202));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12978_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30172), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n17365));
    defparam i12978_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_903 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n29789));
    defparam i1_2_lut_3_lut_adj_903.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_904 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n29785));
    defparam i1_2_lut_3_lut_adj_904.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n17285));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_330_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3561));
    defparam select_330_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_905 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n7_adj_3562));
    defparam i1_2_lut_3_lut_adj_905.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_906 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n29781));
    defparam i1_2_lut_3_lut_adj_906.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_907 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n29777));
    defparam i1_2_lut_3_lut_adj_907.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(n12), .I3(\data_in_frame[0] [5]), .O(n26493));   // verilog/coms.v(76[16:27])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_44_15 (.CI(n24663), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n24664));
    SB_LUT4 i1_2_lut_3_lut_adj_908 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n29801));
    defparam i1_2_lut_3_lut_adj_908.LUT_INIT = 16'he0e0;
    SB_LUT4 add_44_14_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n24662), .O(n2_adj_3563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_909 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n29773));
    defparam i1_2_lut_3_lut_adj_909.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_910 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n7_adj_3564));
    defparam i1_2_lut_3_lut_adj_910.LUT_INIT = 16'he0e0;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_14 (.CI(n24662), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n24663));
    SB_LUT4 i1_2_lut_3_lut_adj_911 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n7_adj_3565));
    defparam i1_2_lut_3_lut_adj_911.LUT_INIT = 16'he0e0;
    SB_LUT4 add_44_13_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n24661), .O(n2_adj_3566)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_912 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n7_adj_3567));
    defparam i1_2_lut_3_lut_adj_912.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17201));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_913 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n7_adj_3568));
    defparam i1_2_lut_3_lut_adj_913.LUT_INIT = 16'he0e0;
    SB_LUT4 i16908_2_lut_3_lut (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n21272));
    defparam i16908_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_4_lut_adj_914 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [1]), .I3(n10_adj_3569), .O(Kp_23__N_832));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_915 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(n30784), .I3(Kp_23__N_794), .O(n30368));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_916 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(n30704), .I3(Kp_23__N_794), .O(n15894));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_917 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_3_lut_adj_917.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n17308));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n17303));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_13 (.CI(n24661), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n24662));
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17199));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_918 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n29769));
    defparam i1_2_lut_3_lut_adj_918.LUT_INIT = 16'he0e0;
    SB_LUT4 i17444_1_lut (.I0(n21813), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1731));
    defparam i17444_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_919 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n29765));
    defparam i1_2_lut_3_lut_adj_919.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_920 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n30575));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_921 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n29761));
    defparam i1_2_lut_3_lut_adj_921.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_922 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n30545));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_922.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_923 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n29757));
    defparam i1_2_lut_3_lut_adj_923.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_924 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n29753));
    defparam i1_2_lut_3_lut_adj_924.LUT_INIT = 16'he0e0;
    SB_LUT4 i12963_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n17350));
    defparam i12963_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_925 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n29749));
    defparam i1_2_lut_3_lut_adj_925.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_926 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n29745));
    defparam i1_2_lut_3_lut_adj_926.LUT_INIT = 16'he0e0;
    SB_LUT4 i12964_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n17351));
    defparam i12964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_12_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n24660), .O(n2_adj_3570)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_927 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n29741));
    defparam i1_2_lut_3_lut_adj_927.LUT_INIT = 16'he0e0;
    SB_LUT4 i12965_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n17352));
    defparam i12965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17198));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_928 (.I0(n54), .I1(n67), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n29733));
    defparam i1_2_lut_3_lut_adj_928.LUT_INIT = 16'he0e0;
    SB_LUT4 i17432_2_lut_4_lut (.I0(n1), .I1(n61), .I2(n133), .I3(\FRAME_MATCHER.state [30]), 
            .O(n21802));
    defparam i17432_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i16909_2_lut_4_lut (.I0(n1), .I1(n61), .I2(n133), .I3(\FRAME_MATCHER.state [29]), 
            .O(n21274));
    defparam i16909_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i17421_2_lut_4_lut (.I0(n1), .I1(n61), .I2(n133), .I3(\FRAME_MATCHER.state [14]), 
            .O(n21790));
    defparam i17421_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_929 (.I0(n1), .I1(n61), .I2(n133), .I3(\FRAME_MATCHER.state [11]), 
            .O(n29565));
    defparam i1_2_lut_4_lut_adj_929.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_930 (.I0(n1), .I1(n13117), .I2(n30199), 
            .I3(\FRAME_MATCHER.state [31]), .O(n29545));
    defparam i1_2_lut_4_lut_adj_930.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_931 (.I0(n1), .I1(n13117), .I2(n30199), 
            .I3(\FRAME_MATCHER.state [27]), .O(n29543));
    defparam i1_2_lut_4_lut_adj_931.LUT_INIT = 16'hea00;
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17197));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17196));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n17307));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_932 (.I0(n1), .I1(n13117), .I2(n30199), 
            .I3(\FRAME_MATCHER.state [23]), .O(n29541));
    defparam i1_2_lut_4_lut_adj_932.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_933 (.I0(n1), .I1(n13117), .I2(n30199), 
            .I3(\FRAME_MATCHER.state [15]), .O(n29539));
    defparam i1_2_lut_4_lut_adj_933.LUT_INIT = 16'hea00;
    SB_CARRY add_44_12 (.CI(n24660), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n24661));
    SB_LUT4 i12966_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n17353));
    defparam i12966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12967_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n17354));
    defparam i12967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12931_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n17318));
    defparam i12931_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17195));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12932_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n17319));
    defparam i12932_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17194));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12968_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n17355));
    defparam i12968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12969_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n17356));
    defparam i12969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12933_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n17320));
    defparam i12933_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12934_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n17321));
    defparam i12934_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12935_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n17322));
    defparam i12935_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12936_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n17323));
    defparam i12936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12970_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30176), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n17357));
    defparam i12970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12937_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n17324));
    defparam i12937_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12938_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30190), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n17325));
    defparam i12938_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_11_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n24659), .O(n2_adj_3571)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_11 (.CI(n24659), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n24660));
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1289));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_10_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n24658), .O(n2_adj_3572)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_934 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[6] [2]), .I3(n15671), .O(n10_adj_3573));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[6] [1]), .I1(n10_adj_3573), .I2(n30404), 
            .I3(GND_net), .O(n15772));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(n30631), .I1(n15772), .I2(n30221), .I3(n15587), 
            .O(n14_adj_3574));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n16139), .I1(n14_adj_3574), .I2(n10_adj_3575), 
            .I3(n16302), .O(Kp_23__N_1405));   // verilog/coms.v(69[16:27])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_44_10 (.CI(n24658), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n24659));
    SB_LUT4 add_44_9_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n24657), .O(n2_adj_3576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n15264), .I2(GND_net), 
            .I3(GND_net), .O(n15224));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_44_9 (.CI(n24657), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n24658));
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17193));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n10_adj_3577));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_44_8_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n24656), .O(n2_adj_3578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n17306));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_935 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_962));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_CARRY add_44_8 (.CI(n24656), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n24657));
    SB_LUT4 i3_2_lut (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3579));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_44_7_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n24655), .O(n2_adj_3580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_7 (.CI(n24655), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n24656));
    SB_LUT4 add_44_6_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n24654), .O(n2_adj_3581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_6 (.CI(n24654), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n24655));
    SB_LUT4 i12947_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n17334));
    defparam i12947_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12948_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n17335));
    defparam i12948_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12949_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n17336));
    defparam i12949_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_936 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15824));
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_5_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n24653), .O(n2_adj_3582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_5 (.CI(n24653), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n24654));
    SB_LUT4 i12950_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n17337));
    defparam i12950_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12951_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n17338));
    defparam i12951_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_44_4_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n24652), .O(n2_adj_3583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17192));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_619_9_lut (.I0(n11438), .I1(byte_transmit_counter[7]), .I2(GND_net), 
            .I3(n24688), .O(n34257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_619_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n24687), .O(n2236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12952_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n17339));
    defparam i12952_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_619_8 (.CI(n24687), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n24688));
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17191));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_619_7_lut (.I0(n11438), .I1(byte_transmit_counter[5]), .I2(GND_net), 
            .I3(n24686), .O(n34256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12953_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n17340));
    defparam i12953_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i9_4_lut (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [28]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [21]), 
            .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_619_7 (.CI(n24686), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n24687));
    SB_CARRY add_44_3 (.CI(n24651), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n24652));
    SB_LUT4 add_619_6_lut (.I0(n11438), .I1(byte_transmit_counter[4]), .I2(GND_net), 
            .I3(n24685), .O(n34258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_706_i1_4_lut (.I0(n21292), .I1(n22052), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n22062));   // verilog/coms.v(147[4] 288[11])
    defparam mux_706_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_adj_937.LUT_INIT = 16'heeee;
    SB_LUT4 i28825_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n22062), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n34460), .O(n34462));   // verilog/coms.v(147[4] 288[11])
    defparam i28825_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i1_4_lut (.I0(n47), .I1(n22054), .I2(n4_c), .I3(n50), .O(n3915));
    defparam i1_4_lut.LUT_INIT = 16'h3032;
    SB_LUT4 i26883_4_lut (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[0] [3]), .O(n32519));
    defparam i26883_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [2]), .O(n38));
    defparam i14_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [6]), .O(n39));
    defparam i15_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [6]), .O(n37));
    defparam i13_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i26879_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [2]), .O(n32515));
    defparam i26879_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_619_6 (.CI(n24685), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n24686));
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n32519), .O(n46));
    defparam i22_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i26881_4_lut (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [2]), .O(n32517));
    defparam i26881_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_3_lut (.I0(n32517), .I1(n46), .I2(n32515), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2428 [3]));
    defparam i23_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2230_3_lut (.I0(n3915), .I1(\FRAME_MATCHER.state [1]), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(GND_net), .O(n5784));
    defparam i2230_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i2_3_lut (.I0(n5784), .I1(\FRAME_MATCHER.state_31__N_2428 [3]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n12917));
    defparam i2_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i12954_3_lut_4_lut (.I0(n10_adj_3550), .I1(n31262), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n17341));
    defparam i12954_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_619_5_lut (.I0(n11438), .I1(byte_transmit_counter[3]), .I2(GND_net), 
            .I3(n24684), .O(n34255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_938 (.I0(n30266), .I1(n30675), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3584));
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_939 (.I0(n27227), .I1(n27225), .I2(n30504), .I3(n6_adj_3584), 
            .O(n26717));
    defparam i4_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16149));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_CARRY add_619_5 (.CI(n24684), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n24685));
    SB_LUT4 i1_4_lut_adj_941 (.I0(\data_in_frame[14] [0]), .I1(n26948), 
            .I2(\data_in_frame[13] [6]), .I3(\data_in_frame[13] [7]), .O(n30504));
    defparam i1_4_lut_adj_941.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_942 (.I0(\data_in_frame[18] [2]), .I1(n30504), 
            .I2(n30672), .I3(n15636), .O(n30591));
    defparam i1_4_lut_adj_942.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_943 (.I0(\data_in_frame[11] [4]), .I1(n16255), 
            .I2(n16360), .I3(n6_adj_3585), .O(n30266));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_944 (.I0(n31605), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30707));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut (.I0(Kp_23__N_1280), .I1(n27261), .I2(\data_in_frame[16] [5]), 
            .I3(\data_in_frame[18] [5]), .O(n30491));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_945 (.I0(n27248), .I1(n30266), .I2(n27225), .I3(n27227), 
            .O(n26635));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_945.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut (.I0(n30591), .I1(\data_in_frame[18] [4]), .I2(n30341), 
            .I3(\data_in_frame[15] [5]), .O(n22_adj_3586));
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut (.I0(n30510), .I1(\data_in_frame[18] [1]), .I2(\data_in_frame[17] [6]), 
            .I3(n15824), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_946 (.I0(n30491), .I1(\data_in_frame[17] [1]), 
            .I2(\data_in_frame[17] [7]), .I3(n30707), .O(n23));
    defparam i9_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n25), .I1(n15982), .I2(n23), .I3(n24), 
            .O(n30660));
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_948 (.I0(\data_in_frame[18] [0]), .I1(n30660), 
            .I2(n26635), .I3(GND_net), .O(n30483));
    defparam i2_3_lut_adj_948.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n13));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_949 (.I0(n30507), .I1(Kp_23__N_1405), .I2(\data_in_frame[15] [3]), 
            .I3(n30483), .O(n15));
    defparam i6_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_950 (.I0(\data_in_frame[19] [7]), .I1(n15), .I2(n13), 
            .I3(n14_adj_3587), .O(n30494));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_951 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10] [5]), 
            .I2(\data_in_frame[13] [0]), .I3(GND_net), .O(n30678));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_951.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_952 (.I0(Kp_23__N_962), .I1(n30235), .I2(\data_in_frame[5] [6]), 
            .I3(GND_net), .O(n30542));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_952.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_953 (.I0(n30678), .I1(\data_in_frame[13] [1]), 
            .I2(n30539), .I3(n30420), .O(n14_adj_3588));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_954 (.I0(n30740), .I1(n14_adj_3588), .I2(n10_adj_3589), 
            .I3(\data_in_frame[15] [2]), .O(n16321));   // verilog/coms.v(72[16:43])
    defparam i7_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30510));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_2_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n2_adj_3533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut (.I0(n26401), .I1(\data_in_frame[11] [7]), .I2(n30648), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_956 (.I0(\data_in_frame[14] [1]), .I1(n16262), 
            .I2(n8), .I3(n30469), .O(n30675));
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_957 (.I0(n30600), .I1(n30675), .I2(GND_net), 
            .I3(GND_net), .O(n27234));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_958 (.I0(n32089), .I1(n32127), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1280));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_959 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n15894), .I3(GND_net), .O(n30648));
    defparam i2_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_960 (.I0(n27227), .I1(Kp_23__N_829), .I2(n30498), 
            .I3(n6_adj_3590), .O(n26948));
    defparam i4_4_lut_adj_960.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_961 (.I0(Kp_23__N_1280), .I1(\data_in_frame[18] [1]), 
            .I2(n27234), .I3(Kp_23__N_1498), .O(n30737));
    defparam i3_4_lut_adj_961.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_962 (.I0(n26948), .I1(n30722), .I2(GND_net), 
            .I3(GND_net), .O(n30651));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_963 (.I0(n30725), .I1(\data_in_frame[11] [3]), 
            .I2(n16360), .I3(n16_adj_3591), .O(n15_adj_3592));
    defparam i6_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_964 (.I0(n15_adj_3592), .I1(\data_in_frame[8] [7]), 
            .I2(n14_adj_3593), .I3(n27225), .O(n27248));
    defparam i8_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_965 (.I0(n30212), .I1(n16139), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n14_adj_3594));   // verilog/coms.v(71[16:42])
    defparam i5_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_966 (.I0(n30263), .I1(n30554), .I2(\data_in_frame[11] [0]), 
            .I3(\data_in_frame[8] [6]), .O(n15_adj_3595));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_967 (.I0(n15_adj_3595), .I1(\data_in_frame[8] [7]), 
            .I2(n14_adj_3594), .I3(\data_in_frame[6] [2]), .O(n15790));   // verilog/coms.v(71[16:42])
    defparam i8_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30554));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_969 (.I0(n15573), .I1(\data_in_frame[6] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n16255));   // verilog/coms.v(77[16:35])
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_970 (.I0(n30480), .I1(\data_in_frame[7] [3]), .I2(\data_in_frame[11] [5]), 
            .I3(n27227), .O(n10_adj_3596));
    defparam i4_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_971 (.I0(\data_in_frame[13] [7]), .I1(n26712), 
            .I2(GND_net), .I3(GND_net), .O(n30469));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_972 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n30235));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_972.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_973 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n14_adj_3597));   // verilog/coms.v(230[9:81])
    defparam i5_3_lut_adj_973.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_974 (.I0(n30235), .I1(\data_in_frame[12] [5]), 
            .I2(n15697), .I3(n15671), .O(n15_adj_3598));   // verilog/coms.v(230[9:81])
    defparam i6_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_975 (.I0(n15_adj_3598), .I1(\data_in_frame[6] [2]), 
            .I2(n14_adj_3597), .I3(\data_in_frame[7] [7]), .O(n15604));   // verilog/coms.v(230[9:81])
    defparam i8_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_976 (.I0(\data_in_frame[15] [3]), .I1(n15604), 
            .I2(GND_net), .I3(GND_net), .O(n30606));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_977 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30397));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_977.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_978 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[9] [2]), .I3(GND_net), .O(n30790));
    defparam i2_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30740));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_980 (.I0(n15746), .I1(\data_in_frame[8] [4]), .I2(\data_in_frame[10] [5]), 
            .I3(n30740), .O(n10_adj_3599));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_981 (.I0(\data_in_frame[6] [3]), .I1(n10_adj_3599), 
            .I2(\data_in_frame[15] [0]), .I3(GND_net), .O(n30232));   // verilog/coms.v(70[16:41])
    defparam i5_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_14__7__I_0_3249_2_lut (.I0(\data_in_frame[14] [7]), 
            .I1(\data_in_frame[14] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1327));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_14__7__I_0_3249_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_982 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[10] [1]), 
            .I2(n30710), .I3(n30758), .O(n30291));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1126_i7_2_lut (.I0(Kp_23__N_962), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3600));   // verilog/coms.v(230[9:81])
    defparam equal_1126_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_983 (.I0(\data_in_frame[14] [4]), .I1(n30704), 
            .I2(n16098), .I3(n30784), .O(n16_adj_3601));
    defparam i6_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_984 (.I0(n30356), .I1(n30758), .I2(\data_in_frame[12] [3]), 
            .I3(n30628), .O(n17_adj_3602));
    defparam i7_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_985 (.I0(n17_adj_3602), .I1(\data_in_frame[7] [4]), 
            .I2(n16_adj_3601), .I3(\data_in_frame[10] [0]), .O(n32127));
    defparam i9_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n15525));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n24651));
    SB_LUT4 i2_3_lut_adj_987 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n30356));
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_988 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[1] [5]), .O(n30404));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_989 (.I0(n30393), .I1(n30575), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n30704));
    defparam i2_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_in_frame[5] [7]), .I1(n30404), .I2(GND_net), 
            .I3(GND_net), .O(n16098));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_991 (.I0(n15894), .I1(\data_in_frame[12] [3]), 
            .I2(n4_adj_3603), .I3(\data_in_frame[14] [5]), .O(n8_adj_3604));
    defparam i1_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30628));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1019));   // verilog/coms.v(83[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(Kp_23__N_1019), .I1(n30628), .I2(\data_in_frame[7] [5]), 
            .I3(\data_in_frame[10] [1]), .O(n12_adj_3605));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[6] [0]), .I1(n12_adj_3605), .I2(n8_adj_3604), 
            .I3(GND_net), .O(n30519));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut (.I0(n30212), .I1(n16094), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_3606));   // verilog/coms.v(83[17:28])
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_993 (.I0(n30356), .I1(\data_in_frame[8] [2]), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[6] [1]), .O(n14_adj_3607));   // verilog/coms.v(83[17:28])
    defparam i6_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_994 (.I0(\data_in_frame[12] [4]), .I1(n14_adj_3607), 
            .I2(n10_adj_3606), .I3(Kp_23__N_1019), .O(n15704));   // verilog/coms.v(83[17:28])
    defparam i7_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_995 (.I0(\data_in_frame[3] [7]), .I1(n30455), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[4] [1]), .O(n15671));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_996 (.I0(n15671), .I1(\data_in_frame[8] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n30263));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_997 (.I0(n15557), .I1(\data_in_frame[0] [0]), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[4] [2]), .O(n15746));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_998 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15587));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_999 (.I0(\data_in_frame[4] [3]), .I1(n30205), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[2] [1]), .O(n16067));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1000 (.I0(n16067), .I1(n30221), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(n15753));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1000.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1001 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[8] [7]), 
            .I2(n15753), .I3(GND_net), .O(n30631));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1001.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1002 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[6] [6]), .I3(GND_net), .O(n14_adj_3608));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_1002.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1003 (.I0(Kp_23__N_829), .I1(n30420), .I2(\data_in_frame[6] [7]), 
            .I3(\data_in_frame[9] [1]), .O(n15_adj_3609));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1004 (.I0(n15_adj_3609), .I1(\data_in_frame[4] [6]), 
            .I2(n14_adj_3608), .I3(\data_in_frame[9] [0]), .O(n15781));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1005 (.I0(n15781), .I1(n30725), .I2(n30631), 
            .I3(n30414), .O(n16146));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(n16146), .I1(n30340), .I2(GND_net), 
            .I3(GND_net), .O(n30341));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(n27165), .I1(\data_in_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27276));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(n15704), .I1(n30519), .I2(GND_net), 
            .I3(GND_net), .O(n26563));
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1009 (.I0(n26388), .I1(n30666), .I2(\data_in_frame[9] [3]), 
            .I3(n10_adj_3596), .O(n26712));
    defparam i5_3_lut_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1010 (.I0(\data_in_frame[16] [1]), .I1(n15982), 
            .I2(\data_in_frame[16] [3]), .I3(\data_in_frame[16] [5]), .O(Kp_23__N_1498));   // verilog/coms.v(83[17:63])
    defparam i3_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1126_i16_2_lut (.I0(Kp_23__N_832), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3591));   // verilog/coms.v(230[9:81])
    defparam equal_1126_i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(n30393), .I1(\data_in_frame[5] [1]), 
            .I2(n26493), .I3(GND_net), .O(n27227));
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n30288), .I1(n30575), .I2(\data_in_frame[5] [4]), 
            .I3(GND_net), .O(n16094));
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(n16094), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30452));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15844));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[1] [3]), .I1(n30288), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3610));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1016 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [2]), .I3(n6_adj_3610), .O(n15697));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\data_in_frame[11] [7]), .I1(n15697), 
            .I2(GND_net), .I3(GND_net), .O(n30609));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1018 (.I0(n15844), .I1(n30452), .I2(n30368), 
            .I3(\data_in_frame[9] [6]), .O(n26401));
    defparam i3_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\data_in_frame[5] [2]), .I1(n16208), 
            .I2(GND_net), .I3(GND_net), .O(n30784));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15557));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1021 (.I0(\data_in_frame[15] [4]), .I1(n15790), 
            .I2(n16146), .I3(GND_net), .O(n15994));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1022 (.I0(\data_in_frame[15] [4]), .I1(n15790), 
            .I2(\data_in_frame[13] [5]), .I3(n27276), .O(n14_adj_3587));   // verilog/coms.v(73[16:43])
    defparam i5_3_lut_4_lut_adj_1022.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1023 (.I0(n15677), .I1(\data_in_frame[2] [6]), 
            .I2(n15557), .I3(\data_in_frame[2] [7]), .O(n14_adj_3611));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1024 (.I0(\data_in_frame[3] [2]), .I1(n14_adj_3611), 
            .I2(n10_adj_3577), .I3(Kp_23__N_823), .O(n30536));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30455));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15725));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i12514_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n16901));
    defparam i12514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12828_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n17215));
    defparam i12828_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1027 (.I0(n15725), .I1(n30455), .I2(n30429), 
            .I3(\data_in_frame[1] [3]), .O(Kp_23__N_794));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1028 (.I0(Kp_23__N_794), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3612));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1029 (.I0(n7_adj_3612), .I1(\data_in_frame[2] [6]), 
            .I2(n30545), .I3(\data_in_frame[0] [4]), .O(n16208));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1030 (.I0(n30536), .I1(\data_in_frame[0] [1]), 
            .I2(Kp_23__N_829), .I3(n30353), .O(n12));   // verilog/coms.v(76[16:27])
    defparam i5_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(n26493), .I1(n16208), .I2(GND_net), 
            .I3(GND_net), .O(n27175));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1032 (.I0(n30536), .I1(n7_adj_3612), .I2(\data_in_frame[2] [4]), 
            .I3(n30545), .O(n10_adj_3569));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1033 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[7] [2]), .I3(GND_net), .O(n30498));
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n16114), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[2] [5]), .O(Kp_23__N_829));   // verilog/coms.v(74[16:43])
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[5] [0]), .I1(n30368), 
            .I2(GND_net), .I3(GND_net), .O(n26388));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1036 (.I0(Kp_23__N_829), .I1(\data_in_frame[14] [2]), 
            .I2(n30498), .I3(GND_net), .O(n14_adj_3613));
    defparam i5_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1037 (.I0(\data_in_frame[11] [7]), .I1(n30666), 
            .I2(Kp_23__N_832), .I3(\data_in_frame[7] [3]), .O(n15_adj_3614));
    defparam i6_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1038 (.I0(n15_adj_3614), .I1(\data_in_frame[4] [7]), 
            .I2(n14_adj_3613), .I3(n26388), .O(n30336));
    defparam i8_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17190));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17189));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1039 (.I0(\data_in_frame[9] [7]), .I1(n16262), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[12] [1]), .O(n30710));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17188));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17187));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17186));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1040 (.I0(n30710), .I1(n30336), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3615));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1041 (.I0(n26401), .I1(n30609), .I2(n30374), 
            .I3(n6_adj_3615), .O(n30600));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3616));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1043 (.I0(n30368), .I1(n30291), .I2(n30609), 
            .I3(n6_adj_3616), .O(n32089));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1044 (.I0(\data_in_frame[16] [0]), .I1(n30426), 
            .I2(Kp_23__N_1498), .I3(n26563), .O(n31605));
    defparam i3_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(n32089), .I1(n30600), .I2(GND_net), 
            .I3(GND_net), .O(n30601));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30353));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17185));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17184));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30205));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1048 (.I0(n30205), .I1(n4_adj_3617), .I2(\data_in_frame[0] [0]), 
            .I3(GND_net), .O(Kp_23__N_823));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1049 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_adj_3617));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1049.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(\data_in_frame[4] [5]), .I1(n16114), 
            .I2(n4_adj_3617), .I3(GND_net), .O(n15573));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(Kp_23__N_823), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16302));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30429));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15677));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_DFFSR tx_transmit_3227 (.Q(\r_SM_Main_2__N_3259[0] ), .C(clk32MHz), 
            .D(n34462), .R(n30807));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17183));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1054 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(n16360), .I3(GND_net), .O(n16139));
    defparam i2_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_LUT4 i11_3_lut (.I0(byte_transmit_counter[2]), .I1(n34331), .I2(n16491), 
            .I3(GND_net), .O(n29349));   // verilog/coms.v(100[12:33])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14056_3_lut (.I0(byte_transmit_counter[3]), .I1(n34255), .I2(n16491), 
            .I3(GND_net), .O(n17517));
    defparam i14056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14062_3_lut (.I0(byte_transmit_counter[4]), .I1(n34258), .I2(n16491), 
            .I3(GND_net), .O(n17518));
    defparam i14062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14058_3_lut (.I0(byte_transmit_counter[5]), .I1(n34256), .I2(n16491), 
            .I3(GND_net), .O(n17519));
    defparam i14058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7187_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n11438));
    defparam i7187_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_1126_i15_2_lut (.I0(Kp_23__N_829), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3618));   // verilog/coms.v(230[9:81])
    defparam equal_1126_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(n27227), .I1(n15_adj_3618), .I2(n30368), .I3(n15697), 
            .O(n28));   // verilog/coms.v(230[9:81])
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i10_4_lut_adj_1055 (.I0(n15573), .I1(n16302), .I2(n16067), 
            .I3(n15894), .O(n26));   // verilog/coms.v(230[9:81])
    defparam i10_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n16094), .I1(n30212), .I2(n16_adj_3591), .I3(n27225), 
            .O(n27));   // verilog/coms.v(230[9:81])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1056 (.I0(n15746), .I1(n7_adj_3600), .I2(n15671), 
            .I3(n16098), .O(n25_adj_3619));   // verilog/coms.v(230[9:81])
    defparam i9_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1057 (.I0(n25_adj_3619), .I1(n27), .I2(n26), 
            .I3(n28), .O(n31_c));   // verilog/coms.v(230[9:81])
    defparam i15_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(n30093), .I1(n30201), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3620));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1059 (.I0(n234), .I1(n30203), .I2(n63_adj_3621), 
            .I3(n6_adj_3620), .O(n22054));
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1060 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(n30793), .O(n30254));
    defparam i1_2_lut_3_lut_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i15_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));
    defparam i15_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(n16139), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30414));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1062 (.I0(\data_in_frame[10] [7]), .I1(n30212), 
            .I2(\data_in_frame[11] [0]), .I3(GND_net), .O(n30539));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1062.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(\data_in_frame[14] [3]), .I1(n26563), .I2(\data_in_frame[14] [4]), 
            .I3(n34), .O(n58));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n30374), .I1(n30232), .I2(n30336), .I3(\data_in_frame[7] [1]), 
            .O(n56_adj_3622));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n27175), .I1(\data_in_frame[8] [6]), .I2(\data_in_frame[11] [2]), 
            .I3(\data_in_frame[12] [4]), .O(n57));
    defparam i24_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut_adj_1063 (.I0(n30722), .I1(n30458), .I2(n30539), 
            .I3(n30414), .O(n55));
    defparam i22_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(\data_in_frame[15] [4]), .I1(n30790), .I2(\data_in_frame[13] [0]), 
            .I3(n15636), .O(n52));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[6] [4]), .I3(n30778), .O(n54_adj_3623));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n30452), .I1(\data_in_frame[14] [1]), .I2(n30359), 
            .I3(\data_in_frame[8] [5]), .O(n53));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n55), .I1(n57), .I2(n56_adj_3622), .I3(n58), 
            .O(n64));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n30528), .I1(n52), .I2(n8_adj_3604), .I3(n26388), 
            .O(n59));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(n59), .I1(n64), .I2(n53), .I3(n54_adj_3623), 
            .O(n27165));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1064 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3624));
    defparam i6_4_lut_adj_1064.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_1065 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [4]), .O(n14_adj_3625));   // verilog/coms.v(232[13:35])
    defparam i6_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 add_619_4_lut (.I0(n11438), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(n24683), .O(n34331)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1066 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3626));
    defparam i5_4_lut_adj_1066.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1067 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3627));   // verilog/coms.v(232[13:35])
    defparam i5_4_lut_adj_1067.LUT_INIT = 16'hfffe;
    SB_LUT4 i16918_4_lut (.I0(n13_adj_3627), .I1(n13_adj_3626), .I2(n14_adj_3625), 
            .I3(n14_adj_3624), .O(n21283));
    defparam i16918_4_lut.LUT_INIT = 16'h32fa;
    SB_CARRY add_619_4 (.CI(n24683), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n24684));
    SB_LUT4 i6_4_lut_adj_1068 (.I0(\data_in_frame[15] [7]), .I1(n15994), 
            .I2(n30663), .I3(n30340), .O(n16_adj_3628));
    defparam i6_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1069 (.I0(\data_in_frame[18] [0]), .I1(n30651), 
            .I2(n30737), .I3(\data_in_frame[15] [6]), .O(n17_adj_3629));
    defparam i7_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1070 (.I0(n30494), .I1(n30663), .I2(\data_in_frame[20] [0]), 
            .I3(n30483), .O(n12_adj_3630));
    defparam i5_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1071 (.I0(n27171), .I1(n30660), .I2(n30494), 
            .I3(\data_in_frame[20] [1]), .O(n31718));
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1072 (.I0(\data_in_frame[18] [4]), .I1(n30326), 
            .I2(\data_in_frame[20] [5]), .I3(n27261), .O(n31188));
    defparam i3_4_lut_adj_1072.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1073 (.I0(\data_in_frame[21] [2]), .I1(n26767), 
            .I2(Kp_23__N_1289), .I3(n26452), .O(n31425));
    defparam i3_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1074 (.I0(\data_in_frame[20] [4]), .I1(n30591), 
            .I2(n30326), .I3(\data_in_frame[16] [2]), .O(n31345));
    defparam i3_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1075 (.I0(n30491), .I1(\data_in_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3631));
    defparam i2_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1076 (.I0(n30778), .I1(n27171), .I2(n30672), 
            .I3(n26712), .O(n14_adj_3632));
    defparam i6_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[18] [7]), .I1(n26930), .I2(n26767), 
            .I3(GND_net), .O(n5_adj_3633));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1077 (.I0(\data_in_frame[20] [3]), .I1(n30737), 
            .I2(n30397), .I3(\data_in_frame[18] [2]), .O(n13_adj_3634));
    defparam i5_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(n30601), .I1(n15525), .I2(n26717), 
            .I3(\data_in_frame[18] [4]), .O(n10_adj_3635));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1079 (.I0(\data_in_frame[20] [6]), .I1(n10_adj_3635), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n31451));
    defparam i5_3_lut_adj_1079.LUT_INIT = 16'h9696;
    SB_LUT4 i26845_4_lut (.I0(n13_adj_3634), .I1(n5_adj_3633), .I2(n14_adj_3632), 
            .I3(n6_adj_3631), .O(n32479));
    defparam i26845_4_lut.LUT_INIT = 16'h1248;
    SB_LUT4 i12829_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n17216));
    defparam i12829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1080 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[15] [0]), .I3(GND_net), .O(n14_adj_3636));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i12830_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n17217));
    defparam i12830_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1081 (.I0(n30603), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[17] [2]), .I3(n30359), .O(n15_adj_3637));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1082 (.I0(n17_adj_3629), .I1(n26717), .I2(n16_adj_3628), 
            .I3(\data_in_frame[20] [2]), .O(n31682));
    defparam i9_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1083 (.I0(\data_in_frame[19] [3]), .I1(n30329), 
            .I2(\data_in_frame[21] [4]), .I3(n26405), .O(n31191));
    defparam i3_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1084 (.I0(n15_adj_3637), .I1(n15790), .I2(n14_adj_3636), 
            .I3(\data_in_frame[19] [5]), .O(n31442));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1085 (.I0(\data_in_frame[21] [3]), .I1(n26452), 
            .I2(n30329), .I3(GND_net), .O(n30595));
    defparam i1_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[21] [5]), .I1(n11), .I2(n30474), 
            .I3(n12_adj_3630), .O(n18_adj_3638));
    defparam i2_4_lut.LUT_INIT = 16'hde7b;
    SB_LUT4 i2_4_lut_adj_1086 (.I0(Kp_23__N_1289), .I1(n26930), .I2(\data_in_frame[21] [0]), 
            .I3(n26767), .O(n31180));
    defparam i2_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i26889_4_lut (.I0(n31345), .I1(n31425), .I2(n31188), .I3(n31718), 
            .O(n32525));
    defparam i26889_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_1087 (.I0(n32479), .I1(\data_in_frame[21] [1]), 
            .I2(n31451), .I3(n26930), .O(n26_adj_3639));
    defparam i10_4_lut_adj_1087.LUT_INIT = 16'hfdf7;
    SB_LUT4 i11_4_lut_adj_1088 (.I0(n30595), .I1(n31442), .I2(n31191), 
            .I3(n31682), .O(n27_adj_3640));
    defparam i11_4_lut_adj_1088.LUT_INIT = 16'hfbff;
    SB_LUT4 i9_4_lut_adj_1089 (.I0(n31180), .I1(n18_adj_3638), .I2(\data_in_frame[21] [7]), 
            .I3(n30516), .O(n25_adj_3641));
    defparam i9_4_lut_adj_1089.LUT_INIT = 16'hfeef;
    SB_LUT4 i15_4_lut_adj_1090 (.I0(n25_adj_3641), .I1(n27_adj_3640), .I2(n26_adj_3639), 
            .I3(n32525), .O(n31_adj_3642));
    defparam i15_4_lut_adj_1090.LUT_INIT = 16'hfeff;
    SB_LUT4 add_619_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n24682), .O(n2236[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16927_2_lut (.I0(n31_adj_3642), .I1(n21283), .I2(GND_net), 
            .I3(GND_net), .O(n21292));
    defparam i16927_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14121_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n21292), .O(n18507));   // verilog/coms.v(110[11:16])
    defparam i14121_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i2_4_lut_adj_1091 (.I0(n12846), .I1(n22054), .I2(n18507), 
            .I3(n4311), .O(n16491));
    defparam i2_4_lut_adj_1091.LUT_INIT = 16'h2220;
    SB_LUT4 i12831_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n17218));
    defparam i12831_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14060_3_lut (.I0(byte_transmit_counter[7]), .I1(n34257), .I2(n16491), 
            .I3(GND_net), .O(n17521));
    defparam i14060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12832_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n17219));
    defparam i12832_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_619_3 (.CI(n24682), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n24683));
    SB_LUT4 i12833_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n17220));
    defparam i12833_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_619_2_lut (.I0(n11438), .I1(byte_transmit_counter[0]), .I2(tx_transmit_N_3151), 
            .I3(GND_net), .O(n34330)) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_619_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3151), 
            .CO(n24682));
    SB_LUT4 i12834_3_lut_4_lut (.I0(n10), .I1(n30180), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n17221));
    defparam i12834_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12899_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n17286));
    defparam i12899_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_33_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n24681), .O(n2_adj_3643)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_32_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n24680), .O(n2_adj_3644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12900_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n17287));
    defparam i12900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_32 (.CI(n24680), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n24681));
    SB_LUT4 add_44_31_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n24679), .O(n2_adj_3645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12901_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n17288));
    defparam i12901_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_31 (.CI(n24679), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n24680));
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17182));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17181));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_30_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n24678), .O(n2_adj_3646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12902_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n17289));
    defparam i12902_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17180));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17179));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17176));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17175));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17174));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17173));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17172));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17171));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17170));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_1092 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[17] [2]), 
            .I2(n30519), .I3(n6_adj_3647), .O(n26405));
    defparam i4_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17167));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17166));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_30 (.CI(n24678), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n24679));
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17163));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17153));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17152));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17150));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n15369));   // verilog/coms.v(253[5:27])
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17148));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3648), .S(n3_adj_3561));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17147));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_330_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_330_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1094 (.I0(n5_adj_3649), .I1(\data_in[3] [2]), .I2(\data_in[3] [7]), 
            .I3(\data_in[0] [1]), .O(n10_adj_3650));
    defparam i2_4_lut_adj_1094.LUT_INIT = 16'hffef;
    SB_LUT4 i6_4_lut_adj_1095 (.I0(\data_in[2] [0]), .I1(\data_in[1] [2]), 
            .I2(\data_in[1] [6]), .I3(\data_in[0] [5]), .O(n14_adj_3651));
    defparam i6_4_lut_adj_1095.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1096 (.I0(\data_in[2] [5]), .I1(n14_adj_3651), 
            .I2(n10_adj_3650), .I3(\data_in[2] [6]), .O(n15283));
    defparam i7_4_lut_adj_1096.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1097 (.I0(n15283), .I1(\data_in[0] [7]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_3652));
    defparam i6_4_lut_adj_1097.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37044));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37044_bdd_4_lut (.I0(n37044), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37047));
    defparam n37044_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31378 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37038));
    defparam byte_transmit_counter_0__bdd_4_lut_31378.LUT_INIT = 16'he4aa;
    SB_LUT4 n37038_bdd_4_lut (.I0(n37038), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37041));
    defparam n37038_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1098 (.I0(n15355), .I1(\data_in[0] [2]), .I2(\data_in[3] [3]), 
            .I3(\data_in[3] [1]), .O(n17_adj_3653));
    defparam i7_4_lut_adj_1098.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1099 (.I0(n17_adj_3653), .I1(\data_in[2] [3]), 
            .I2(n16_adj_3652), .I3(\data_in[3] [5]), .O(n63_adj_3554));
    defparam i9_4_lut_adj_1099.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1100 (.I0(\data_in[3] [0]), .I1(n15427), .I2(n15283), 
            .I3(\data_in[2] [2]), .O(n16_adj_3654));
    defparam i6_4_lut_adj_1100.LUT_INIT = 16'hfffe;
    SB_LUT4 i12903_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n17290));
    defparam i12903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1101 (.I0(\data_in[2] [4]), .I1(\data_in[1] [0]), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n17_adj_3655));
    defparam i7_4_lut_adj_1101.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1102 (.I0(n17_adj_3655), .I1(\data_in[0] [6]), 
            .I2(n16_adj_3654), .I3(\data_in[1] [4]), .O(n63_adj_3553));
    defparam i9_4_lut_adj_1102.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_3_lut (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i17023_4_lut (.I0(n10_adj_3656), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n15421), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i17023_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n32541), .I2(n32542), .I3(byte_transmit_counter[2]), .O(n37026));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 add_44_29_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n24677), .O(n2_adj_3657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n37026_bdd_4_lut (.I0(n37026), .I1(n32545), .I2(n32544), .I3(byte_transmit_counter[2]), 
            .O(n37029));
    defparam n37026_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31364 (.I0(byte_transmit_counter[1]), 
            .I1(n32550), .I2(n32551), .I3(byte_transmit_counter[2]), .O(n37020));
    defparam byte_transmit_counter_1__bdd_4_lut_31364.LUT_INIT = 16'he4aa;
    SB_LUT4 n37020_bdd_4_lut (.I0(n37020), .I1(n32548), .I2(n32547), .I3(byte_transmit_counter[2]), 
            .O(n37023));
    defparam n37020_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31373 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37014));
    defparam byte_transmit_counter_0__bdd_4_lut_31373.LUT_INIT = 16'he4aa;
    SB_LUT4 n37014_bdd_4_lut (.I0(n37014), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37017));
    defparam n37014_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31359 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3549), .I2(n34278), .I3(byte_transmit_counter[2]), 
            .O(n37008));
    defparam byte_transmit_counter_1__bdd_4_lut_31359.LUT_INIT = 16'he4aa;
    SB_LUT4 i27007_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n32644));
    defparam i27007_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12904_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n17291));
    defparam i12904_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(byte_transmit_counter[7]), .I1(n21899), 
            .I2(byte_transmit_counter[6]), .I3(byte_transmit_counter[5]), 
            .O(n22044));
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(n15239), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3658));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'heeee;
    SB_LUT4 i17019_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3658), .I3(\FRAME_MATCHER.i [1]), .O(n740));   // verilog/coms.v(157[9:60])
    defparam i17019_4_lut.LUT_INIT = 16'h3230;
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17146));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17145));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n37008_bdd_4_lut (.I0(n37008), .I1(n17_adj_3547), .I2(n16_adj_3546), 
            .I3(byte_transmit_counter[2]), .O(n37011));
    defparam n37008_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31354 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n36996));
    defparam byte_transmit_counter_0__bdd_4_lut_31354.LUT_INIT = 16'he4aa;
    SB_LUT4 n36996_bdd_4_lut (.I0(n36996), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n36999));
    defparam n36996_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17143));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17142));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17139));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17138));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17137));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17136));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17135));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_29 (.CI(n24677), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n24678));
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17133));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31349 (.I0(byte_transmit_counter[1]), 
            .I1(n34176), .I2(n5_c), .I3(byte_transmit_counter[2]), .O(n36984));
    defparam byte_transmit_counter_1__bdd_4_lut_31349.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31329 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3543), .I2(n34175), .I3(byte_transmit_counter[2]), 
            .O(n36978));
    defparam byte_transmit_counter_1__bdd_4_lut_31329.LUT_INIT = 16'he4aa;
    SB_LUT4 n36978_bdd_4_lut (.I0(n36978), .I1(n17_adj_3542), .I2(n16_adj_3541), 
            .I3(byte_transmit_counter[2]), .O(n36981));
    defparam n36978_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_1105 (.I0(n15358), .I1(n21813), .I2(n15264), 
            .I3(GND_net), .O(n6_adj_3659));
    defparam i1_3_lut_adj_1105.LUT_INIT = 16'hc8c8;
    SB_LUT4 i4_4_lut_adj_1106 (.I0(n63_adj_3660), .I1(n15494), .I2(n15502), 
            .I3(n6_adj_3659), .O(n2421));
    defparam i4_4_lut_adj_1106.LUT_INIT = 16'h8000;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [19]), .O(n42));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17132));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i15_4_lut_adj_1107 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [27]), .I3(\FRAME_MATCHER.i [10]), .O(n40));
    defparam i15_4_lut_adj_1107.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [13]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1108 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(\FRAME_MATCHER.i [11]), .O(n39_adj_3661));
    defparam i14_4_lut_adj_1108.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38_adj_3662));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3663));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12905_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n17292));
    defparam i12905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12906_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30176), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n17293));
    defparam i12906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31324 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3540), .I2(n34172), .I3(byte_transmit_counter[2]), 
            .O(n36972));
    defparam byte_transmit_counter_1__bdd_4_lut_31324.LUT_INIT = 16'he4aa;
    SB_LUT4 n36972_bdd_4_lut (.I0(n36972), .I1(n17_adj_3539), .I2(n16_adj_3538), 
            .I3(byte_transmit_counter[2]), .O(n36975));
    defparam n36972_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31319 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3537), .I2(n34171), .I3(byte_transmit_counter[2]), 
            .O(n36966));
    defparam byte_transmit_counter_1__bdd_4_lut_31319.LUT_INIT = 16'he4aa;
    SB_LUT4 n36966_bdd_4_lut (.I0(n36966), .I1(n17), .I2(n16), .I3(byte_transmit_counter[2]), 
            .O(n36969));
    defparam n36966_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31314 (.I0(byte_transmit_counter[1]), 
            .I1(n19), .I2(n34170), .I3(byte_transmit_counter[2]), .O(n36960));
    defparam byte_transmit_counter_1__bdd_4_lut_31314.LUT_INIT = 16'he4aa;
    SB_LUT4 i23_4_lut_adj_1109 (.I0(n39_adj_3661), .I1(n41), .I2(n40), 
            .I3(n42), .O(n48));
    defparam i23_4_lut_adj_1109.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [23]), .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1110 (.I0(n43), .I1(n48), .I2(n37_adj_3663), 
            .I3(n38_adj_3662), .O(n15421));
    defparam i24_4_lut_adj_1110.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1111 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3664));
    defparam i4_4_lut_adj_1111.LUT_INIT = 16'hfdff;
    SB_LUT4 add_44_3_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n24651), .O(n2_adj_3648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_adj_1112 (.I0(\data_in[2] [7]), .I1(n10_adj_3664), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n15424));
    defparam i5_3_lut_adj_1112.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3665));
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'heeee;
    SB_LUT4 i26831_4_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(\data_in[1] [5]), 
            .I3(\data_in[2] [2]), .O(n32465));
    defparam i26831_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1114 (.I0(n32465), .I1(n7_adj_3665), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n15355));
    defparam i5_4_lut_adj_1114.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_2_lut_adj_1115 (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3666));
    defparam i2_2_lut_adj_1115.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3667));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(\data_in[3] [6]), .I1(n14_adj_3667), 
            .I2(n10_adj_3666), .I3(\data_in[2] [1]), .O(n15427));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_2_lut_adj_1118 (.I0(\data_in[1] [3]), .I1(\data_in[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3668));
    defparam i3_2_lut_adj_1118.LUT_INIT = 16'hdddd;
    SB_LUT4 i9_4_lut_adj_1119 (.I0(\data_in[3] [7]), .I1(n15427), .I2(\data_in[2] [6]), 
            .I3(\data_in[0] [5]), .O(n22_adj_3669));
    defparam i9_4_lut_adj_1119.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_3_lut_adj_1120 (.I0(\data_in[2] [5]), .I1(\data_in[1] [2]), 
            .I2(n15355), .I3(GND_net), .O(n20_adj_3670));
    defparam i7_3_lut_adj_1120.LUT_INIT = 16'hf7f7;
    SB_LUT4 i11_4_lut_adj_1121 (.I0(n15424), .I1(n22_adj_3669), .I2(n16_adj_3668), 
            .I3(\data_in[0] [1]), .O(n24_adj_3671));
    defparam i11_4_lut_adj_1121.LUT_INIT = 16'hfeff;
    SB_LUT4 i12_4_lut_adj_1122 (.I0(\data_in[2] [0]), .I1(n24_adj_3671), 
            .I2(n20_adj_3670), .I3(\data_in[3] [2]), .O(n63));
    defparam i12_4_lut_adj_1122.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut_adj_1123 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n15493), .I3(GND_net), .O(n15494));   // verilog/coms.v(195[5:24])
    defparam i2_3_lut_adj_1123.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_adj_1124 (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_3553), 
            .I2(n63_adj_3554), .I3(GND_net), .O(n18493));   // verilog/coms.v(110[11:16])
    defparam i1_3_lut_adj_1124.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_355_Select_2_i5_4_lut (.I0(n2857), .I1(n15504), .I2(n63), 
            .I3(n18493), .O(n5));
    defparam select_355_Select_2_i5_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i1_rep_134_2_lut (.I0(n63), .I1(n18493), .I2(GND_net), .I3(GND_net), 
            .O(n37539));   // verilog/coms.v(110[11:16])
    defparam i1_rep_134_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17131));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17130));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17129));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17127));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_28_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n24676), .O(n2_adj_3673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_28 (.CI(n24676), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n24677));
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17126));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12891_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n17278));
    defparam i12891_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21269), .O(n30187));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17124));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n36960_bdd_4_lut (.I0(n36960), .I1(n17_adj_3674), .I2(n16_adj_3675), 
            .I3(byte_transmit_counter[2]), .O(n36963));
    defparam n36960_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11_3_lut_adj_1125 (.I0(byte_transmit_counter[0]), .I1(n34330), 
            .I2(n16491), .I3(GND_net), .O(n29343));   // verilog/coms.v(100[12:33])
    defparam i11_3_lut_adj_1125.LUT_INIT = 16'hcaca;
    SB_LUT4 i17022_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15239), .I3(\FRAME_MATCHER.i [31]), .O(n2857));
    defparam i17022_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i2014_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3656));
    defparam i2014_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i12892_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n17279));
    defparam i12892_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1126 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21269), .O(n31262));
    defparam i2_2_lut_3_lut_4_lut_adj_1126.LUT_INIT = 16'h8000;
    SB_LUT4 add_44_27_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n24675), .O(n2_adj_3676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_27 (.CI(n24675), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n24676));
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17262));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12893_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n17280));
    defparam i12893_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12894_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n17281));
    defparam i12894_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_26_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n24674), .O(n2_adj_3677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_26 (.CI(n24674), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n24675));
    SB_LUT4 add_44_25_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n24673), .O(n2_adj_3678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_25 (.CI(n24673), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n24674));
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n17284));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n17283));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n17282));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n17281));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n17280));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17279));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17278));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17277));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17276));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3583), .S(n3_adj_3679));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3582), .S(n3_adj_3680));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3581), .S(n3_adj_3681));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3580), .S(n3_adj_3682));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3578), .S(n3_adj_3683));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3576), .S(n3_adj_3684));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3572), .S(n3_adj_3685));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3571), .S(n3_adj_3686));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3570), .S(n3_adj_3687));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3566), .S(n3_adj_3688));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3563), .S(n3_adj_3689));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3556), .S(n3_adj_3690));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3545), .S(n3_adj_3691));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3536), .S(n3_adj_3692));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3535), .S(n3_adj_3693));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3534), .S(n3_adj_3694));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3695));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3696), .S(n3_adj_3697));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3698), .S(n3_adj_3699));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3700), .S(n3_adj_3701));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3702), .S(n3_adj_3703));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3678), .S(n3_adj_3704));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3677), .S(n3_adj_3705));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3676), .S(n3_adj_3706));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3673), .S(n3_adj_3707));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3657), .S(n3_adj_3708));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3646), .S(n3_adj_3709));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3645), .S(n3_adj_3710));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3644), .S(n3_adj_3711));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3643), .S(n3_adj_3712));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17122));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17121));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17120));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n16553), .D(n31387));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n16553), .D(n31499));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n16553), .D(n31154));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n16553), .D(n31813));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n16553), .D(n31828));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n16553), .D(n31232));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n16553), .D(n31697));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n16553), .D(n31402));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n16553), .D(n32201));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n16553), .D(n32039));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n16553), .D(n31333));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n16553), .D(n31193));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n16553), .D(n31184));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n16553), .D(n30323));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n16553), .D(n30344));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n16553), .D(n31393));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17275));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n17333));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n29603), .S(n37190));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n29613), .S(n29609));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n29733), .S(n29655));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n29741), .S(n29617));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n29745), .S(n29619));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n29749), .S(n29653));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n29753), .S(n29651));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n29757), .S(n29649));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n29761), .S(n29621));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n29765), .S(n29565));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n29769), .S(n29647));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n56), .S(n29597));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n21272), .S(n21790));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_3568), .S(n29539));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n7_adj_3567), .S(n8_adj_3713));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n7_adj_3565), .S(n8_adj_3714));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_3564), .S(n8_adj_3715));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n29773), .S(n29623));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n29801), .S(n29667));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n29777), .S(n29645));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n29781), .S(n29643));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_3562), .S(n29541));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n29785), .S(n29641));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n29789), .S(n29639));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n7_adj_3560), .S(n8_adj_3716));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_3559), .S(n29543));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n29793), .S(n29637));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n7_adj_3558), .S(n21274));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n29797), .S(n21802));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7), .S(n29545));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17119));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_24_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n24672), .O(n2_adj_3702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17115));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_1127 (.I0(n15753), .I1(n15772), .I2(\data_in_frame[12] [7]), 
            .I3(n30678), .O(n10_adj_3717));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17113));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17110));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17109));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17107));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17105));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17104));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17099));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n17086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n17085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk32MHz), 
           .D(n17084));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_1128 (.I0(\data_in_frame[14] [7]), .I1(n10_adj_3717), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n30362));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31309 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3718), .I2(n34169), .I3(byte_transmit_counter[2]), 
            .O(n36954));
    defparam byte_transmit_counter_1__bdd_4_lut_31309.LUT_INIT = 16'he4aa;
    SB_LUT4 i12895_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n17282));
    defparam i12895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1129 (.I0(n30734), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3719));   // verilog/coms.v(69[16:27])
    defparam i2_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17083));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17082));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17081));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17079));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n17332));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17274));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n17305));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17074));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17073));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17072));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12896_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n17283));
    defparam i12896_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12897_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n17284));
    defparam i12897_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17071));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i11_4_lut_adj_1130 (.I0(\FRAME_MATCHER.state [20]), .I1(n22), 
            .I2(n16_adj_3579), .I3(\FRAME_MATCHER.state [25]), .O(n24_adj_3720));
    defparam i11_4_lut_adj_1130.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17273));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n17331));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_24 (.CI(n24672), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n24673));
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17270));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17070));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n17304));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17069));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12898_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30180), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n17285));
    defparam i12898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n36954_bdd_4_lut (.I0(n36954), .I1(n17_adj_3721), .I2(n16_adj_3722), 
            .I3(byte_transmit_counter[2]), .O(n36957));
    defparam n36954_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1131 (.I0(n30606), .I1(n30362), .I2(\data_in_frame[17] [4]), 
            .I3(\data_in_frame[17] [3]), .O(n14_adj_3723));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1132 (.I0(\FRAME_MATCHER.state [18]), .I1(n24_adj_3720), 
            .I2(n20), .I3(\FRAME_MATCHER.state [19]), .O(n30093));
    defparam i12_4_lut_adj_1132.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n17330));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_23_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n24671), .O(n2_adj_3700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n17329));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n17328));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n17327));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n17326));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n17325));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n17324));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n17323));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n17322));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n17321));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n17320));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17068));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1133 (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n30201));
    defparam i3_4_lut_adj_1133.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(GND_net), .I3(GND_net), .O(n63_adj_3621));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1135 (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n234));
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1136 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [15]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n10_adj_3724));
    defparam i4_4_lut_adj_1136.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1137 (.I0(\FRAME_MATCHER.state [12]), .I1(n10_adj_3724), 
            .I2(\FRAME_MATCHER.state [11]), .I3(GND_net), .O(n30203));
    defparam i5_3_lut_adj_1137.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1138 (.I0(n63_adj_3621), .I1(n30201), .I2(n30093), 
            .I3(n6_adj_3725), .O(n15264));   // verilog/coms.v(206[5:16])
    defparam i4_4_lut_adj_1138.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n15361));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'hbbbb;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17067));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_23 (.CI(n24671), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n24672));
    SB_LUT4 i2_3_lut_4_lut_adj_1140 (.I0(\FRAME_MATCHER.state [1]), .I1(n15361), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n15264), .O(n15502));   // verilog/coms.v(244[5:25])
    defparam i2_3_lut_4_lut_adj_1140.LUT_INIT = 16'hffdf;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31339 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n36948));
    defparam byte_transmit_counter_0__bdd_4_lut_31339.LUT_INIT = 16'he4aa;
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_1141 (.I0(n15501), .I1(n15361), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n15264), .O(n21813));
    defparam i2_4_lut_adj_1141.LUT_INIT = 16'haaa8;
    SB_LUT4 n36948_bdd_4_lut (.I0(n36948), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n36951));
    defparam n36948_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1142 (.I0(Kp_23__N_1405), .I1(n14_adj_3723), .I2(n10_adj_3719), 
            .I3(n15994), .O(n30516));   // verilog/coms.v(69[16:27])
    defparam i7_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 equal_120_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10));   // verilog/coms.v(154[7:23])
    defparam equal_120_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n17269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17066));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17267));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17265));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n17319));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17063));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n17318));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17062));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n17317));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17060));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17053));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n17052));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n17051));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n17050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n17049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n17048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17047));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n17046));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_114_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_3550));   // verilog/coms.v(154[7:23])
    defparam equal_114_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n17040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n17039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n17038));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n17037));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n17036));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n17035));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12871_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n17258));
    defparam i12871_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n17034));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_22_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n24670), .O(n2_adj_3698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n17033));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12874_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n17261));
    defparam i12874_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n17032));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n17031));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n17030));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n17029));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n17028));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n17027));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n17026));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n17025));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n17024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n17023));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n17022));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n17021));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n17020));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n17019));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n16772));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12872_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n17259));
    defparam i12872_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n16770));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n17018));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_1143 (.I0(n16318), .I1(n15824), .I2(n16321), 
            .I3(Kp_23__N_1327), .O(n12_adj_3726));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i12873_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n17260));
    defparam i12873_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17258));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12867_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n17254));
    defparam i12867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n16967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n16966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n16965));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12868_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n17255));
    defparam i12868_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n16964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n16963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n16962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n16961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n16960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n16959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n16958));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n16957));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n16956));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n16955));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n16954));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n16953));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n16952));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n16951));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n16950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n16949));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n16948));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n16947));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n16946));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n16944));   // verilog/coms.v(126[12] 289[6])
    SB_DFF LED_3230 (.Q(LED_c), .C(clk32MHz), .D(n30948));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12869_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n17256));
    defparam i12869_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12870_3_lut_4_lut (.I0(n10), .I1(n30190), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n17257));
    defparam i12870_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12917_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n17304));
    defparam i12917_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12918_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n17305));
    defparam i12918_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n29611));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n16903));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n16902));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n16901));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n16900));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n16899));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12919_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n17306));
    defparam i12919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12920_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n17307));
    defparam i12920_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12916_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n17303));
    defparam i12916_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12907_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n17294));
    defparam i12907_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12921_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n17308));
    defparam i12921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12922_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n17309));
    defparam i12922_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12908_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n17295));
    defparam i12908_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1144 (.I0(n26405), .I1(n12_adj_3726), .I2(\data_in_frame[19] [4]), 
            .I3(\data_in_frame[19] [3]), .O(n30474));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i12915_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30168), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n17302));
    defparam i12915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1145 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21269), .O(n30172));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1145.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1146 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21269), .O(n30168));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1146.LUT_INIT = 16'hdfff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1147 (.I0(n21269), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n30190));
    defparam i2_2_lut_3_lut_4_lut_adj_1147.LUT_INIT = 16'hff7f;
    SB_LUT4 i12909_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n17296));
    defparam i12909_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1148 (.I0(n21269), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n30176));
    defparam i2_2_lut_3_lut_4_lut_adj_1148.LUT_INIT = 16'hfff7;
    SB_CARRY add_44_4 (.CI(n24652), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n24653));
    SB_LUT4 i12910_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n17297));
    defparam i12910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1149 (.I0(n15704), .I1(n30542), .I2(n30232), 
            .I3(\data_in_frame[6] [2]), .O(n16318));   // verilog/coms.v(70[16:41])
    defparam i3_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30634));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17264));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_22 (.CI(n24670), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n24671));
    SB_LUT4 i12911_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n17298));
    defparam i12911_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12912_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n17299));
    defparam i12912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n17316));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n17315));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12913_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n17300));
    defparam i12913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_21_lut (.I0(n1731), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n24669), .O(n2_adj_3696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1151 (.I0(\data_in_frame[19] [2]), .I1(n30634), 
            .I2(\data_in_frame[14] [7]), .I3(n16318), .O(n10_adj_3727));
    defparam i4_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i12914_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30172), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n17301));
    defparam i12914_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1152 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21269), .O(n30164));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1152.LUT_INIT = 16'hfbff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31300 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n36942));
    defparam byte_transmit_counter_0__bdd_4_lut_31300.LUT_INIT = 16'he4aa;
    SB_LUT4 n36942_bdd_4_lut (.I0(n36942), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n36945));
    defparam n36942_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12835_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n17222));
    defparam i12835_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12836_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n17223));
    defparam i12836_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12837_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n17224));
    defparam i12837_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1153 (.I0(n21269), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n30180));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1153.LUT_INIT = 16'hfffd;
    SB_LUT4 i12838_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n17225));
    defparam i12838_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12839_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n17226));
    defparam i12839_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12840_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n17227));
    defparam i12840_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12841_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n17228));
    defparam i12841_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12842_3_lut_4_lut (.I0(n10), .I1(n30176), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n17229));
    defparam i12842_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31295 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n36936));
    defparam byte_transmit_counter_0__bdd_4_lut_31295.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1019_i24_3_lut (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4311), .I3(GND_net), .O(n4335));
    defparam mux_1019_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i1_3_lut (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4311), .I3(GND_net), .O(n4312));
    defparam mux_1019_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i23_3_lut (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4311), .I3(GND_net), .O(n4334));
    defparam mux_1019_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i22_3_lut (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4311), .I3(GND_net), .O(n4333));
    defparam mux_1019_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i21_3_lut (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4311), .I3(GND_net), .O(n4332));
    defparam mux_1019_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i20_3_lut (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4311), .I3(GND_net), .O(n4331));
    defparam mux_1019_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i19_3_lut (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4311), .I3(GND_net), .O(n4330));
    defparam mux_1019_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i18_3_lut (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4311), .I3(GND_net), .O(n4329));
    defparam mux_1019_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n36936_bdd_4_lut (.I0(n36936), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n36939));
    defparam n36936_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31290 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n36930));
    defparam byte_transmit_counter_0__bdd_4_lut_31290.LUT_INIT = 16'he4aa;
    SB_LUT4 n36930_bdd_4_lut (.I0(n36930), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n36933));
    defparam n36930_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31285 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n36924));
    defparam byte_transmit_counter_0__bdd_4_lut_31285.LUT_INIT = 16'he4aa;
    SB_LUT4 n36924_bdd_4_lut (.I0(n36924), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n36927));
    defparam n36924_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31280 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n36918));
    defparam byte_transmit_counter_0__bdd_4_lut_31280.LUT_INIT = 16'he4aa;
    SB_LUT4 n36918_bdd_4_lut (.I0(n36918), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n36921));
    defparam n36918_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1154 (.I0(n3915), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n5784), .I3(GND_net), .O(n16553));
    defparam i1_2_lut_3_lut_adj_1154.LUT_INIT = 16'h0202;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31275 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n36912));
    defparam byte_transmit_counter_0__bdd_4_lut_31275.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1155 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[5] [6]), .O(n30522));
    defparam i2_3_lut_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1019_i17_3_lut (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4311), .I3(GND_net), .O(n4328));
    defparam mux_1019_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i16_3_lut (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4311), .I3(GND_net), .O(n4327));
    defparam mux_1019_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1156 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[7] [1]), .O(n1237));
    defparam i1_2_lut_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 n36912_bdd_4_lut (.I0(n36912), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n36915));
    defparam n36912_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31270 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n36906));
    defparam byte_transmit_counter_0__bdd_4_lut_31270.LUT_INIT = 16'he4aa;
    SB_LUT4 n36906_bdd_4_lut (.I0(n36906), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n36909));
    defparam n36906_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1157 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(n30793), .I3(GND_net), .O(n15506));
    defparam i1_2_lut_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31265 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n36900));
    defparam byte_transmit_counter_0__bdd_4_lut_31265.LUT_INIT = 16'he4aa;
    SB_LUT4 n36900_bdd_4_lut (.I0(n36900), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n36903));
    defparam n36900_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[16] [5]), .I1(n16356), .I2(\data_out_frame[18] [7]), 
            .I3(n27213), .O(n10_adj_3728));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31260 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n36882));
    defparam byte_transmit_counter_0__bdd_4_lut_31260.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1158 (.I0(\data_out_frame[7] [2]), .I1(n30793), 
            .I2(n30548), .I3(n30365), .O(n15054));
    defparam i2_3_lut_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1159 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [5]), .I3(GND_net), .O(n30548));
    defparam i1_2_lut_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i15_3_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4311), .I3(GND_net), .O(n4326));
    defparam mux_1019_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i14_3_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4311), .I3(GND_net), .O(n4325));
    defparam mux_1019_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n36882_bdd_4_lut (.I0(n36882), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n36885));
    defparam n36882_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1019_i13_3_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4311), .I3(GND_net), .O(n4324));
    defparam mux_1019_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1160 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[5] [6]), .O(n6_adj_3729));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1019_i12_3_lut (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4311), .I3(GND_net), .O(n4323));
    defparam mux_1019_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1161 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(n15863), .I3(n30224), .O(n30698));
    defparam i1_2_lut_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1019_i11_3_lut (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4311), .I3(GND_net), .O(n4322));
    defparam mux_1019_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(\data_out_frame[15] [0]), .I1(n15863), 
            .I2(n30224), .I3(GND_net), .O(n27167));
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i10_3_lut (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4311), .I3(GND_net), .O(n4321));
    defparam mux_1019_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1163 (.I0(n16214), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[13] [5]), .I3(GND_net), .O(n30781));
    defparam i1_2_lut_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i9_3_lut (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4311), .I3(GND_net), .O(n4320));
    defparam mux_1019_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i8_3_lut (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4311), .I3(GND_net), .O(n4319));
    defparam mux_1019_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1164 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(n30588), .I3(GND_net), .O(n6_adj_3730));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i7_3_lut (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4311), .I3(GND_net), .O(n4318));
    defparam mux_1019_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1165 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[11] [0]), .O(n30588));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1166 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[6] [6]), 
            .I2(n30770), .I3(GND_net), .O(n30559));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1167 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n30770));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i6_3_lut (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4311), .I3(GND_net), .O(n4317));
    defparam mux_1019_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1168 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n30315));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n30695));
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1019_i5_3_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4311), .I3(GND_net), .O(n4316));
    defparam mux_1019_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i4_3_lut (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4311), .I3(GND_net), .O(n4315));
    defparam mux_1019_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1019_i3_3_lut (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4311), .I3(GND_net), .O(n4314));
    defparam mux_1019_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_1170 (.I0(n21540), .I1(n18518), .I2(n22054), 
            .I3(GND_net), .O(n31259));
    defparam i3_3_lut_adj_1170.LUT_INIT = 16'hfbfb;
    SB_LUT4 mux_1019_i2_3_lut (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4311), .I3(GND_net), .O(n4313));
    defparam mux_1019_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1171 (.I0(n15880), .I1(\data_out_frame[14] [7]), 
            .I2(n15630), .I3(GND_net), .O(n6_adj_3731));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n16_adj_3732));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1172 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n30701), .I3(GND_net), .O(n6_adj_3733));
    defparam i1_2_lut_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1173 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [5]), 
            .I2(n10_adj_3734), .I3(n30565), .O(n30572));
    defparam i5_3_lut_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1174 (.I0(\data_out_frame[20] [2]), .I1(n30322), 
            .I2(n26487), .I3(n30441), .O(n31184));
    defparam i2_3_lut_4_lut_adj_1174.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1175 (.I0(\FRAME_MATCHER.state[3] ), .I1(n2421), 
            .I2(n13117), .I3(n67), .O(n29613));
    defparam i1_3_lut_4_lut_adj_1175.LUT_INIT = 16'haa80;
    SB_LUT4 i1_2_lut_3_lut_adj_1176 (.I0(n15495), .I1(n740), .I2(n13117), 
            .I3(GND_net), .O(n1));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_1176.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1177 (.I0(\data_in_frame[6] [6]), .I1(Kp_23__N_823), 
            .I2(\data_in_frame[4] [4]), .I3(n15573), .O(n16360));
    defparam i1_2_lut_3_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1178 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[15] [7]), 
            .I2(n26635), .I3(GND_net), .O(n30778));
    defparam i1_2_lut_3_lut_adj_1178.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1179 (.I0(\FRAME_MATCHER.state [1]), .I1(n15264), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n15361), .O(n15504));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_4_lut_adj_1179.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_adj_1180 (.I0(\FRAME_MATCHER.state [1]), .I1(n15264), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n15369), .O(n63_adj_3660));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_4_lut_adj_1180.LUT_INIT = 16'hffef;
    SB_LUT4 i17459_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n15493), .I3(n21813), .O(n2430));   // verilog/coms.v(148[5:9])
    defparam i17459_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i12960_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n17347));
    defparam i12960_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12961_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n17348));
    defparam i12961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_adj_1181 (.I0(n63), .I1(n740), .I2(n31), .I3(n15495), 
            .O(n5_adj_3));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut_adj_1181.LUT_INIT = 16'ha0a2;
    SB_LUT4 i17395_2_lut_3_lut (.I0(n63), .I1(n740), .I2(n93[1]), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2396 [1]));   // verilog/coms.v(157[6] 159[9])
    defparam i17395_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i31196_2_lut_3_lut (.I0(\r_SM_Main_2__N_3259[0] ), .I1(tx_active), 
            .I2(n22044), .I3(GND_net), .O(tx_transmit_N_3151));   // verilog/coms.v(126[12] 289[6])
    defparam i31196_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_3_lut_adj_1182 (.I0(\r_SM_Main_2__N_3259[0] ), .I1(tx_active), 
            .I2(n22044), .I3(GND_net), .O(n961));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1182.LUT_INIT = 16'hefef;
    SB_LUT4 i12928_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n17315));
    defparam i12928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12929_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n17316));
    defparam i12929_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1183 (.I0(n30417), .I1(n10_adj_3727), .I2(\data_in_frame[17] [0]), 
            .I3(GND_net), .O(n30329));
    defparam i5_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i12930_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n17317));
    defparam i12930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(n26452), .I1(n30329), .I2(GND_net), 
            .I3(GND_net), .O(n30594));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i12923_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n17310));
    defparam i12923_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12924_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n17311));
    defparam i12924_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12925_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n17312));
    defparam i12925_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12926_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n17313));
    defparam i12926_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12962_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n17349));
    defparam i12962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1185 (.I0(\data_in_frame[5] [0]), .I1(n30368), 
            .I2(n30666), .I3(n30648), .O(n6_adj_3590));
    defparam i1_2_lut_3_lut_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i12927_3_lut_4_lut (.I0(n10_adj_3550), .I1(n30164), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n17314));
    defparam i12927_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i25324_3_lut_4_lut (.I0(n15369), .I1(n15493), .I2(LED_c), 
            .I3(n13117), .O(n30948));   // verilog/coms.v(148[5:9])
    defparam i25324_3_lut_4_lut.LUT_INIT = 16'he0ee;
    SB_LUT4 i12859_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n17246));
    defparam i12859_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12860_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n17247));
    defparam i12860_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12861_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n17248));
    defparam i12861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12955_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n17342));
    defparam i12955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12956_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n17343));
    defparam i12956_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12862_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n17249));
    defparam i12862_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12863_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n17250));
    defparam i12863_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12864_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n17251));
    defparam i12864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12865_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n17252));
    defparam i12865_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12866_3_lut_4_lut (.I0(n10), .I1(n30164), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n17253));
    defparam i12866_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3722));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3721));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12513_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[0] ), .O(n16900));
    defparam i12513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3736));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29215_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34853));   // verilog/coms.v(104[34:55])
    defparam i29215_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3737));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26902_4_lut (.I0(n19_adj_3736), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n32539));
    defparam i26902_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26903_3_lut (.I0(n36999), .I1(n32539), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32540));
    defparam i26903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26940_4_lut (.I0(n5_adj_3737), .I1(n34853), .I2(n32644), 
            .I3(byte_transmit_counter[0]), .O(n32577));
    defparam i26940_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26942_4_lut (.I0(n32577), .I1(n32540), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32579));
    defparam i26942_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26941_3_lut (.I0(n36909), .I1(n36903), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32578));
    defparam i26941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3738));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29211_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34849));   // verilog/coms.v(104[34:55])
    defparam i29211_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3739));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26899_4_lut (.I0(n19_adj_3738), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n32536));
    defparam i26899_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26900_3_lut (.I0(n37047), .I1(n32536), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32537));
    defparam i26900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26937_4_lut (.I0(n5_adj_3739), .I1(n34849), .I2(n32644), 
            .I3(byte_transmit_counter[0]), .O(n32574));
    defparam i26937_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26939_4_lut (.I0(n32574), .I1(n32537), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32576));
    defparam i26939_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26938_3_lut (.I0(n36921), .I1(n36915), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32575));
    defparam i26938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12515_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n16902));
    defparam i12515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12516_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [0]), 
            .I3(PWMLimit[0]), .O(n16903));
    defparam i12516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n34844));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3740));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26934_4_lut (.I0(n5_adj_3740), .I1(byte_transmit_counter[0]), 
            .I2(n32644), .I3(n34844), .O(n32571));
    defparam i26934_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26936_4_lut (.I0(n32571), .I1(n36957), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32573));
    defparam i26936_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26935_3_lut (.I0(n36933), .I1(n36927), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32572));
    defparam i26935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12557_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [7]), 
            .I3(gearBoxRatio[23]), .O(n16944));
    defparam i12557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30158_3_lut (.I0(n37017), .I1(n36885), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n35797));
    defparam i30158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30162_3_lut (.I0(n36987), .I1(n35797), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n35801));   // verilog/coms.v(104[34:55])
    defparam i30162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30163_4_lut (.I0(n35801), .I1(n36963), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i30163_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12559_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [6]), 
            .I3(gearBoxRatio[22]), .O(n16946));
    defparam i12559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28885_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n34271));   // verilog/coms.v(104[34:55])
    defparam i28885_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n34271), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3741));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3742));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12560_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [5]), 
            .I3(gearBoxRatio[21]), .O(n16947));
    defparam i12560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i26931_3_lut (.I0(n5_adj_3742), .I1(n6_adj_3741), .I2(n32644), 
            .I3(GND_net), .O(n32568));
    defparam i26931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26933_4_lut (.I0(n32568), .I1(n36969), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32570));
    defparam i26933_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26932_3_lut (.I0(n36945), .I1(n36939), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32569));
    defparam i26932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12561_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [4]), 
            .I3(gearBoxRatio[20]), .O(n16948));
    defparam i12561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29256_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n34268));   // verilog/coms.v(104[34:55])
    defparam i29256_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(n34268), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3743));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3744));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26928_3_lut (.I0(n5_adj_3744), .I1(n6_adj_3743), .I2(n32644), 
            .I3(GND_net), .O(n32565));
    defparam i26928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26930_4_lut (.I0(n32565), .I1(n36975), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32567));
    defparam i26930_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12562_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [3]), 
            .I3(gearBoxRatio[19]), .O(n16949));
    defparam i12562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i26929_3_lut (.I0(n37041), .I1(n36951), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n32566));
    defparam i26929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12563_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [2]), 
            .I3(gearBoxRatio[18]), .O(n16950));
    defparam i12563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12564_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [1]), 
            .I3(gearBoxRatio[17]), .O(n16951));
    defparam i12564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12565_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[17] [0]), 
            .I3(gearBoxRatio[16]), .O(n16952));
    defparam i12565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12957_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n17344));
    defparam i12957_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12566_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [7]), 
            .I3(gearBoxRatio[15]), .O(n16953));
    defparam i12566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29188_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34825));   // verilog/coms.v(104[34:55])
    defparam i29188_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i12567_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [6]), 
            .I3(gearBoxRatio[14]), .O(n16954));
    defparam i12567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3745));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26925_4_lut (.I0(n5_adj_3745), .I1(n34825), .I2(n32644), 
            .I3(byte_transmit_counter[0]), .O(n32562));
    defparam i26925_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26927_4_lut (.I0(n32562), .I1(n36981), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n32564));
    defparam i26927_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12568_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [5]), 
            .I3(gearBoxRatio[13]), .O(n16955));
    defparam i12568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12569_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [4]), 
            .I3(gearBoxRatio[12]), .O(n16956));
    defparam i12569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12570_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [3]), 
            .I3(gearBoxRatio[11]), .O(n16957));
    defparam i12570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12571_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [2]), 
            .I3(gearBoxRatio[10]), .O(n16958));
    defparam i12571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12572_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [1]), 
            .I3(gearBoxRatio[9]), .O(n16959));
    defparam i12572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1186 (.I0(n30474), .I1(n30594), .I2(n30516), 
            .I3(n30494), .O(n26930));
    defparam i3_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i12573_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[18] [0]), 
            .I3(gearBoxRatio[8]), .O(n16960));
    defparam i12573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12574_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [7]), 
            .I3(gearBoxRatio[7]), .O(n16961));
    defparam i12574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12958_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n17345));
    defparam i12958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12575_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [6]), 
            .I3(gearBoxRatio[6]), .O(n16962));
    defparam i12575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12576_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [5]), 
            .I3(gearBoxRatio[5]), .O(n16963));
    defparam i12576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12577_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [4]), 
            .I3(gearBoxRatio[4]), .O(n16964));
    defparam i12577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12578_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [3]), 
            .I3(gearBoxRatio[3]), .O(n16965));
    defparam i12578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12579_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [2]), 
            .I3(gearBoxRatio[2]), .O(n16966));
    defparam i12579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12959_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30180), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n17346));
    defparam i12959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12580_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [1]), 
            .I3(gearBoxRatio[1]), .O(n16967));
    defparam i12580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[14] [6]), .I1(n15704), 
            .I2(GND_net), .I3(GND_net), .O(n30603));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1188 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n15421), .I3(\FRAME_MATCHER.i [4]), .O(n15239));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1188.LUT_INIT = 16'hfffe;
    SB_LUT4 i12385_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[19] [0]), 
            .I3(gearBoxRatio[0]), .O(n16772));
    defparam i12385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12690_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[1] ), .O(n17077));
    defparam i12690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1189 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n10_adj_3552));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_adj_1189.LUT_INIT = 16'hefef;
    SB_LUT4 i12691_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[2] ), .O(n17078));
    defparam i12691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29204_2_lut (.I0(\data_out_frame[22] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34169));
    defparam i29204_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3718));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1190 (.I0(\data_in_frame[19] [1]), .I1(n30603), 
            .I2(n15604), .I3(Kp_23__N_1280), .O(n16_adj_3746));
    defparam i6_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i17173_4_lut (.I0(n21283), .I1(n31_adj_3642), .I2(n31_c), 
            .I3(\FRAME_MATCHER.state [1]), .O(n21540));
    defparam i17173_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1191 (.I0(n5784), .I1(n21540), .I2(\FRAME_MATCHER.state_31__N_2428 [3]), 
            .I3(n5782), .O(n16549));
    defparam i1_4_lut_adj_1191.LUT_INIT = 16'ha022;
    SB_LUT4 i7_4_lut_adj_1192 (.I0(n30426), .I1(n30761), .I2(n16149), 
            .I3(n30707), .O(n17_adj_3747));
    defparam i7_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1193 (.I0(n17_adj_3747), .I1(\data_in_frame[18] [7]), 
            .I2(n16_adj_3746), .I3(\data_in_frame[16] [3]), .O(n26452));
    defparam i9_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1194 (.I0(n30601), .I1(n30417), .I2(\data_in_frame[19] [0]), 
            .I3(\data_in_frame[16] [4]), .O(n26767));
    defparam i3_4_lut_adj_1194.LUT_INIT = 16'h9669;
    SB_LUT4 i12692_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[3] ), .O(n17079));
    defparam i12692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_in_frame[15] [7]), .I1(n26635), 
            .I2(GND_net), .I3(GND_net), .O(n30624));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i12693_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[4] ), .O(n17080));
    defparam i12693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12694_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[5] ), .O(n17081));
    defparam i12694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12695_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[6] ), .O(n17082));
    defparam i12695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12696_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[7] ), .O(n17083));
    defparam i12696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13003_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n17390));
    defparam i13003_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16906_2_lut_3_lut (.I0(n21813), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n21269));
    defparam i16906_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\FRAME_MATCHER.state [26]), .I1(n32330), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3716));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1197 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n15224), .O(n15501));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1197.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut_adj_1198 (.I0(\FRAME_MATCHER.state [12]), .I1(n10_adj_3724), 
            .I2(\FRAME_MATCHER.state [11]), .I3(n234), .O(n6_adj_3725));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_4_lut_adj_1198.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1199 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n15358));   // verilog/coms.v(225[5:23])
    defparam i1_2_lut_3_lut_adj_1199.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1200 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n15493), .I3(GND_net), .O(n15495));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_1200.LUT_INIT = 16'hfbfb;
    SB_LUT4 i17529_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[3]), 
            .O(n21899));
    defparam i17529_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\FRAME_MATCHER.state [18]), .I1(n32330), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3715));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1202 (.I0(\data_in[1] [3]), .I1(\data_in[2] [7]), 
            .I2(n10_adj_3664), .I3(\data_in[3] [4]), .O(n5_adj_3649));
    defparam i1_2_lut_4_lut_adj_1202.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\FRAME_MATCHER.state [17]), .I1(n32330), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3714));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_1204 (.I0(n61), .I1(n15495), .I2(n133), .I3(n13185), 
            .O(n32330));
    defparam i2_4_lut_adj_1204.LUT_INIT = 16'h0405;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\FRAME_MATCHER.state [16]), .I1(n32330), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3713));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1206 (.I0(n2421), .I1(n2857), .I2(n15504), .I3(GND_net), 
            .O(n30199));
    defparam i1_3_lut_adj_1206.LUT_INIT = 16'habab;
    SB_LUT4 i13004_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n17391));
    defparam i13004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13005_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n17392));
    defparam i13005_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13006_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n17393));
    defparam i13006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13007_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n17394));
    defparam i13007_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13008_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n17395));
    defparam i13008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1207 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n15264), .I3(GND_net), .O(n15493));   // verilog/coms.v(195[5:24])
    defparam i1_2_lut_3_lut_adj_1207.LUT_INIT = 16'hfefe;
    SB_LUT4 i13009_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n17396));
    defparam i13009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1208 (.I0(\data_in_frame[14] [7]), .I1(n10_adj_3717), 
            .I2(\data_in_frame[15] [1]), .I3(n30634), .O(n6_adj_3647));
    defparam i1_2_lut_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_1209 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n12846));
    defparam i1_4_lut_4_lut_adj_1209.LUT_INIT = 16'h2034;
    SB_LUT4 i1_2_lut_3_lut_adj_1210 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[14] [6]), 
            .I2(n30291), .I3(GND_net), .O(n34));
    defparam i1_2_lut_3_lut_adj_1210.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1211 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [7]), 
            .I2(n26712), .I3(GND_net), .O(n30722));
    defparam i1_2_lut_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(Kp_23__N_823), .I1(\data_in_frame[4] [4]), 
            .I2(n15573), .I3(GND_net), .O(n30458));
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 equal_1126_i9_3_lut_4_lut (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(n30429), .O(n30212));   // verilog/coms.v(230[9:81])
    defparam equal_1126_i9_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1213 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n16114));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1214 (.I0(\data_in_frame[9] [4]), .I1(n26493), 
            .I2(n16208), .I3(GND_net), .O(n30666));
    defparam i1_2_lut_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i13010_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [1]), 
            .I3(PWMLimit[1]), .O(n17397));
    defparam i13010_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13011_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [2]), 
            .I3(PWMLimit[2]), .O(n17398));
    defparam i13011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13012_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [3]), 
            .I3(PWMLimit[3]), .O(n17399));
    defparam i13012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13013_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [4]), 
            .I3(PWMLimit[4]), .O(n17400));
    defparam i13013_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13014_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [5]), 
            .I3(PWMLimit[5]), .O(n17401));
    defparam i13014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1215 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[7] [5]), 
            .I2(\data_in_frame[7] [4]), .I3(\data_in_frame[7] [6]), .O(n30374));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1216 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n30288));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1217 (.I0(n27227), .I1(Kp_23__N_832), .I2(\data_in_frame[4] [7]), 
            .I3(\data_in_frame[7] [3]), .O(n16262));   // verilog/coms.v(77[16:35])
    defparam i2_3_lut_4_lut_adj_1217.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1218 (.I0(Kp_23__N_794), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[1] [0]), .O(n30393));   // verilog/coms.v(68[16:69])
    defparam i2_3_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1219 (.I0(n27165), .I1(\data_in_frame[15] [5]), 
            .I2(n16146), .I3(n30340), .O(n30426));
    defparam i1_2_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1220 (.I0(Kp_23__N_823), .I1(\data_in_frame[4] [4]), 
            .I2(\data_in_frame[6] [5]), .I3(n16067), .O(n30725));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1221 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(n15746), .I3(\data_in_frame[8] [6]), .O(n30420));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1222 (.I0(\data_in_frame[6] [3]), .I1(n15671), 
            .I2(\data_in_frame[8] [5]), .I3(GND_net), .O(n30221));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1223 (.I0(\data_in_frame[5] [7]), .I1(n30404), 
            .I2(\data_in_frame[10] [2]), .I3(GND_net), .O(n4_adj_3603));
    defparam i1_2_lut_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1224 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[16] [4]), .I3(\data_in_frame[16] [2]), .O(n15982));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n30761));
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1226 (.I0(Kp_23__N_962), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[12] [2]), .I3(\data_in_frame[9] [6]), .O(n30758));
    defparam i2_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(n740), .I1(n13117), .I2(GND_net), .I3(GND_net), 
            .O(n13185));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h4444;
    SB_LUT4 i13015_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [6]), 
            .I3(PWMLimit[6]), .O(n17402));
    defparam i13015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i113_3_lut (.I0(n15502), .I1(n961), .I2(n13117), .I3(GND_net), 
            .O(n54));   // verilog/coms.v(113[11:12])
    defparam i113_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut_adj_1228 (.I0(n15504), .I1(n2857), .I2(n13117), .I3(GND_net), 
            .O(n61));   // verilog/coms.v(216[5:21])
    defparam i1_3_lut_adj_1228.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[13] [4]), .I3(GND_net), .O(n15636));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1230 (.I0(n15501), .I1(n3761), .I2(n13117), .I3(GND_net), 
            .O(n67));   // verilog/coms.v(244[5:25])
    defparam i1_3_lut_adj_1230.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(n2421), .I1(n13117), .I2(GND_net), 
            .I3(GND_net), .O(n133));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h8888;
    SB_LUT4 i13016_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[7] [7]), 
            .I3(PWMLimit[7]), .O(n17403));
    defparam i13016_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1232 (.I0(\FRAME_MATCHER.state[3] ), .I1(n61), 
            .I2(n1), .I3(n54), .O(n7_adj_3748));   // verilog/coms.v(113[11:12])
    defparam i1_4_lut_adj_1232.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_1233 (.I0(n15358), .I1(n7_adj_3748), .I2(n15224), 
            .I3(\FRAME_MATCHER.state_31__N_2428 [3]), .O(n29609));   // verilog/coms.v(113[11:12])
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'hcdcc;
    SB_LUT4 i2_3_lut_4_lut_adj_1234 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[15] [3]), 
            .I2(n15604), .I3(\data_in_frame[15] [2]), .O(n30359));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i13017_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [0]), 
            .I3(PWMLimit[8]), .O(n17404));
    defparam i13017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(\data_in_frame[7] [1]), .I1(n15573), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n30480));
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i25267_2_lut (.I0(n15501), .I1(n3761), .I2(GND_net), .I3(GND_net), 
            .O(n30890));
    defparam i25267_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32579), .I3(n32578), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i2_3_lut_4_lut_adj_1236 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[12] [7]), .O(n30528));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 select_355_Select_1_i5_4_lut (.I0(n63), .I1(n15504), .I2(n2857), 
            .I3(n93[1]), .O(n5_adj_3749));
    defparam select_355_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i5_3_lut_4_lut_adj_1237 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[7] [1]), .I3(n16255), .O(n14_adj_3593));
    defparam i5_3_lut_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1238 (.I0(n93[1]), .I1(n5_adj_3749), .I2(n30890), 
            .I3(n63), .O(n6_adj_3750));
    defparam i2_4_lut_adj_1238.LUT_INIT = 16'hcecf;
    SB_LUT4 i3_4_lut_adj_1239 (.I0(n15494), .I1(n6_adj_3750), .I2(\FRAME_MATCHER.state_31__N_2396 [1]), 
            .I3(n15495), .O(n37190));
    defparam i3_4_lut_adj_1239.LUT_INIT = 16'hddfd;
    SB_LUT4 i13018_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [1]), 
            .I3(PWMLimit[9]), .O(n17405));
    defparam i13018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32576), .I3(n32575), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13019_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [2]), 
            .I3(PWMLimit[10]), .O(n17406));
    defparam i13019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(n26493), .I1(n16208), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n27225));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1241 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[19] [6]), .I3(n16321), .O(n30734));
    defparam i2_3_lut_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1242 (.I0(Kp_23__N_962), .I1(n30235), .I2(\data_in_frame[5] [6]), 
            .I3(n16302), .O(n10_adj_3589));   // verilog/coms.v(72[16:43])
    defparam i2_2_lut_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(n22_adj_3586), 
            .I2(\data_in_frame[18] [7]), .I3(\data_in_frame[18] [6]), .O(n25));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1243 (.I0(n30343), .I1(n30716), .I2(\data_out_frame[20] [6]), 
            .I3(GND_net), .O(n31393));
    defparam i2_3_lut_adj_1243.LUT_INIT = 16'h6969;
    SB_LUT4 i13020_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [3]), 
            .I3(PWMLimit[11]), .O(n17407));
    defparam i13020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(n30450), .I1(n30343), .I2(GND_net), 
            .I3(GND_net), .O(n30344));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(n30450), .I1(n30322), .I2(GND_net), 
            .I3(GND_net), .O(n30323));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1246 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[7] [2]), .I3(\data_in_frame[9] [2]), .O(n6_adj_3585));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(n30302), .I1(n16389), .I2(\data_out_frame[20] [0]), 
            .I3(n30582), .O(n10_adj_3751));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1248 (.I0(\data_out_frame[19] [6]), .I1(n10_adj_3751), 
            .I2(\data_out_frame[20] [1]), .I3(GND_net), .O(n31333));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1248.LUT_INIT = 16'h6969;
    SB_LUT4 i13021_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [4]), 
            .I3(PWMLimit[12]), .O(n17408));
    defparam i13021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(n26487), .I1(n30441), .I2(GND_net), 
            .I3(GND_net), .O(n27271));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1250 (.I0(\data_out_frame[18] [0]), .I1(n30691), 
            .I2(n30257), .I3(n30781), .O(n16_adj_3752));
    defparam i6_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1251 (.I0(n30447), .I1(n30752), .I2(\data_out_frame[6] [4]), 
            .I3(n30565), .O(n17_adj_3753));
    defparam i7_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1252 (.I0(n17_adj_3753), .I1(n30298), .I2(n16_adj_3752), 
            .I3(\data_out_frame[15] [6]), .O(n30441));
    defparam i9_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1253 (.I0(n15781), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[16] [0]), .I3(n26717), .O(n30672));
    defparam i2_3_lut_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_1254 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n4_c));
    defparam i1_4_lut_4_lut_adj_1254.LUT_INIT = 16'h1110;
    SB_LUT4 i3_4_lut_adj_1255 (.I0(\data_out_frame[19] [7]), .I1(n30572), 
            .I2(n30302), .I3(\data_out_frame[17] [3]), .O(n15085));
    defparam i3_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30565));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1257 (.I0(n15760), .I1(n30695), .I2(\data_out_frame[17] [7]), 
            .I3(n26362), .O(n10_adj_3734));
    defparam i4_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1258 (.I0(n15085), .I1(\data_out_frame[16] [7]), 
            .I2(n30582), .I3(n27213), .O(n18_adj_3754));
    defparam i7_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1259 (.I0(n26378), .I1(n18_adj_3754), .I2(n30435), 
            .I3(n30764), .O(n20_adj_3755));
    defparam i9_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n18518));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'h1010;
    SB_LUT4 i10_4_lut_adj_1261 (.I0(n15_adj_3756), .I1(n20_adj_3755), .I2(n27167), 
            .I3(n27271), .O(n32039));
    defparam i10_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1262 (.I0(n32039), .I1(n16389), .I2(n30572), 
            .I3(n6_adj_3733), .O(n32201));
    defparam i4_4_lut_adj_1262.LUT_INIT = 16'h9669;
    SB_LUT4 i28823_2_lut_3_lut (.I0(n22054), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n34460));
    defparam i28823_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30284));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut_adj_1264 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_3757));
    defparam i4_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1265 (.I0(\data_out_frame[20] [4]), .I1(n15034), 
            .I2(n27257), .I3(\data_out_frame[16] [1]), .O(n13_adj_3758));
    defparam i5_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32573), .I3(n32572), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32570), .I3(n32569), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i7_4_lut_adj_1266 (.I0(n13_adj_3758), .I1(n32059), .I2(n12_adj_3757), 
            .I3(n16042), .O(n30450));
    defparam i7_4_lut_adj_1266.LUT_INIT = 16'h9669;
    SB_LUT4 i25195_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n22054), .I3(n2_adj_3759), .O(n30807));
    defparam i25195_4_lut_4_lut.LUT_INIT = 16'hfbf8;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(n30787), .I1(n30208), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3760));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1268 (.I0(n30691), .I1(n30728), .I2(\data_out_frame[15] [7]), 
            .I3(n30438), .O(n12_adj_3761));
    defparam i5_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1269 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[6] [6]), 
            .I2(n12_adj_3761), .I3(n8_adj_3760), .O(n6_adj_3762));
    defparam i1_4_lut_adj_1269.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1270 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[16] [1]), 
            .I2(n27257), .I3(n6_adj_3762), .O(n32059));
    defparam i4_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1271 (.I0(n30731), .I1(n30350), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3763));
    defparam i2_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1272 (.I0(\data_out_frame[20] [5]), .I1(n27257), 
            .I2(n6_adj_3763), .I3(n30645), .O(n30343));
    defparam i1_4_lut_adj_1272.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n26487), .I1(\data_out_frame[20] [3]), 
            .I2(n32059), .I3(GND_net), .O(n30322));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h6969;
    SB_LUT4 i13022_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [5]), 
            .I3(PWMLimit[13]), .O(n17409));
    defparam i13022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n2_adj_3759));
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1275 (.I0(\data_in_frame[16] [3]), .I1(n30600), 
            .I2(n30675), .I3(GND_net), .O(n27261));
    defparam i1_2_lut_3_lut_adj_1275.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n30322), .I1(n30343), .I2(n30371), 
            .I3(n6_adj_3548), .O(n26378));
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1277 (.I0(\data_in_frame[13] [1]), .I1(n30554), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[10] [5]), .O(n10_adj_3575));   // verilog/coms.v(69[16:27])
    defparam i2_2_lut_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32561), .I3(n37029), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i4_4_lut_adj_1278 (.I0(n30701), .I1(n26487), .I2(n26378), 
            .I3(n30716), .O(n10_adj_3764));
    defparam i4_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1279 (.I0(n30657), .I1(n10_adj_3764), .I2(n27001), 
            .I3(GND_net), .O(n31402));
    defparam i5_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1280 (.I0(n30746), .I1(n30208), .I2(\data_out_frame[8] [5]), 
            .I3(n30559), .O(n15624));   // verilog/coms.v(72[16:27])
    defparam i2_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i13023_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [6]), 
            .I3(PWMLimit[14]), .O(n17410));
    defparam i13023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13024_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[6] [7]), 
            .I3(PWMLimit[15]), .O(n17411));
    defparam i13024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(\data_out_frame[17] [2]), .I1(n30657), 
            .I2(n30486), .I3(n30392), .O(n31697));
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1282 (.I0(n15880), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[15] [2]), .I3(\data_out_frame[13] [0]), 
            .O(n12_adj_3765));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1283 (.I0(\data_out_frame[13] [1]), .I1(n12_adj_3765), 
            .I2(n30617), .I3(n1595), .O(n16389));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32564), .I3(n37023), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i3_4_lut_adj_1284 (.I0(\data_out_frame[15] [1]), .I1(n16389), 
            .I2(\data_out_frame[19] [4]), .I3(n15541), .O(n30486));
    defparam i3_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1285 (.I0(\data_out_frame[17] [3]), .I1(n30533), 
            .I2(n30486), .I3(\data_out_frame[17] [1]), .O(n31232));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1286 (.I0(\data_out_frame[19] [3]), .I1(n30224), 
            .I2(n16377), .I3(n6_adj_3544), .O(n30533));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_out_frame[15] [1]), .I1(n30669), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3766));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1288 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(n30533), .I3(n6_adj_3766), .O(n31828));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(n31361), .I1(n30669), .I2(n30501), 
            .I3(\data_out_frame[17] [1]), .O(n31813));
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'h9669;
    SB_LUT4 i13025_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [0]), 
            .I3(PWMLimit[16]), .O(n17412));
    defparam i13025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(n15532), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15986));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i13026_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [1]), 
            .I3(PWMLimit[17]), .O(n17413));
    defparam i13026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1291 (.I0(n15986), .I1(n30513), .I2(n1967), .I3(\data_out_frame[19] [1]), 
            .O(n31154));
    defparam i3_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1292 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(n30548), .I3(\data_out_frame[6] [2]), .O(n18_adj_3767));
    defparam i7_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1293 (.I0(n27173), .I1(n18_adj_3767), .I2(n30365), 
            .I3(n30743), .O(n20_adj_3768));
    defparam i9_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1294 (.I0(n30681), .I1(n20_adj_3768), .I2(n16_adj_3732), 
            .I3(n30377), .O(n16246));
    defparam i10_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(\data_out_frame[14] [7]), .I1(n15630), 
            .I2(GND_net), .I3(GND_net), .O(n30435));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1296 (.I0(\data_out_frame[15] [0]), .I1(n15863), 
            .I2(\data_out_frame[14] [6]), .I3(n6_adj_3731), .O(n15541));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1297 (.I0(\data_out_frame[14] [6]), .I1(n30597), 
            .I2(n30333), .I3(n27179), .O(n31361));
    defparam i3_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1298 (.I0(\data_out_frame[16] [4]), .I1(n31361), 
            .I2(\data_out_frame[19] [0]), .I3(GND_net), .O(n26497));
    defparam i2_3_lut_adj_1298.LUT_INIT = 16'h6969;
    SB_LUT4 i13027_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [2]), 
            .I3(PWMLimit[18]), .O(n17414));
    defparam i13027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(n30585), .I1(n30315), .I2(\data_out_frame[6] [3]), 
            .I3(\data_out_frame[5] [7]), .O(n15630));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(\data_out_frame[18] [5]), .I1(n16042), 
            .I2(GND_net), .I3(GND_net), .O(n30568));
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n32567), .I3(n32566), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13028_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [3]), 
            .I3(PWMLimit[19]), .O(n17415));
    defparam i13028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1301 (.I0(n30764), .I1(n15054), .I2(n15630), 
            .I3(n26497), .O(n15_adj_3769));
    defparam i6_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1302 (.I0(n15_adj_3769), .I1(n16217), .I2(n14), 
            .I3(n30568), .O(n27001));
    defparam i8_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15766));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h6666;
    SB_LUT4 i1211_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1967));   // verilog/coms.v(69[16:27])
    defparam i1211_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1304 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[18] [4]), .I3(\data_out_frame[18] [3]), 
            .O(n30731));
    defparam i3_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1305 (.I0(\data_out_frame[17] [0]), .I1(n15532), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n30333));
    defparam i2_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n15760));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30501));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30743));
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30691));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1310 (.I0(n30559), .I1(n30691), .I2(\data_out_frame[13] [2]), 
            .I3(n30281), .O(n12_adj_3770));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1311 (.I0(\data_out_frame[7] [0]), .I1(n12_adj_3770), 
            .I2(n30749), .I3(\data_out_frame[6] [7]), .O(n16214));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30298));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i13029_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [4]), 
            .I3(PWMLimit[20]), .O(n17416));
    defparam i13029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1313 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [7]), 
            .I2(n30315), .I3(n6_adj_3730), .O(n1595));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1314 (.I0(n1595), .I1(n30687), .I2(n30276), .I3(GND_net), 
            .O(n30746));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30728));
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30752));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1317 (.I0(n30637), .I1(n30728), .I2(\data_out_frame[15] [5]), 
            .I3(n30562), .O(n12_adj_3771));
    defparam i5_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1318 (.I0(\data_out_frame[13] [3]), .I1(n12_adj_3771), 
            .I2(n30752), .I3(\data_out_frame[8] [5]), .O(n26362));
    defparam i6_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\data_out_frame[16] [0]), .I1(n26362), 
            .I2(GND_net), .I3(GND_net), .O(n30260));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(n15054), .I1(n30461), .I2(GND_net), 
            .I3(GND_net), .O(n27257));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1321 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3772));
    defparam i2_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i13030_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [5]), 
            .I3(PWMLimit[21]), .O(n17417));
    defparam i13030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1322 (.I0(n7_adj_3772), .I1(n15034), .I2(n27257), 
            .I3(n30260), .O(n26487));
    defparam i4_4_lut_adj_1322.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1323 (.I0(\data_out_frame[5] [3]), .I1(n30579), 
            .I2(\data_out_frame[12] [0]), .I3(n30254), .O(n18_adj_3773));   // verilog/coms.v(73[16:43])
    defparam i7_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3774));   // verilog/coms.v(73[16:43])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1324 (.I0(n1237), .I1(n18_adj_3773), .I2(\data_out_frame[14] [1]), 
            .I3(\data_out_frame[9] [6]), .O(n20_adj_3775));   // verilog/coms.v(73[16:43])
    defparam i9_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1325 (.I0(\data_out_frame[13] [7]), .I1(n20_adj_3775), 
            .I2(n16_adj_3774), .I3(\data_out_frame[5] [4]), .O(n16042));   // verilog/coms.v(73[16:43])
    defparam i10_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i13031_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [6]), 
            .I3(PWMLimit[22]), .O(n17418));
    defparam i13031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13032_3_lut_4_lut (.I0(n21292), .I1(n63_adj_3660), .I2(\data_in_frame[5] [7]), 
            .I3(PWMLimit[23]), .O(n17419));
    defparam i13032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12851_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n17238));
    defparam i12851_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12852_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n17239));
    defparam i12852_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12853_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n17240));
    defparam i12853_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1326 (.I0(n16042), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30350));
    defparam i1_2_lut_adj_1326.LUT_INIT = 16'h6666;
    SB_LUT4 i12854_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n17241));
    defparam i12854_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12855_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n17242));
    defparam i12855_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1327 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[10] [2]), 
            .I2(n30525), .I3(n30218), .O(n12_adj_3776));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1328 (.I0(\data_out_frame[9] [7]), .I1(n12_adj_3776), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[12] [3]), .O(n30224));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(n15863), .I1(n30224), .I2(GND_net), 
            .I3(GND_net), .O(n26562));
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1330 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [7]), 
            .I2(n30384), .I3(\data_out_frame[8] [7]), .O(n30684));
    defparam i3_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30318));
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3777));
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i12856_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n17243));
    defparam i12856_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1333 (.I0(n30551), .I1(n30318), .I2(n30684), 
            .I3(n6_adj_3777), .O(n30461));
    defparam i4_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1334 (.I0(n30254), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[15] [6]), .I3(\data_out_frame[16] [0]), 
            .O(n30787));
    defparam i3_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1335 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n30687));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30438));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15651));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30377));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1339 (.I0(n30377), .I1(\data_out_frame[6] [4]), 
            .I2(n15651), .I3(\data_out_frame[8] [5]), .O(n30617));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1340 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30276));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30749));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30719));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1343 (.I0(\data_out_frame[9] [1]), .I1(n30749), 
            .I2(n30276), .I3(\data_out_frame[9] [2]), .O(n30562));
    defparam i3_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30525));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30384));
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30465));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1347 (.I0(n16226), .I1(n30465), .I2(n16426), 
            .I3(\data_out_frame[14] [2]), .O(n30645));
    defparam i3_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1348 (.I0(n30444), .I1(n30522), .I2(\data_out_frame[14] [3]), 
            .I3(\data_out_frame[10] [1]), .O(n12_adj_3778));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1349 (.I0(\data_out_frame[12] [2]), .I1(n12_adj_3778), 
            .I2(n30579), .I3(\data_out_frame[12] [1]), .O(n16356));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1350 (.I0(n15704), .I1(n30519), .I2(n32127), 
            .I3(\data_in_frame[16] [6]), .O(n30417));
    defparam i1_2_lut_3_lut_4_lut_adj_1350.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30585));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1352 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30208));
    defparam i1_2_lut_adj_1352.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1353 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n30381));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(\data_out_frame[12] [5]), .I1(n15886), 
            .I2(GND_net), .I3(GND_net), .O(n30407));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1355 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[6] [0]), .I3(n6_adj_3729), .O(n15880));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i12857_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n17244));
    defparam i12857_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30305));
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1357 (.I0(n16335), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [3]), .I3(n30305), .O(n10_adj_3779));
    defparam i4_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1358 (.I0(\data_out_frame[8] [1]), .I1(n10_adj_3779), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n15886));
    defparam i5_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1359 (.I0(n15886), .I1(n30411), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n15863));
    defparam i2_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i12858_3_lut_4_lut (.I0(n10), .I1(n30168), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n17245));
    defparam i12858_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12843_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n17230));
    defparam i12843_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30250));
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i12844_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n17231));
    defparam i12844_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1361 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[9] [1]), .I3(GND_net), .O(n30281));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1362 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(n30208), .I3(n30381), .O(n14_adj_3780));
    defparam i6_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1363 (.I0(n1112), .I1(n1256), .I2(\data_out_frame[7] [2]), 
            .I3(\data_out_frame[5] [2]), .O(n13_adj_3781));
    defparam i5_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1364 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[11] [6]), .I3(\data_out_frame[10] [5]), 
            .O(n14_adj_3782));
    defparam i6_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1365 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[11] [7]), .I3(\data_out_frame[11] [2]), 
            .O(n13_adj_3783));
    defparam i5_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1366 (.I0(n13_adj_3781), .I1(n30585), .I2(n14_adj_3780), 
            .I3(GND_net), .O(n12_adj_3784));
    defparam i2_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i12845_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n17232));
    defparam i12845_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1367 (.I0(n30384), .I1(n12_adj_3784), .I2(n13_adj_3783), 
            .I3(n14_adj_3782), .O(n16_adj_3785));
    defparam i6_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1368 (.I0(n30525), .I1(n30465), .I2(n30562), 
            .I3(n30719), .O(n17_adj_3786));
    defparam i7_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1369 (.I0(n17_adj_3786), .I1(n30617), .I2(n16_adj_3785), 
            .I3(n30767), .O(n32150));
    defparam i9_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1370 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[15] [2]), 
            .I2(n30438), .I3(n18), .O(n30));
    defparam i13_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1371 (.I0(n15532), .I1(n30687), .I2(n30787), 
            .I3(n30461), .O(n28_adj_3787));
    defparam i11_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1372 (.I0(n30281), .I1(n27179), .I2(n16377), 
            .I3(\data_out_frame[15] [5]), .O(n29));
    defparam i12_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1373 (.I0(n30684), .I1(n30698), .I2(n32150), 
            .I3(n30350), .O(n27_adj_3788));
    defparam i10_4_lut_adj_1373.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1374 (.I0(n27_adj_3788), .I1(n29), .I2(n28_adj_3787), 
            .I3(n30), .O(n32152));
    defparam i16_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1375 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(n26487), .I3(n30434), .O(n54_adj_3789));
    defparam i23_4_lut_adj_1375.LUT_INIT = 16'h9669;
    SB_LUT4 i12846_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n17233));
    defparam i12846_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21_4_lut_adj_1376 (.I0(n30695), .I1(n30260), .I2(n30501), 
            .I3(\data_out_frame[19] [3]), .O(n52_adj_3790));
    defparam i21_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1377 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[11] [3]), .I3(n32152), .O(n53_adj_3791));
    defparam i22_4_lut_adj_1377.LUT_INIT = 16'h9669;
    SB_LUT4 i20_4_lut_adj_1378 (.I0(\data_out_frame[18] [2]), .I1(n30781), 
            .I2(\data_out_frame[19] [5]), .I3(n30746), .O(n51));
    defparam i20_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1379 (.I0(n30333), .I1(n30731), .I2(n1967), 
            .I3(\data_out_frame[9] [3]), .O(n48_adj_3792));
    defparam i17_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1380 (.I0(n30250), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[17] [6]), .I3(\data_out_frame[5] [1]), .O(n50_adj_3793));
    defparam i19_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1381 (.I0(n16048), .I1(n30770), .I2(\data_out_frame[19] [4]), 
            .I3(n30588), .O(n49));
    defparam i18_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n51), .I1(n53_adj_3791), .I2(n52_adj_3790), 
            .I3(n54_adj_3789), .O(n60));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1382 (.I0(n15766), .I1(n48_adj_3792), .I2(n30793), 
            .I3(\data_out_frame[13] [6]), .O(n55_adj_3794));
    defparam i24_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n55_adj_3794), .I1(n60), .I2(n49), .I3(n50_adj_3793), 
            .O(n27213));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1383 (.I0(\data_out_frame[16] [5]), .I1(n16356), 
            .I2(\data_out_frame[18] [7]), .I3(GND_net), .O(n30597));
    defparam i2_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 n36984_bdd_4_lut_4_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(n36984), .O(n36987));
    defparam n36984_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_LUT4 i6_4_lut_adj_1384 (.I0(n30392), .I1(\data_out_frame[16] [6]), 
            .I2(n26562), .I3(n27001), .O(n14_adj_3795));
    defparam i6_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1385 (.I0(\data_out_frame[20] [7]), .I1(n14_adj_3795), 
            .I2(n10_adj_3728), .I3(\data_out_frame[15] [1]), .O(n31499));
    defparam i7_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i12847_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n17234));
    defparam i12847_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30637));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30447));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i12848_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n17235));
    defparam i12848_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1388 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_1388.LUT_INIT = 16'h6666;
    SB_LUT4 i12849_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n17236));
    defparam i12849_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12850_3_lut_4_lut (.I0(n10), .I1(n30172), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n17237));
    defparam i12850_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1389 (.I0(\data_out_frame[7] [2]), .I1(n30793), 
            .I2(GND_net), .I3(GND_net), .O(n30681));
    defparam i1_2_lut_adj_1389.LUT_INIT = 16'h6666;
    SB_LUT4 i12995_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n17382));
    defparam i12995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1390 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30294));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1391 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n30365));
    defparam i2_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1392 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n31635));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1393 (.I0(\data_out_frame[11] [6]), .I1(n30294), 
            .I2(n31635), .I3(n15506), .O(n16226));
    defparam i3_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1394 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n30257));
    defparam i2_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1395 (.I0(n16226), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[13] [7]), .I3(n30365), .O(n30551));
    defparam i3_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i12996_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n17383));
    defparam i12996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1396 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16048));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1397 (.I0(n1237), .I1(n30551), .I2(n30257), .I3(\data_out_frame[13] [6]), 
            .O(n15034));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i500_2_lut (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1256));   // verilog/coms.v(83[17:28])
    defparam i500_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12997_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n17384));
    defparam i12997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1398 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30444));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1398.LUT_INIT = 16'h6666;
    SB_LUT4 i356_2_lut (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1112));   // verilog/coms.v(74[16:27])
    defparam i356_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1399 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16335));
    defparam i1_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1400 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(n1256), .I3(\data_out_frame[6] [0]), .O(n30218));
    defparam i3_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1401 (.I0(\data_out_frame[10] [2]), .I1(n30218), 
            .I2(n30522), .I3(\data_out_frame[5] [4]), .O(n30411));
    defparam i1_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i12998_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n17385));
    defparam i12998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12999_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n17386));
    defparam i12999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13000_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n17387));
    defparam i13000_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13001_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n17388));
    defparam i13001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1402 (.I0(\data_out_frame[5] [3]), .I1(n1112), 
            .I2(n30444), .I3(\data_out_frame[7] [6]), .O(n12_adj_3796));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1403 (.I0(\data_out_frame[5] [2]), .I1(n12_adj_3796), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[10] [0]), .O(n16426));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1404 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[12] [2]), 
            .I2(n16426), .I3(n30411), .O(n30767));
    defparam i3_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i13002_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30190), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n17389));
    defparam i13002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1405 (.I0(n15034), .I1(n16048), .I2(\data_out_frame[14] [0]), 
            .I3(\data_out_frame[18] [4]), .O(n30612));
    defparam i3_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i12987_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n17374));
    defparam i12987_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12988_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n17375));
    defparam i12988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\data_out_frame[16] [3]), .I1(n30434), 
            .I2(GND_net), .I3(GND_net), .O(n16217));
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'h9999;
    SB_LUT4 i12989_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n17376));
    defparam i12989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30371));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i2228_2_lut (.I0(n3915), .I1(\FRAME_MATCHER.state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n5782));
    defparam i2228_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12990_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n17377));
    defparam i12990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12991_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n17378));
    defparam i12991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_330_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3712));
    defparam select_330_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3711));
    defparam select_330_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3710));
    defparam select_330_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3709));
    defparam select_330_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3708));
    defparam select_330_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3707));
    defparam select_330_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3706));
    defparam select_330_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3705));
    defparam select_330_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3704));
    defparam select_330_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3703));
    defparam select_330_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3701));
    defparam select_330_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3699));
    defparam select_330_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3697));
    defparam select_330_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3695));
    defparam select_330_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3694));
    defparam select_330_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3693));
    defparam select_330_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3692));
    defparam select_330_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3691));
    defparam select_330_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3690));
    defparam select_330_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3689));
    defparam select_330_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3688));
    defparam select_330_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3687));
    defparam select_330_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3686));
    defparam select_330_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3685));
    defparam select_330_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3684));
    defparam select_330_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3683));
    defparam select_330_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12992_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n17379));
    defparam i12992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_330_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3682));
    defparam select_330_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3681));
    defparam select_330_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_330_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3680));
    defparam select_330_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12993_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n17380));
    defparam i12993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_330_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2430), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3679));
    defparam select_330_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12994_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30164), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n17381));
    defparam i12994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[17] [0]), .I1(n15541), 
            .I2(n15532), .I3(\data_out_frame[16] [6]), .O(n30669));
    defparam i1_2_lut_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1409 (.I0(n15880), .I1(\data_out_frame[12] [5]), 
            .I2(n15886), .I3(n15863), .O(n27179));
    defparam i1_2_lut_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1410 (.I0(n15880), .I1(\data_out_frame[12] [5]), 
            .I2(n15886), .I3(\data_out_frame[13] [0]), .O(n27173));
    defparam i1_2_lut_3_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i12979_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n17366));
    defparam i12979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12980_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n17367));
    defparam i12980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1411 (.I0(\data_out_frame[14] [4]), .I1(n30767), 
            .I2(n15863), .I3(n30224), .O(n15532));
    defparam i1_2_lut_3_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_3_lut_4_lut (.I0(\data_out_frame[16] [3]), .I1(n30434), 
            .I2(n30612), .I3(n30513), .O(n15_adj_3756));   // verilog/coms.v(69[16:27])
    defparam i4_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12981_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n17368));
    defparam i12981_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3675));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3674));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12982_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n17369));
    defparam i12982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12983_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n17370));
    defparam i12983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12984_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n17371));
    defparam i12984_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12985_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n17372));
    defparam i12985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12986_3_lut_4_lut (.I0(n10_adj_3552), .I1(n30168), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n17373));
    defparam i12986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12876_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n17263));
    defparam i12876_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12877_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n17264));
    defparam i12877_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12878_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n17265));
    defparam i12878_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12879_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n17266));
    defparam i12879_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12880_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n17267));
    defparam i12880_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12881_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n17268));
    defparam i12881_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12882_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n17269));
    defparam i12882_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12875_3_lut_4_lut (.I0(n10), .I1(n30187), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n17262));
    defparam i12875_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12883_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n17270));
    defparam i12883_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1412 (.I0(n15781), .I1(n27248), .I2(\data_in_frame[13] [4]), 
            .I3(GND_net), .O(n30340));
    defparam i1_2_lut_3_lut_adj_1412.LUT_INIT = 16'h6969;
    SB_LUT4 i12884_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n17271));
    defparam i12884_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12885_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n17272));
    defparam i12885_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12886_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n17273));
    defparam i12886_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12887_3_lut_4_lut (.I0(n10), .I1(n31262), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n17274));
    defparam i12887_3_lut_4_lut.LUT_INIT = 16'hfb40;
    uart_tx tx (.GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .tx_data({tx_data}), .tx_o(tx_o), .tx_enable(tx_enable), .\r_SM_Main_2__N_3259[0] (\r_SM_Main_2__N_3259[0] ), 
            .tx_active(tx_active)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.n16816(n16816), .r_Bit_Index({r_Bit_Index}), .clk32MHz(clk32MHz), 
            .n16819(n16819), .n29853(n29853), .rx_data_ready(rx_data_ready), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3185[2] (\r_SM_Main_2__N_3185[2] ), 
            .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .PIN_13_N_65(PIN_13_N_65), 
            .VCC_net(VCC_net), .n16600(n16600), .n16687(n16687), .n4573(n4573), 
            .n17013(n17013), .rx_data({rx_data}), .n16841(n16841), .n16840(n16840), 
            .n16839(n16839), .n16835(n16835), .n16825(n16825), .n16824(n16824), 
            .n16823(n16823), .n21347(n21347), .n4(n4), .n4_adj_1(n4_adj_4), 
            .n15244(n15244), .n15373(n15373), .n4_adj_2(n4_adj_5)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (GND_net, clk32MHz, VCC_net, tx_data, tx_o, tx_enable, 
            \r_SM_Main_2__N_3259[0] , tx_active) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input [7:0]tx_data;
    output tx_o;
    output tx_enable;
    input \r_SM_Main_2__N_3259[0] ;
    output tx_active;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [8:0]n312;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n24700, n24701, n24699, n24698, n24697, n17531;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n16813, n29897, n17478;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n16585, n23819, n24696, n13047;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n23902, n16606, n31428, n10, n5, n37002, n37005, n24703, 
        n24702, n29961, n29903, n15, n31835, n36891, n23926, n17, 
        n46, n4, n34339, n10_adj_3532, n36888;
    
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n24700), .O(n312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n24700), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n24701));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n24699), .O(n312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n24699), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n24700));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n24698), .O(n312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n24698), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n24699));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n24697), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17531));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n16813));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n29897));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n17478));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .E(n16585), 
            .D(n312[8]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .E(n16585), 
            .D(n312[7]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .E(n16585), 
            .D(n312[6]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .E(n16585), 
            .D(n312[5]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .E(n16585), 
            .D(n312[4]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .E(n16585), 
            .D(n312[3]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .E(n16585), 
            .D(n312[2]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .E(n16585), 
            .D(n312[1]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_4 (.CI(n24697), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n24698));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n24696), .O(n312[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n24696), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n24697));
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n312[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n24696));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(\r_SM_Main_2__N_3259[0] ), .O(n13047));   // verilog/uart_tx.v(31[16:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i31192_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(n23902), 
            .I3(r_SM_Main[2]), .O(n23819));   // verilog/uart_tx.v(31[16:25])
    defparam i31192_3_lut_4_lut.LUT_INIT = 16'h00f1;
    SB_LUT4 i19_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16585));
    defparam i19_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(n16585), 
            .D(n312[0]), .R(n23819));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i19621_4_lut (.I0(n16606), .I1(r_SM_Main[1]), .I2(r_Bit_Index[1]), 
            .I3(r_Bit_Index[0]), .O(n16813));   // verilog/uart_tx.v(31[16:25])
    defparam i19621_4_lut.LUT_INIT = 16'h58d0;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[2]), .O(n31428));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(n31428), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[8]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n23902));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/uart_tx.v(33[16:27])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n23902), .O(n16606));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i19603_4_lut (.I0(n16606), .I1(r_SM_Main[1]), .I2(r_Bit_Index[2]), 
            .I3(n5), .O(n17531));   // verilog/uart_tx.v(31[16:25])
    defparam i19603_4_lut.LUT_INIT = 16'h58d0;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n37002));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37002_bdd_4_lut (.I0(n37002), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n37005));
    defparam n37002_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_3_lut (.I0(n16606), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29897));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13047), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n24703), .O(n312[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n24702), .O(n312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n29961));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n29903));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n15));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_9 (.CI(n24702), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n24703));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n24701), .O(n312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n31835));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_8 (.CI(n24701), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n24702));
    SB_LUT4 i19611_3_lut (.I0(n37005), .I1(n36891), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n23926));   // verilog/uart_tx.v(33[16:27])
    defparam i19611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut (.I0(n23926), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(133[8:12])
    defparam i33_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i32_3_lut (.I0(n17), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n15));   // verilog/TinyFPGA_B.v(133[8:12])
    defparam i32_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_2_lut_adj_860 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3259[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n46));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h4444;
    SB_LUT4 i12_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(n46), .I3(n4), 
            .O(n29903));   // verilog/uart_tx.v(31[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i29298_2_lut (.I0(n23902), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34339));   // verilog/uart_tx.v(33[16:27])
    defparam i29298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24_4_lut (.I0(\r_SM_Main_2__N_3259[0] ), .I1(n34339), .I2(r_SM_Main[1]), 
            .I3(n5), .O(n10_adj_3532));   // verilog/uart_tx.v(33[16:27])
    defparam i24_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n23902), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n17478));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0078;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_31344 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n36888));
    defparam r_Bit_Index_0__bdd_4_lut_31344.LUT_INIT = 16'he4aa;
    SB_LUT4 n36888_bdd_4_lut (.I0(n36888), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n36891));
    defparam n36888_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(n23902), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i3_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(n23902), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main[1]), .O(n31835));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_3_lut_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(n10_adj_3532), .I2(n23902), 
            .I3(r_SM_Main[0]), .O(n29961));   // verilog/uart_tx.v(33[16:27])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0544;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n16816, r_Bit_Index, clk32MHz, n16819, n29853, rx_data_ready, 
            r_SM_Main, \r_SM_Main_2__N_3185[2] , GND_net, r_Rx_Data, 
            PIN_13_N_65, VCC_net, n16600, n16687, n4573, n17013, 
            rx_data, n16841, n16840, n16839, n16835, n16825, n16824, 
            n16823, n21347, n4, n4_adj_1, n15244, n15373, n4_adj_2) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n16816;
    output [2:0]r_Bit_Index;
    input clk32MHz;
    input n16819;
    input n29853;
    output rx_data_ready;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3185[2] ;
    input GND_net;
    output r_Rx_Data;
    input PIN_13_N_65;
    input VCC_net;
    output n16600;
    output n16687;
    output n4573;
    input n17013;
    output [7:0]rx_data;
    input n16841;
    input n16840;
    input n16839;
    input n16835;
    input n16825;
    input n16824;
    input n16823;
    output n21347;
    output n4;
    output n4_adj_1;
    output n15244;
    output n15373;
    output n4_adj_2;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n16865;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n16871, n16874, n17509, n16883, n17507, n16929, n16940, 
        n17493, n17468, n31843, n34160, n23242, n34285, n24695;
    wire [31:0]n194;
    
    wire n24694, r_Rx_Data_R, n34277, n24693, n34276, n24692, n24691, 
        n24690, n24689, n6, n251, n30091, n4_c, n244, n4_adj_3525;
    wire [2:0]r_SM_Main_2__N_3188;
    
    wire n6_adj_3526, n223_adj_3527, n245, n266, n6_adj_3528, n16908, 
        n15249, n37035, n37032, n34263;
    
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n16816));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n16819));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n16865));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n16871));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n16874));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n17509));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n16883));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n17507));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n16929));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n16940));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17493));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n29853));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n17468));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3185[2] ), 
            .R(n31843));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i25215_4_lut (.I0(r_SM_Main[2]), .I1(n34160), .I2(\r_SM_Main_2__N_3185[2] ), 
            .I3(r_SM_Main[1]), .O(n23242));   // verilog/uart_rx.v(36[17:26])
    defparam i25215_4_lut.LUT_INIT = 16'hafee;
    SB_LUT4 add_62_9_lut (.I0(n23242), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n24695), .O(n34285)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n24694), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_65));   // verilog/uart_rx.v(41[10] 45[8])
    SB_CARRY add_62_8 (.CI(n24694), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n24695));
    SB_LUT4 add_62_7_lut (.I0(n23242), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n24693), .O(n34277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n24693), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n24694));
    SB_LUT4 add_62_6_lut (.I0(n23242), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n24692), .O(n34276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n24692), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n24693));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n24691), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n24691), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n24692));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n24690), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n24690), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n24691));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n24689), .O(n194[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n24689), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n24690));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n24689));
    SB_LUT4 i2_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n31843));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_adj_848 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n6));
    defparam i2_3_lut_adj_848.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_849 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(GND_net), .O(n251));
    defparam i2_3_lut_adj_849.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[5]), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[4]), .O(n30091));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[3]), .I1(n30091), .I2(n251), .I3(GND_net), 
            .O(\r_SM_Main_2__N_3185[2] ));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3185[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n16600));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i12338_3_lut (.I0(n16600), .I1(n6), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n16687));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12338_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1222_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4573));   // verilog/uart_rx.v(102[36:51])
    defparam i1222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_850 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(\r_SM_Main_2__N_3185[2] ), 
            .I3(GND_net), .O(n244));   // verilog/uart_rx.v(36[17:26])
    defparam i1_3_lut_adj_850.LUT_INIT = 16'hecec;
    SB_LUT4 i19070_4_lut (.I0(n4_adj_3525), .I1(n244), .I2(r_SM_Main[1]), 
            .I3(n4_c), .O(n17468));   // verilog/uart_rx.v(36[17:26])
    defparam i19070_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_3188[0]), .O(n6_adj_3526));
    defparam i1_4_lut.LUT_INIT = 16'h0501;
    SB_LUT4 i14222_4_lut (.I0(n16687), .I1(n6_adj_3526), .I2(n16600), 
            .I3(r_Bit_Index[0]), .O(n17493));
    defparam i14222_4_lut.LUT_INIT = 16'h0530;
    SB_LUT4 i29367_4_lut (.I0(r_Clock_Count[0]), .I1(n23242), .I2(n194[0]), 
            .I3(n223_adj_3527), .O(n16929));
    defparam i29367_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_851 (.I0(n245), .I1(r_Rx_Data), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3525));   // verilog/uart_rx.v(41[10] 45[8])
    defparam i1_2_lut_adj_851.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_852 (.I0(n30091), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(GND_net), .O(n266));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_852.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_853 (.I0(n266), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[0]), .O(n245));
    defparam i3_4_lut_adj_853.LUT_INIT = 16'hbfff;
    SB_LUT4 i2_2_lut (.I0(n245), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_3528));   // verilog/uart_rx.v(36[17:26])
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_854 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n6_adj_3528), 
            .I3(r_SM_Main[0]), .O(n223_adj_3527));   // verilog/uart_rx.v(36[17:26])
    defparam i1_4_lut_adj_854.LUT_INIT = 16'h3233;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n17013));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n16908));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n16841));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n16840));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n16839));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n16835));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n16825));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n16824));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n16823));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i18956_3_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n34276), 
            .I3(r_Clock_Count[4]), .O(n16874));
    defparam i18956_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_4_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n194[2]), 
            .I3(r_Clock_Count[2]), .O(n16865));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hc480;
    SB_LUT4 i12484_4_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n194[3]), 
            .I3(r_Clock_Count[3]), .O(n16871));
    defparam i12484_4_lut_4_lut.LUT_INIT = 16'hc480;
    SB_LUT4 i12553_4_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n194[1]), 
            .I3(r_Clock_Count[1]), .O(n16940));
    defparam i12553_4_lut_4_lut.LUT_INIT = 16'hc480;
    SB_LUT4 i1_4_lut_4_lut_adj_855 (.I0(n223_adj_3527), .I1(n23242), .I2(n194[6]), 
            .I3(r_Clock_Count[6]), .O(n16883));
    defparam i1_4_lut_4_lut_adj_855.LUT_INIT = 16'hc480;
    SB_LUT4 i16982_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n21347));
    defparam i16982_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18988_3_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n34277), 
            .I3(r_Clock_Count[5]), .O(n17509));
    defparam i18988_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 equal_130_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_130_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_132_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_132_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i19020_3_lut_4_lut (.I0(n223_adj_3527), .I1(n23242), .I2(n34285), 
            .I3(r_Clock_Count[7]), .O(n17507));
    defparam i19020_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_adj_856 (.I0(r_Bit_Index[0]), .I1(n15249), .I2(GND_net), 
            .I3(GND_net), .O(n15244));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_856.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_857 (.I0(r_SM_Main[2]), .I1(n37035), .I2(GND_net), 
            .I3(GND_net), .O(n16908));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut_adj_858 (.I0(r_SM_Main[0]), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(\r_SM_Main_2__N_3185[2] ), .O(n15249));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i3_4_lut_adj_858.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_859 (.I0(r_Bit_Index[0]), .I1(n15249), .I2(GND_net), 
            .I3(GND_net), .O(n15373));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_859.LUT_INIT = 16'heeee;
    SB_LUT4 equal_134_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_134_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28978_2_lut_3_lut (.I0(n245), .I1(r_Rx_Data), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n34160));   // verilog/uart_rx.v(36[17:26])
    defparam i28978_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(\r_SM_Main_2__N_3185[2] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(r_Bit_Index[0]), .O(r_SM_Main_2__N_3188[0]));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(\r_SM_Main_2__N_3185[2] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main_2__N_3188[0]), .I3(r_SM_Main[0]), .O(n37032));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 n37032_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n34263), 
            .I3(n37032), .O(n37035));   // verilog/uart_rx.v(30[17:26])
    defparam n37032_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i28908_2_lut_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(n266), .O(n34263));
    defparam i28908_2_lut_4_lut.LUT_INIT = 16'hff7f;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n17466, encoder1_position, clk32MHz, 
            n17465, n17464, n17463, n17462, n17461, n17460, n17459, 
            n17458, n17457, n17456, n17455, n17454, n17453, n17452, 
            n17451, n17450, n17449, n17448, n17447, n17446, n17445, 
            n17444, data_o, GND_net, n2571, count_enable, n16906, 
            n17479, reg_B, n31841, PIN_7_c_1, PIN_6_c_0, n16918) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17466;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n17465;
    input n17464;
    input n17463;
    input n17462;
    input n17461;
    input n17460;
    input n17459;
    input n17458;
    input n17457;
    input n17456;
    input n17455;
    input n17454;
    input n17453;
    input n17452;
    input n17451;
    input n17450;
    input n17449;
    input n17448;
    input n17447;
    input n17446;
    input n17445;
    input n17444;
    output [1:0]data_o;
    input GND_net;
    output [23:0]n2571;
    output count_enable;
    input n16906;
    input n17479;
    output [1:0]reg_B;
    output n31841;
    input PIN_7_c_1;
    input PIN_6_c_0;
    input n16918;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, count_direction, n2561, n24850, n24849, 
        n24848, n24847, n24846, n24845, n24844, n24843, n24842, 
        n24841, n24840, n24839, n24838, n24837, n24836, n24835, 
        n24834, n24833, n24832, n24831, n24830, n24829, n24828, 
        n24827;
    
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n17466));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n17465));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n17464));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n17463));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n17462));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n17461));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n17460));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n17459));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n17458));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n17457));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n17456));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n17455));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n17454));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n17453));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n17452));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n17451));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n17450));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n17449));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n17448));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n17447));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n17446));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n17445));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n17444));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_586_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2561), 
            .I3(n24850), .O(n2571[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_586_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2561), 
            .I3(n24849), .O(n2571[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_24 (.CI(n24849), .I0(encoder1_position[22]), .I1(n2561), 
            .CO(n24850));
    SB_LUT4 add_586_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2561), 
            .I3(n24848), .O(n2571[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_23 (.CI(n24848), .I0(encoder1_position[21]), .I1(n2561), 
            .CO(n24849));
    SB_LUT4 add_586_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2561), 
            .I3(n24847), .O(n2571[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_22 (.CI(n24847), .I0(encoder1_position[20]), .I1(n2561), 
            .CO(n24848));
    SB_LUT4 add_586_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2561), 
            .I3(n24846), .O(n2571[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_21 (.CI(n24846), .I0(encoder1_position[19]), .I1(n2561), 
            .CO(n24847));
    SB_LUT4 add_586_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2561), 
            .I3(n24845), .O(n2571[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_20 (.CI(n24845), .I0(encoder1_position[18]), .I1(n2561), 
            .CO(n24846));
    SB_LUT4 add_586_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2561), 
            .I3(n24844), .O(n2571[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_19 (.CI(n24844), .I0(encoder1_position[17]), .I1(n2561), 
            .CO(n24845));
    SB_LUT4 add_586_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2561), 
            .I3(n24843), .O(n2571[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_18 (.CI(n24843), .I0(encoder1_position[16]), .I1(n2561), 
            .CO(n24844));
    SB_LUT4 add_586_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2561), 
            .I3(n24842), .O(n2571[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_17 (.CI(n24842), .I0(encoder1_position[15]), .I1(n2561), 
            .CO(n24843));
    SB_LUT4 add_586_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2561), 
            .I3(n24841), .O(n2571[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_16 (.CI(n24841), .I0(encoder1_position[14]), .I1(n2561), 
            .CO(n24842));
    SB_LUT4 add_586_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2561), 
            .I3(n24840), .O(n2571[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_15 (.CI(n24840), .I0(encoder1_position[13]), .I1(n2561), 
            .CO(n24841));
    SB_LUT4 add_586_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2561), 
            .I3(n24839), .O(n2571[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_14 (.CI(n24839), .I0(encoder1_position[12]), .I1(n2561), 
            .CO(n24840));
    SB_LUT4 add_586_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2561), 
            .I3(n24838), .O(n2571[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_13 (.CI(n24838), .I0(encoder1_position[11]), .I1(n2561), 
            .CO(n24839));
    SB_LUT4 add_586_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2561), 
            .I3(n24837), .O(n2571[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_12 (.CI(n24837), .I0(encoder1_position[10]), .I1(n2561), 
            .CO(n24838));
    SB_LUT4 add_586_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2561), 
            .I3(n24836), .O(n2571[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_11 (.CI(n24836), .I0(encoder1_position[9]), .I1(n2561), 
            .CO(n24837));
    SB_LUT4 add_586_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2561), 
            .I3(n24835), .O(n2571[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_10 (.CI(n24835), .I0(encoder1_position[8]), .I1(n2561), 
            .CO(n24836));
    SB_LUT4 add_586_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2561), 
            .I3(n24834), .O(n2571[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_9 (.CI(n24834), .I0(encoder1_position[7]), .I1(n2561), 
            .CO(n24835));
    SB_LUT4 add_586_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2561), 
            .I3(n24833), .O(n2571[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_8 (.CI(n24833), .I0(encoder1_position[6]), .I1(n2561), 
            .CO(n24834));
    SB_LUT4 add_586_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2561), 
            .I3(n24832), .O(n2571[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_7 (.CI(n24832), .I0(encoder1_position[5]), .I1(n2561), 
            .CO(n24833));
    SB_LUT4 add_586_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2561), 
            .I3(n24831), .O(n2571[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_586_6 (.CI(n24831), .I0(encoder1_position[4]), .I1(n2561), 
            .CO(n24832));
    SB_LUT4 add_586_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2561), 
            .I3(n24830), .O(n2571[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_5 (.CI(n24830), .I0(encoder1_position[3]), .I1(n2561), 
            .CO(n24831));
    SB_LUT4 add_586_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2561), 
            .I3(n24829), .O(n2571[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_4 (.CI(n24829), .I0(encoder1_position[2]), .I1(n2561), 
            .CO(n24830));
    SB_LUT4 add_586_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2561), 
            .I3(n24828), .O(n2571[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_3 (.CI(n24828), .I0(encoder1_position[1]), .I1(n2561), 
            .CO(n24829));
    SB_LUT4 add_586_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n24827), .O(n2571[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_586_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_586_2 (.CI(n24827), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n24828));
    SB_CARRY add_586_1 (.CI(GND_net), .I0(n2561), .I1(n2561), .CO(n24827));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n16906));   // quad.v(35[10] 41[6])
    SB_LUT4 i888_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2561));   // quad.v(37[5] 40[8])
    defparam i888_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n17479(n17479), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .GND_net(GND_net), .n31841(n31841), .PIN_7_c_1(PIN_7_c_1), 
            .PIN_6_c_0(PIN_6_c_0), .n16918(n16918)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n17479, data_o, clk32MHz, reg_B, GND_net, 
            n31841, PIN_7_c_1, PIN_6_c_0, n16918) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n17479;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n31841;
    input PIN_7_c_1;
    input PIN_6_c_0;
    input n16918;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3420;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17479));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n31841), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i20126_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20126_1_lut.LUT_INIT = 16'h5555;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_7_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1132__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n31841));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_6_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1132__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1132__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16918));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i20135_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20135_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i20128_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20128_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n17442, encoder0_position, clk32MHz, 
            n17441, n17440, n17439, n17438, n17437, n17436, n17435, 
            n17434, n17433, n17432, n17431, n17430, n17429, n17428, 
            n17427, n17426, n17425, n17424, n17423, n17422, n17421, 
            n17420, data_o, n2621, GND_net, count_enable, n16904, 
            n17467, reg_B, n31114, PIN_2_c_1, PIN_1_c_0, n16907) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17442;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n17441;
    input n17440;
    input n17439;
    input n17438;
    input n17437;
    input n17436;
    input n17435;
    input n17434;
    input n17433;
    input n17432;
    input n17431;
    input n17430;
    input n17429;
    input n17428;
    input n17427;
    input n17426;
    input n17425;
    input n17424;
    input n17423;
    input n17422;
    input n17421;
    input n17420;
    output [1:0]data_o;
    output [23:0]n2621;
    input GND_net;
    output count_enable;
    input n16904;
    input n17467;
    output [1:0]reg_B;
    output n31114;
    input PIN_2_c_1;
    input PIN_1_c_0;
    input n16907;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2617, n24727, n24726, n24725, n24724, 
        n24723, n24722, n24721, n24720, n24719, n24718, n24717, 
        n24716, n24715, n24714, n24713, n24712, n24711, n24710, 
        n24709, n24708, n24707, n24706, n24705, count_direction, 
        n24704;
    
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n17442));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n17441));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n17440));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n17439));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n17438));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n17437));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n17436));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n17435));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n17434));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n17433));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n17432));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n17431));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n17430));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n17429));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n17428));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n17427));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n17426));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n17425));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n17424));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n17423));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n17422));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n17421));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n17420));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_612_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2617), 
            .I3(n24727), .O(n2621[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_612_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2617), 
            .I3(n24726), .O(n2621[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_24 (.CI(n24726), .I0(encoder0_position[22]), .I1(n2617), 
            .CO(n24727));
    SB_LUT4 add_612_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2617), 
            .I3(n24725), .O(n2621[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_23 (.CI(n24725), .I0(encoder0_position[21]), .I1(n2617), 
            .CO(n24726));
    SB_LUT4 add_612_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2617), 
            .I3(n24724), .O(n2621[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_22 (.CI(n24724), .I0(encoder0_position[20]), .I1(n2617), 
            .CO(n24725));
    SB_LUT4 add_612_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2617), 
            .I3(n24723), .O(n2621[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_21 (.CI(n24723), .I0(encoder0_position[19]), .I1(n2617), 
            .CO(n24724));
    SB_LUT4 add_612_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2617), 
            .I3(n24722), .O(n2621[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_20 (.CI(n24722), .I0(encoder0_position[18]), .I1(n2617), 
            .CO(n24723));
    SB_LUT4 add_612_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2617), 
            .I3(n24721), .O(n2621[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_19 (.CI(n24721), .I0(encoder0_position[17]), .I1(n2617), 
            .CO(n24722));
    SB_LUT4 add_612_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2617), 
            .I3(n24720), .O(n2621[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_18 (.CI(n24720), .I0(encoder0_position[16]), .I1(n2617), 
            .CO(n24721));
    SB_LUT4 add_612_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2617), 
            .I3(n24719), .O(n2621[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_17 (.CI(n24719), .I0(encoder0_position[15]), .I1(n2617), 
            .CO(n24720));
    SB_LUT4 add_612_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2617), 
            .I3(n24718), .O(n2621[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_16 (.CI(n24718), .I0(encoder0_position[14]), .I1(n2617), 
            .CO(n24719));
    SB_LUT4 add_612_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2617), 
            .I3(n24717), .O(n2621[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_15 (.CI(n24717), .I0(encoder0_position[13]), .I1(n2617), 
            .CO(n24718));
    SB_LUT4 add_612_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2617), 
            .I3(n24716), .O(n2621[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_14 (.CI(n24716), .I0(encoder0_position[12]), .I1(n2617), 
            .CO(n24717));
    SB_LUT4 add_612_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2617), 
            .I3(n24715), .O(n2621[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_612_13 (.CI(n24715), .I0(encoder0_position[11]), .I1(n2617), 
            .CO(n24716));
    SB_LUT4 add_612_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2617), 
            .I3(n24714), .O(n2621[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_12 (.CI(n24714), .I0(encoder0_position[10]), .I1(n2617), 
            .CO(n24715));
    SB_LUT4 add_612_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2617), 
            .I3(n24713), .O(n2621[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_11 (.CI(n24713), .I0(encoder0_position[9]), .I1(n2617), 
            .CO(n24714));
    SB_LUT4 add_612_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2617), 
            .I3(n24712), .O(n2621[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_10 (.CI(n24712), .I0(encoder0_position[8]), .I1(n2617), 
            .CO(n24713));
    SB_LUT4 add_612_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2617), 
            .I3(n24711), .O(n2621[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_9 (.CI(n24711), .I0(encoder0_position[7]), .I1(n2617), 
            .CO(n24712));
    SB_LUT4 add_612_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2617), 
            .I3(n24710), .O(n2621[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_8 (.CI(n24710), .I0(encoder0_position[6]), .I1(n2617), 
            .CO(n24711));
    SB_LUT4 add_612_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2617), 
            .I3(n24709), .O(n2621[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_7 (.CI(n24709), .I0(encoder0_position[5]), .I1(n2617), 
            .CO(n24710));
    SB_LUT4 add_612_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2617), 
            .I3(n24708), .O(n2621[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_6 (.CI(n24708), .I0(encoder0_position[4]), .I1(n2617), 
            .CO(n24709));
    SB_LUT4 add_612_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2617), 
            .I3(n24707), .O(n2621[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_5 (.CI(n24707), .I0(encoder0_position[3]), .I1(n2617), 
            .CO(n24708));
    SB_LUT4 add_612_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2617), 
            .I3(n24706), .O(n2621[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_4 (.CI(n24706), .I0(encoder0_position[2]), .I1(n2617), 
            .CO(n24707));
    SB_LUT4 add_612_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2617), 
            .I3(n24705), .O(n2621[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_3 (.CI(n24705), .I0(encoder0_position[1]), .I1(n2617), 
            .CO(n24706));
    SB_LUT4 add_612_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n24704), .O(n2621[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_612_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_612_2 (.CI(n24704), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n24705));
    SB_CARRY add_612_1 (.CI(GND_net), .I0(n2617), .I1(n2617), .CO(n24704));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n16904));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i887_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2617));   // quad.v(37[5] 40[8])
    defparam i887_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n17467(n17467), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .GND_net(GND_net), .n31114(n31114), 
            .PIN_2_c_1(PIN_2_c_1), .PIN_1_c_0(PIN_1_c_0), .n16907(n16907)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n17467, data_o, clk32MHz, reg_B, GND_net, 
            n31114, PIN_2_c_1, PIN_1_c_0, n16907) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n17467;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n31114;
    input PIN_2_c_1;
    input PIN_1_c_0;
    input n16907;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3420;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17467));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n31114), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i20104_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20104_1_lut.LUT_INIT = 16'h5555;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_2_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1131__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n31114));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_1_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1131__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1131__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3420));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16907));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i20113_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20113_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i20106_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20106_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (pwm_setpoint, \half_duty_new[0] , 
            CLK_c, PIN_19_c_0, GND_net, VCC_net, n925, \half_duty[0][1] , 
            n17487, \half_duty[0][7] , n17486, \half_duty[0][6] , n17485, 
            \half_duty[0][5] , n17484, \half_duty[0][4] , n17483, \half_duty[0][3] , 
            n17482, \half_duty[0][2] , n17481, \half_duty_new[7] , \half_duty_new[6] , 
            \half_duty_new[5] , \half_duty_new[4] , \half_duty_new[3] , 
            \half_duty_new[2] , \half_duty_new[1] , \half_duty[0][0] , 
            n16936) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input [22:0]pwm_setpoint;
    output \half_duty_new[0] ;
    input CLK_c;
    output PIN_19_c_0;
    input GND_net;
    input VCC_net;
    output n925;
    output \half_duty[0][1] ;
    input n17487;
    output \half_duty[0][7] ;
    input n17486;
    output \half_duty[0][6] ;
    input n17485;
    output \half_duty[0][5] ;
    input n17484;
    output \half_duty[0][4] ;
    input n17483;
    output \half_duty[0][3] ;
    input n17482;
    output \half_duty[0][2] ;
    input n17481;
    output \half_duty_new[7] ;
    output \half_duty_new[6] ;
    output \half_duty_new[5] ;
    output \half_duty_new[4] ;
    output \half_duty_new[3] ;
    output \half_duty_new[2] ;
    output \half_duty_new[1] ;
    output \half_duty[0][0] ;
    input n16936;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n24903;
    wire [22:0]n5538;
    
    wire n24904, n24902, n24901, n24900, n24899, n24898, n24897, 
        n24896, n24895;
    wire [9:0]half_duty_new_9__N_600;
    
    wire pwm_out_0__N_518, n16531, n24894, n24893, n24892, n24891, 
        n24890, n24889, n24888, n10, n24647;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n24887, n24648, n9, n24646;
    wire [10:0]n49;
    
    wire pause_counter_0__N_548, n24886;
    wire [10:0]pwm_out_0__N_523;
    
    wire n24885, n24884, n8, n24645, n24883, n24882, n7, n24644, 
        n24881, n6, n24643, n5, n24642, n5_adj_3522, n20, n16, 
        n24880, n4, n24641, n24879, n24878, n24877, n24876, n24875, 
        n3, n24640, n24874, n2, n24639, n1, n30927, pause_counter_0, 
        n24649, pwm_out_0__N_522, n20_adj_3523, n19, n6_adj_3524, 
        n32443, n32513, n22, n21, n14, n12, n13, n25518, n25517, 
        n25516, n25515, n25514, n25513, n25512, n25511, n25510, 
        n25509, n24916, n24915, n24914, n24913, n24912, n24911, 
        n24910, n24909, n24908, n24907, n24906, n24905;
    
    SB_CARRY add_2006_11 (.CI(n24903), .I0(n5538[9]), .I1(pwm_setpoint[9]), 
            .CO(n24904));
    SB_CARRY add_2006_10 (.CI(n24902), .I0(n5538[8]), .I1(pwm_setpoint[8]), 
            .CO(n24903));
    SB_CARRY add_2006_9 (.CI(n24901), .I0(n5538[7]), .I1(pwm_setpoint[7]), 
            .CO(n24902));
    SB_CARRY add_2006_8 (.CI(n24900), .I0(n5538[6]), .I1(pwm_setpoint[6]), 
            .CO(n24901));
    SB_CARRY add_2006_7 (.CI(n24899), .I0(n5538[5]), .I1(pwm_setpoint[5]), 
            .CO(n24900));
    SB_CARRY add_2006_6 (.CI(n24898), .I0(n5538[4]), .I1(pwm_setpoint[4]), 
            .CO(n24899));
    SB_CARRY add_2006_5 (.CI(n24897), .I0(n5538[3]), .I1(pwm_setpoint[3]), 
            .CO(n24898));
    SB_CARRY add_2006_4 (.CI(n24896), .I0(n5538[2]), .I1(pwm_setpoint[2]), 
            .CO(n24897));
    SB_CARRY add_2006_3 (.CI(n24895), .I0(n5538[1]), .I1(pwm_setpoint[1]), 
            .CO(n24896));
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_600[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n16531), .D(pwm_out_0__N_518));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2006_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n24895));
    SB_LUT4 add_2014_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n24894), .O(n5538[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2014_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n24893), .O(n5538[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_22 (.CI(n24893), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n24894));
    SB_LUT4 add_2014_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n24892), .O(n5538[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_21 (.CI(n24892), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n24893));
    SB_LUT4 add_2014_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n24891), .O(n5538[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_20 (.CI(n24891), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n24892));
    SB_LUT4 add_2014_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n24890), .O(n5538[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_19 (.CI(n24890), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n24891));
    SB_LUT4 add_2014_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n24889), .O(n5538[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_18 (.CI(n24889), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n24890));
    SB_LUT4 add_2014_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n24888), .O(n5538[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_19_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n24647), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2014_17 (.CI(n24888), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n24889));
    SB_LUT4 add_2014_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n24887), .O(n5538[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_19_11 (.CI(n24647), .I0(VCC_net), .I1(VCC_net), 
            .CO(n24648));
    SB_LUT4 pwm_out_0__I_19_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n24646), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2014_16 (.CI(n24887), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n24888));
    SB_CARRY pwm_out_0__I_19_10 (.CI(n24646), .I0(GND_net), .I1(VCC_net), 
            .CO(n24647));
    SB_DFFESR count_0__1130__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[10]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[9]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[8]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[7]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[6]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 add_2014_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n24886), .O(n5538[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2014_15 (.CI(n24886), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n24887));
    SB_DFFESR count_0__1130__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[5]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 add_2014_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n24885), .O(n5538[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_14 (.CI(n24885), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n24886));
    SB_LUT4 add_2014_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n24884), .O(n5538[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1130__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[4]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n17487));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n17486));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0][5] ), .C(CLK_c), .D(n17485));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n17484));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n17483));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n17482));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n17481));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1130__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[3]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[2]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[1]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1130__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_548), 
            .D(n49[0]), .R(n925));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_2014_13 (.CI(n24884), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n24885));
    SB_LUT4 pwm_out_0__I_19_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_523[7]), 
            .I3(n24645), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_2014_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n24883), .O(n5538[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2014_12 (.CI(n24883), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n24884));
    SB_LUT4 add_2014_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n24882), .O(n5538[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_11 (.CI(n24882), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n24883));
    SB_CARRY pwm_out_0__I_19_9 (.CI(n24645), .I0(GND_net), .I1(pwm_out_0__N_523[7]), 
            .CO(n24646));
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_out_0__I_19_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_523[6]), 
            .I3(n24644), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_19_8 (.CI(n24644), .I0(VCC_net), .I1(pwm_out_0__N_523[6]), 
            .CO(n24645));
    SB_LUT4 add_2014_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n24881), .O(n5538[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_19_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_523[5]), 
            .I3(n24643), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_19_7 (.CI(n24643), .I0(GND_net), .I1(pwm_out_0__N_523[5]), 
            .CO(n24644));
    SB_LUT4 pwm_out_0__I_19_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_523[4]), 
            .I3(n24642), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 half_duty_0__9__I_0_47_i5_2_lut (.I0(\half_duty[0][4] ), .I1(\count[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3522));   // vhdl/pwm.vhd(80[8:31])
    defparam half_duty_0__9__I_0_47_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut (.I0(n5_adj_3522), .I1(n20), .I2(n16), .I3(\count[0] [10]), 
            .O(pwm_out_0__N_518));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY pwm_out_0__I_19_6 (.CI(n24642), .I0(GND_net), .I1(pwm_out_0__N_523[4]), 
            .CO(n24643));
    SB_CARRY add_2014_10 (.CI(n24881), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n24882));
    SB_LUT4 add_2014_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n24880), .O(n5538[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_19_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_523[3]), 
            .I3(n24641), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2014_9 (.CI(n24880), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n24881));
    SB_LUT4 add_2014_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n24879), .O(n5538[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_19_5 (.CI(n24641), .I0(GND_net), .I1(pwm_out_0__N_523[3]), 
            .CO(n24642));
    SB_CARRY add_2014_8 (.CI(n24879), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n24880));
    SB_LUT4 add_2014_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n24878), .O(n5538[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_7 (.CI(n24878), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n24879));
    SB_LUT4 add_2014_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n24877), .O(n5538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_6 (.CI(n24877), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n24878));
    SB_LUT4 add_2014_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n24876), .O(n5538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_5 (.CI(n24876), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n24877));
    SB_LUT4 add_2014_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n24875), .O(n5538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_19_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_523[2]), 
            .I3(n24640), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2014_4 (.CI(n24875), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n24876));
    SB_LUT4 add_2014_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n24874), .O(n5538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_19_4 (.CI(n24640), .I0(GND_net), .I1(pwm_out_0__N_523[2]), 
            .CO(n24641));
    SB_CARRY add_2014_3 (.CI(n24874), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n24875));
    SB_LUT4 add_2014_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2014_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2014_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n24874));
    SB_LUT4 pwm_out_0__I_19_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_523[1]), 
            .I3(n24639), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_19_3 (.CI(n24639), .I0(GND_net), .I1(pwm_out_0__N_523[1]), 
            .CO(n24640));
    SB_LUT4 pwm_out_0__I_19_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_523[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_19_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_19_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_523[0]), 
            .CO(n24639));
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0][5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i7_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[6]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n30927));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_600[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_600[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(\half_duty_new[5] ), .C(CLK_c), .D(half_duty_new_9__N_600[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_600[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_600[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_600[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_600[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_19_12 (.CI(n24648), .I0(VCC_net), .I1(VCC_net), 
            .CO(n24649));
    SB_CARRY pwm_out_0__I_19_13 (.CI(n24649), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_522));
    SB_LUT4 i8_4_lut (.I0(\count[0] [6]), .I1(\count[0] [0]), .I2(\count[0] [10]), 
            .I3(\count[0] [4]), .O(n20_adj_3523));
    defparam i8_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i7_4_lut (.I0(pause_counter_0), .I1(\count[0] [9]), .I2(\count[0] [8]), 
            .I3(\count[0] [7]), .O(n19));
    defparam i7_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut (.I0(\count[0] [3]), .I1(n19), .I2(n20_adj_3523), 
            .I3(GND_net), .O(n6_adj_3524));
    defparam i1_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4_4_lut (.I0(\count[0] [2]), .I1(\count[0] [5]), .I2(\count[0] [1]), 
            .I3(n6_adj_3524), .O(n925));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_548));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26809_2_lut (.I0(n8), .I1(n9), .I2(GND_net), .I3(GND_net), 
            .O(n32443));
    defparam i26809_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26877_4_lut (.I0(n2), .I1(n5), .I2(n4), .I3(n7), .O(n32513));
    defparam i26877_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_845 (.I0(\count[0] [10]), .I1(n32513), .I2(n32443), 
            .I3(n6), .O(n22));
    defparam i10_4_lut_adj_845.LUT_INIT = 16'h0002;
    SB_LUT4 i9_4_lut (.I0(n10), .I1(n3), .I2(n1), .I3(pwm_out_0__N_522), 
            .O(n21));
    defparam i9_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut (.I0(n21), .I1(pause_counter_0), .I2(pwm_out_0__N_518), 
            .I3(n22), .O(n16531));
    defparam i1_4_lut.LUT_INIT = 16'h2303;
    SB_LUT4 i3_4_lut (.I0(\half_duty[0][6] ), .I1(\half_duty[0][5] ), .I2(\count[0] [6]), 
            .I3(\count[0] [5]), .O(n14));   // vhdl/pwm.vhd(80[8:31])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_846 (.I0(\half_duty[0][7] ), .I1(\half_duty[0][3] ), 
            .I2(\count[0] [7]), .I3(\count[0] [3]), .O(n12));   // vhdl/pwm.vhd(80[8:31])
    defparam i1_4_lut_adj_846.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut (.I0(\half_duty[0][2] ), .I1(\half_duty[0][1] ), .I2(\count[0] [2]), 
            .I3(\count[0] [1]), .O(n13));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i5_3_lut (.I0(\half_duty[0][0] ), .I1(\count[0] [9]), .I2(\count[0] [0]), 
            .I3(GND_net), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i31217_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_518), .I2(GND_net), 
            .I3(GND_net), .O(n30927));
    defparam i31217_2_lut.LUT_INIT = 16'h1111;
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n16936));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 count_0__1130_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n25518), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1130_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n25517), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_11 (.CI(n25517), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n25518));
    SB_LUT4 count_0__1130_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n25516), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_10 (.CI(n25516), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n25517));
    SB_LUT4 count_0__1130_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n25515), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_9 (.CI(n25515), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n25516));
    SB_LUT4 count_0__1130_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n25514), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_8 (.CI(n25514), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n25515));
    SB_LUT4 count_0__1130_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n25513), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_7 (.CI(n25513), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n25514));
    SB_LUT4 count_0__1130_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n25512), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_6 (.CI(n25512), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n25513));
    SB_LUT4 count_0__1130_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n25511), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_5 (.CI(n25511), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n25512));
    SB_LUT4 count_0__1130_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n25510), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_4 (.CI(n25510), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n25511));
    SB_LUT4 count_0__1130_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n25509), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_3 (.CI(n25509), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n25510));
    SB_LUT4 count_0__1130_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1130_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1130_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n25509));
    SB_LUT4 add_2006_24_lut (.I0(GND_net), .I1(n5538[22]), .I2(pwm_setpoint[22]), 
            .I3(n24916), .O(half_duty_new_9__N_600[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2006_23_lut (.I0(GND_net), .I1(n5538[21]), .I2(pwm_setpoint[21]), 
            .I3(n24915), .O(half_duty_new_9__N_600[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_23 (.CI(n24915), .I0(n5538[21]), .I1(pwm_setpoint[21]), 
            .CO(n24916));
    SB_LUT4 add_2006_22_lut (.I0(GND_net), .I1(n5538[20]), .I2(pwm_setpoint[20]), 
            .I3(n24914), .O(half_duty_new_9__N_600[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_22 (.CI(n24914), .I0(n5538[20]), .I1(pwm_setpoint[20]), 
            .CO(n24915));
    SB_LUT4 add_2006_21_lut (.I0(GND_net), .I1(n5538[19]), .I2(pwm_setpoint[19]), 
            .I3(n24913), .O(half_duty_new_9__N_600[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_21 (.CI(n24913), .I0(n5538[19]), .I1(pwm_setpoint[19]), 
            .CO(n24914));
    SB_LUT4 add_2006_20_lut (.I0(GND_net), .I1(n5538[18]), .I2(pwm_setpoint[18]), 
            .I3(n24912), .O(half_duty_new_9__N_600[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_20 (.CI(n24912), .I0(n5538[18]), .I1(pwm_setpoint[18]), 
            .CO(n24913));
    SB_LUT4 add_2006_19_lut (.I0(GND_net), .I1(n5538[17]), .I2(pwm_setpoint[17]), 
            .I3(n24911), .O(half_duty_new_9__N_600[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_19 (.CI(n24911), .I0(n5538[17]), .I1(pwm_setpoint[17]), 
            .CO(n24912));
    SB_LUT4 add_2006_18_lut (.I0(GND_net), .I1(n5538[16]), .I2(pwm_setpoint[16]), 
            .I3(n24910), .O(half_duty_new_9__N_600[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_18 (.CI(n24910), .I0(n5538[16]), .I1(pwm_setpoint[16]), 
            .CO(n24911));
    SB_LUT4 add_2006_17_lut (.I0(GND_net), .I1(n5538[15]), .I2(pwm_setpoint[15]), 
            .I3(n24909), .O(half_duty_new_9__N_600[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2006_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2006_17 (.CI(n24909), .I0(n5538[15]), .I1(pwm_setpoint[15]), 
            .CO(n24910));
    SB_CARRY add_2006_16 (.CI(n24908), .I0(n5538[14]), .I1(pwm_setpoint[14]), 
            .CO(n24909));
    SB_CARRY add_2006_15 (.CI(n24907), .I0(n5538[13]), .I1(pwm_setpoint[13]), 
            .CO(n24908));
    SB_CARRY add_2006_14 (.CI(n24906), .I0(n5538[12]), .I1(pwm_setpoint[12]), 
            .CO(n24907));
    SB_CARRY add_2006_13 (.CI(n24905), .I0(n5538[11]), .I1(pwm_setpoint[11]), 
            .CO(n24906));
    SB_CARRY add_2006_12 (.CI(n24904), .I0(n5538[10]), .I1(pwm_setpoint[10]), 
            .CO(n24905));
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_523[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut_adj_847 (.I0(\count[0] [8]), .I1(n13), .I2(n12), 
            .I3(n14), .O(n20));   // vhdl/pwm.vhd(80[8:31])
    defparam i9_4_lut_adj_847.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[1] , GND_net, \Kp[0] , \Kp[2] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , PWMLimit, setpoint, 
            duty, clk32MHz, motor_state, VCC_net, n36858) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input \Kp[1] ;
    input GND_net;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input [23:0]PWMLimit;
    input [23:0]setpoint;
    output [23:0]duty;
    input clk32MHz;
    input [23:0]motor_state;
    input VCC_net;
    output n36858;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n107, n38, n180, n253, n326, n399, n472, n545, n110, 
        n41, n183, n256, n329;
    wire [23:0]n1;
    
    wire n402, n475, n548, n113, n44, n186, n259, n332, n405, 
        n478, n551, n116, n47, n189, n262, n335, n408, n481, 
        n554, n119, n50;
    wire [23:0]n1_adj_3521;
    
    wire n192, n265, n338, n411, n484, n557, n122, n53, n195, 
        n268, n341, n414, n487, n560, n125, n41_adj_3422, n56, 
        n39, n45, n37, n29, n31, n43, n23_adj_3423, n25_adj_3424, 
        n35, n33, n11, n13, n15, n27, n9_adj_3425, n17, n19, 
        n21, n34879, n34873, n12, n30, n34391, n34888, n35411;
    wire [23:0]duty_23__N_3291;
    
    wire n35978, n198, n35610, n36047;
    wire [23:0]\PID_CONTROLLER.err_23__N_3315 ;
    
    wire n271, n6_adj_3426, n35644, n35645, n16, n24_adj_3427, n34858, 
        n8_adj_3428, n34855, n35688, n35242, n4_adj_3429, n35640, 
        n35641, n344, n417, n34869, n6_adj_3430;
    wire [3:0]n8576;
    wire [4:0]n8569;
    
    wire n204, n10, n34867, n36008, n35244, n36124;
    wire [1:0]n8587;
    
    wire n36125, n131, n62, n36086, n34860, n35919, n35250, n36030, 
        duty_23__N_3363;
    wire [23:0]n103;
    
    wire n39_adj_3431, n4_adj_3432;
    wire [2:0]n8582;
    
    wire n490, n12_adj_3433, n8_adj_3434, n41_adj_3436, n11_adj_3437, 
        n45_adj_3438, n6_adj_3439, n43_adj_3440, n24565, n37_adj_3441, 
        n18, n29_adj_3443, n31_adj_3444, n23_adj_3446, n25_adj_3447, 
        n35_adj_3449, n13_adj_3450, n11_adj_3452, n13_adj_3453, n27_adj_3454, 
        n4_adj_3455, n31625, n15_adj_3456, n33_adj_3457, n9_adj_3458, 
        n17_adj_3460, n19_adj_3461, n21_adj_3462, n34813, n34806, 
        n12_adj_3464, n10_adj_3465, n30_adj_3466, n34839, n35383, 
        n35379, n35972, n35594, n36045, n16_adj_3468, n6_adj_3469, 
        n35634, n35635, n8_adj_3470, n24_adj_3471, n34792, n34790, 
        n35690, n35252, n4_adj_3472, n35632, n35633, n34802, n34800, 
        n36010, n35254, n36126, n36127, n36082, n34794, n35921, 
        n35260, n36032, n102;
    wire [23:0]duty_23__N_3339;
    
    wire n24795, n24794, n24793, n24792, n24791, n24790, n24789, 
        n24788, n24787, n24786, n24785, n24784, n24783, n24782, 
        n24781, n24780, n24779, n24778, n24777, n24776;
    wire [5:0]n8561;
    
    wire n25888, n25887, n25886, n25885, n25884;
    wire [6:0]n8552;
    
    wire n25883, n25882, n25881, n25880, n25879, n25878;
    wire [7:0]n8542;
    
    wire n25877, n25876, n25875, n24775, n24774, n24773, n25874, 
        n25873, n25872, n25871, n24772;
    wire [8:0]n8531;
    
    wire n25870, n25869, n25868, n25867, n25866, n25865, n25864, 
        n24771, n24770, n24769, n24768, n25863;
    wire [9:0]n8519;
    
    wire n25862, n25861, n25860, n25859, n25858, n25857, n25856, 
        n25855, n25854;
    wire [10:0]n8506;
    
    wire n25853, n25852, n24767, n25851, n25850, n25849, n25848, 
        n24766, n25847, n24765, n25846, n25845, n25844;
    wire [11:0]n8492;
    
    wire n25843, n25842, n25841, n25840, n25839, n25838, n25837, 
        n25836, n25835, n25834, n25833;
    wire [12:0]n8477;
    
    wire n25832, n25831, n25830, n25829, n25828, n25827, n542, 
        n25826, n469, n25825, n396, n25824, n24764, n323, n25823, 
        n250, n25822, n177, n25821, n35_adj_3490, n104_adj_3491;
    wire [13:0]n8461;
    
    wire n25820, n25819, n24763, n25818, n25817, n25816, n25815, 
        n25814, n539, n25813, n466, n25812, n24762, n393, n25811, 
        n24761, n320, n25810, n24760, n24759, n24758, n24757, 
        n247, n25809, n24756, n24755, n24754, n24753, n24752, 
        n24751, n174, n25808, n32, n101;
    wire [14:0]n8444;
    
    wire n25807, n25806, n25805, n25804, n25803, n25802, n25801, 
        n25800, n536, n25799, n463, n25798, n390, n25797, n317, 
        n25796, n244, n25795, n171, n25794, n29_adj_3506, n98;
    wire [15:0]n8426;
    
    wire n25793, n25792, n25791, n25790, n25789, n25788, n25787, 
        n25786, n25785, n533, n25784, n460, n25783, n387, n25782, 
        n314, n25781, n241, n25780, n168, n25779, n26, n95;
    wire [16:0]n8407;
    
    wire n25778, n25777, n25776, n25775, n25774, n25773, n25772, 
        n25771, n25770, n25769, n530, n25768, n457, n25767, n384, 
        n25766, n311, n25765, n238, n25764, n165, n25763, n23_adj_3507, 
        n92;
    wire [17:0]n8387;
    
    wire n25762, n25761, n25760, n25759, n25758, n25757, n25756, 
        n25755, n25754, n25753, n25752, n527, n25751, n454, n25750, 
        n381, n25749, n308, n25748, n235, n25747, n162, n25746, 
        n20_adj_3508, n89;
    wire [18:0]n8366;
    
    wire n25745, n25744, n25743, n25742, n25741, n25740, n25739, 
        n25738, n25737, n25736, n25735, n25734, n524, n25733, 
        n451, n25732, n378, n25731, n305, n25730, n232, n25729, 
        n159, n25728, n17_adj_3509, n86, n4_adj_3510;
    wire [19:0]n8344;
    
    wire n25727, n25726, n25725, n25724, n25723, n25722, n25721, 
        n25720, n25719, n25718, n25717, n25716, n25715, n521, 
        n25714, n448, n25713, n375, n25712, n302, n25711, n229, 
        n25710, n156, n25709, n14_adj_3511, n83;
    wire [20:0]n8321;
    
    wire n25708, n25707, n25706, n25705, n25704, n25703, n25702, 
        n25701, n25700, n25699, n25698, n25697, n25696, n25695, 
        n518, n25694, n445, n25693, n24463, n372, n25692, n299, 
        n25691, n226, n25690, n153, n25689, n11_adj_3512, n80, 
        n34262;
    wire [21:0]n8297;
    
    wire n25688;
    wire [47:0]n28;
    
    wire n25687, n25686, n25685, n25684, n25683, n25682, n25681, 
        n25680, n25679, n25678, n25677, n25676, n24750, n25675, 
        n25674, n25673, n512, n25672, n439, n25671, n366, n25670, 
        n293, n25669, n220, n25668, n147, n25667, n5_adj_3517, 
        n74_adj_3518, n25666, n25665, n25664, n25663, n25662, n25661, 
        n25660, n25659, n25658, n25657, n25656, n25655, n25654, 
        n25653, n25652, n515, n25651, n442, n25650, n369, n25649, 
        n296, n25648, n223, n25647, n150, n25646, n8_adj_3519, 
        n77, n24540;
    
    SB_LUT4 mult_4_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[0]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[1]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[2]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[3]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3422));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_4_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3423));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3424));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3425));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29241_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9_adj_3425), 
            .O(n34879));
    defparam i29241_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29235_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n34873));
    defparam i29235_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(duty[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29250_4_lut (.I0(n13), .I1(n11), .I2(n9_adj_3425), .I3(n34391), 
            .O(n34888));
    defparam i29250_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29773_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n34888), 
            .O(n35411));
    defparam i29773_4_lut.LUT_INIT = 16'heeef;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3291[0]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 i30339_4_lut (.I0(n25_adj_3424), .I1(n23_adj_3423), .I2(n21), 
            .I3(n35411), .O(n35978));
    defparam i30339_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_4_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29971_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n35978), 
            .O(n35610));
    defparam i29971_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30408_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n35610), 
            .O(n36047));
    defparam i30408_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [0]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 mult_4_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30005_3_lut (.I0(n6_adj_3426), .I1(duty[10]), .I2(n21), .I3(GND_net), 
            .O(n35644));   // verilog/motorControl.v(43[10:25])
    defparam i30005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30006_3_lut (.I0(n35644), .I1(duty[11]), .I2(n23_adj_3423), 
            .I3(GND_net), .O(n35645));   // verilog/motorControl.v(43[10:25])
    defparam i30006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(duty[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_3427));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29220_4_lut (.I0(n43), .I1(n25_adj_3424), .I2(n23_adj_3423), 
            .I3(n34879), .O(n34858));
    defparam i29220_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30049_4_lut (.I0(n24_adj_3427), .I1(n8_adj_3428), .I2(n45), 
            .I3(n34855), .O(n35688));   // verilog/motorControl.v(43[10:25])
    defparam i30049_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29604_3_lut (.I0(n35645), .I1(duty[12]), .I2(n25_adj_3424), 
            .I3(GND_net), .O(n35242));   // verilog/motorControl.v(43[10:25])
    defparam i29604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(PWMLimit[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(duty[0]), .O(n4_adj_3429));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30001_3_lut (.I0(n4_adj_3429), .I1(duty[13]), .I2(n27), .I3(GND_net), 
            .O(n35640));   // verilog/motorControl.v(43[10:25])
    defparam i30001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30002_3_lut (.I0(n35640), .I1(duty[14]), .I2(n29), .I3(GND_net), 
            .O(n35641));   // verilog/motorControl.v(43[10:25])
    defparam i30002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29231_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n34873), 
            .O(n34869));
    defparam i29231_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i2_4_lut (.I0(n6_adj_3430), .I1(\Kp[4] ), .I2(n8576[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8569[3]));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_4_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30369_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n34867), 
            .O(n36008));   // verilog/motorControl.v(43[10:25])
    defparam i30369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29606_3_lut (.I0(n35641), .I1(duty[15]), .I2(n31), .I3(GND_net), 
            .O(n35244));   // verilog/motorControl.v(43[10:25])
    defparam i29606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30485_4_lut (.I0(n35244), .I1(n36008), .I2(n35), .I3(n34869), 
            .O(n36124));   // verilog/motorControl.v(43[10:25])
    defparam i30485_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i20234_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8587[0]));   // verilog/motorControl.v(41[17:23])
    defparam i20234_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i30486_3_lut (.I0(n36124), .I1(duty[18]), .I2(n37), .I3(GND_net), 
            .O(n36125));   // verilog/motorControl.v(43[10:25])
    defparam i30486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30447_3_lut (.I0(n36125), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n36086));   // verilog/motorControl.v(43[10:25])
    defparam i30447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29222_4_lut (.I0(n43), .I1(n41_adj_3422), .I2(n39), .I3(n36047), 
            .O(n34860));
    defparam i29222_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30280_4_lut (.I0(n35242), .I1(n35688), .I2(n45), .I3(n34858), 
            .O(n35919));   // verilog/motorControl.v(43[10:25])
    defparam i30280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29612_3_lut (.I0(n36086), .I1(duty[20]), .I2(n41_adj_3422), 
            .I3(GND_net), .O(n35250));   // verilog/motorControl.v(43[10:25])
    defparam i29612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30391_4_lut (.I0(n35250), .I1(n35919), .I2(n45), .I3(n34860), 
            .O(n36030));   // verilog/motorControl.v(43[10:25])
    defparam i30391_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30392_3_lut (.I0(n36030), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3363));   // verilog/motorControl.v(43[10:25])
    defparam i30392_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_7_i39_2_lut (.I0(duty[19]), .I1(n103[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3431));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_840 (.I0(n4_adj_3432), .I1(\Kp[3] ), .I2(n8582[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8576[2]));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut_adj_840.LUT_INIT = 16'h965a;
    SB_LUT4 mult_4_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_841 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_3433));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut_adj_841.LUT_INIT = 16'h9c50;
    SB_LUT4 i20170_4_lut (.I0(n8576[2]), .I1(\Kp[4] ), .I2(n6_adj_3430), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_3434));   // verilog/motorControl.v(41[17:23])
    defparam i20170_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 LessThan_7_i41_2_lut (.I0(duty[20]), .I1(n103[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3436));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_3437));   // verilog/motorControl.v(41[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_7_i45_2_lut (.I0(duty[22]), .I1(n103[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3438));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i20201_4_lut (.I0(n8582[1]), .I1(\Kp[3] ), .I2(n4_adj_3432), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_3439));   // verilog/motorControl.v(41[17:23])
    defparam i20201_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 LessThan_7_i43_2_lut (.I0(duty[21]), .I1(n103[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3440));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i20236_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n24565));   // verilog/motorControl.v(41[17:23])
    defparam i20236_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_7_i37_2_lut (.I0(duty[18]), .I1(n103[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3441));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3439), .I1(n11_adj_3437), .I2(n8_adj_3434), 
            .I3(n12_adj_3433), .O(n18));   // verilog/motorControl.v(41[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_7_i29_2_lut (.I0(duty[14]), .I1(n103[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3443));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i31_2_lut (.I0(duty[15]), .I1(n103[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3444));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i23_2_lut (.I0(duty[11]), .I1(n103[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3446));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i25_2_lut (.I0(duty[12]), .I1(n103[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3447));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i35_2_lut (.I0(duty[17]), .I1(n103[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3449));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_3450));   // verilog/motorControl.v(41[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_7_i11_2_lut (.I0(duty[5]), .I1(n103[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3452));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i13_2_lut (.I0(duty[6]), .I1(n103[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3453));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i27_2_lut (.I0(duty[13]), .I1(n103[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3454));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(n13_adj_3450), .I1(n18), .I2(n24565), .I3(n4_adj_3455), 
            .O(n31625));   // verilog/motorControl.v(41[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_7_i15_2_lut (.I0(duty[7]), .I1(n103[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3456));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i33_2_lut (.I0(duty[16]), .I1(n103[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3457));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i9_2_lut (.I0(duty[4]), .I1(n103[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3458));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i17_2_lut (.I0(duty[8]), .I1(n103[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3460));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i19_2_lut (.I0(duty[9]), .I1(n103[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3461));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i21_2_lut (.I0(duty[10]), .I1(n103[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3462));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[4]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29176_4_lut (.I0(n21_adj_3462), .I1(n19_adj_3461), .I2(n17_adj_3460), 
            .I3(n9_adj_3458), .O(n34813));
    defparam i29176_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29169_4_lut (.I0(n27_adj_3454), .I1(n15_adj_3456), .I2(n13_adj_3453), 
            .I3(n11_adj_3452), .O(n34806));
    defparam i29169_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_7_i12_3_lut (.I0(n103[7]), .I1(n103[16]), .I2(n33_adj_3457), 
            .I3(GND_net), .O(n12_adj_3464));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i10_3_lut (.I0(n103[5]), .I1(n103[6]), .I2(n13_adj_3453), 
            .I3(GND_net), .O(n10_adj_3465));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[5]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_7_i30_3_lut (.I0(n12_adj_3464), .I1(n103[17]), .I2(n35_adj_3449), 
            .I3(GND_net), .O(n30_adj_3466));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29745_4_lut (.I0(n13_adj_3453), .I1(n11_adj_3452), .I2(n9_adj_3458), 
            .I3(n34839), .O(n35383));
    defparam i29745_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[6]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29741_4_lut (.I0(n19_adj_3461), .I1(n17_adj_3460), .I2(n15_adj_3456), 
            .I3(n35383), .O(n35379));
    defparam i29741_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30333_4_lut (.I0(n25_adj_3447), .I1(n23_adj_3446), .I2(n21_adj_3462), 
            .I3(n35379), .O(n35972));
    defparam i30333_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29955_4_lut (.I0(n31_adj_3444), .I1(n29_adj_3443), .I2(n27_adj_3454), 
            .I3(n35972), .O(n35594));
    defparam i29955_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30406_4_lut (.I0(n37_adj_3441), .I1(n35_adj_3449), .I2(n33_adj_3457), 
            .I3(n35594), .O(n36045));
    defparam i30406_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_7_i16_3_lut (.I0(n103[9]), .I1(n103[21]), .I2(n43_adj_3440), 
            .I3(GND_net), .O(n16_adj_3468));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29995_3_lut (.I0(n6_adj_3469), .I1(n103[10]), .I2(n21_adj_3462), 
            .I3(GND_net), .O(n35634));   // verilog/motorControl.v(45[19:35])
    defparam i29995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29996_3_lut (.I0(n35634), .I1(n103[11]), .I2(n23_adj_3446), 
            .I3(GND_net), .O(n35635));   // verilog/motorControl.v(45[19:35])
    defparam i29996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i8_3_lut (.I0(n103[4]), .I1(n103[8]), .I2(n17_adj_3460), 
            .I3(GND_net), .O(n8_adj_3470));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i24_3_lut (.I0(n16_adj_3468), .I1(n103[22]), .I2(n45_adj_3438), 
            .I3(GND_net), .O(n24_adj_3471));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29155_4_lut (.I0(n43_adj_3440), .I1(n25_adj_3447), .I2(n23_adj_3446), 
            .I3(n34813), .O(n34792));
    defparam i29155_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30051_4_lut (.I0(n24_adj_3471), .I1(n8_adj_3470), .I2(n45_adj_3438), 
            .I3(n34790), .O(n35690));   // verilog/motorControl.v(45[19:35])
    defparam i30051_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29614_3_lut (.I0(n35635), .I1(n103[12]), .I2(n25_adj_3447), 
            .I3(GND_net), .O(n35252));   // verilog/motorControl.v(45[19:35])
    defparam i29614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i4_4_lut (.I0(n103[0]), .I1(n103[1]), .I2(duty[1]), 
            .I3(duty[0]), .O(n4_adj_3472));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i29993_3_lut (.I0(n4_adj_3472), .I1(n103[13]), .I2(n27_adj_3454), 
            .I3(GND_net), .O(n35632));   // verilog/motorControl.v(45[19:35])
    defparam i29993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29994_3_lut (.I0(n35632), .I1(n103[14]), .I2(n29_adj_3443), 
            .I3(GND_net), .O(n35633));   // verilog/motorControl.v(45[19:35])
    defparam i29994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[7]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29165_4_lut (.I0(n33_adj_3457), .I1(n31_adj_3444), .I2(n29_adj_3443), 
            .I3(n34806), .O(n34802));
    defparam i29165_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30371_4_lut (.I0(n30_adj_3466), .I1(n10_adj_3465), .I2(n35_adj_3449), 
            .I3(n34800), .O(n36010));   // verilog/motorControl.v(45[19:35])
    defparam i30371_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29616_3_lut (.I0(n35633), .I1(n103[15]), .I2(n31_adj_3444), 
            .I3(GND_net), .O(n35254));   // verilog/motorControl.v(45[19:35])
    defparam i29616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30487_4_lut (.I0(n35254), .I1(n36010), .I2(n35_adj_3449), 
            .I3(n34802), .O(n36126));   // verilog/motorControl.v(45[19:35])
    defparam i30487_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30488_3_lut (.I0(n36126), .I1(n103[18]), .I2(n37_adj_3441), 
            .I3(GND_net), .O(n36127));   // verilog/motorControl.v(45[19:35])
    defparam i30488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30443_3_lut (.I0(n36127), .I1(n103[19]), .I2(n39_adj_3431), 
            .I3(GND_net), .O(n36082));   // verilog/motorControl.v(45[19:35])
    defparam i30443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[8]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29157_4_lut (.I0(n43_adj_3440), .I1(n41_adj_3436), .I2(n39_adj_3431), 
            .I3(n36045), .O(n34794));
    defparam i29157_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30282_4_lut (.I0(n35252), .I1(n35690), .I2(n45_adj_3438), 
            .I3(n34792), .O(n35921));   // verilog/motorControl.v(45[19:35])
    defparam i30282_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[9]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29622_3_lut (.I0(n36082), .I1(n103[20]), .I2(n41_adj_3436), 
            .I3(GND_net), .O(n35260));   // verilog/motorControl.v(45[19:35])
    defparam i29622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30393_4_lut (.I0(n35260), .I1(n35921), .I2(n45_adj_3438), 
            .I3(n34794), .O(n36032));   // verilog/motorControl.v(45[19:35])
    defparam i30393_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[10]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30394_3_lut (.I0(n36032), .I1(duty[23]), .I2(n103[23]), .I3(GND_net), 
            .O(n102));   // verilog/motorControl.v(45[19:35])
    defparam i30394_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_9_i1_4_lut (.I0(\PID_CONTROLLER.err [0]), .I1(n103[0]), 
            .I2(n102), .I3(\Kp[0] ), .O(duty_23__N_3339[0]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i1_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 duty_23__I_0_18_i1_3_lut (.I0(duty_23__N_3339[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[0]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[11]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_3521[23]), .I3(n24795), .O(\PID_CONTROLLER.err_23__N_3315 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[12]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_3521[22]), .I3(n24794), .O(\PID_CONTROLLER.err_23__N_3315 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n24794), .I0(motor_state[22]), 
            .I1(n1_adj_3521[22]), .CO(n24795));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_3521[21]), .I3(n24793), .O(\PID_CONTROLLER.err_23__N_3315 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n24793), .I0(motor_state[21]), 
            .I1(n1_adj_3521[21]), .CO(n24794));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_3521[20]), .I3(n24792), .O(\PID_CONTROLLER.err_23__N_3315 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[13]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n24792), .I0(motor_state[20]), 
            .I1(n1_adj_3521[20]), .CO(n24793));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_3521[19]), .I3(n24791), .O(\PID_CONTROLLER.err_23__N_3315 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n24791), .I0(motor_state[19]), 
            .I1(n1_adj_3521[19]), .CO(n24792));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_3521[18]), .I3(n24790), .O(\PID_CONTROLLER.err_23__N_3315 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n24790), .I0(motor_state[18]), 
            .I1(n1_adj_3521[18]), .CO(n24791));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_3521[17]), .I3(n24789), .O(\PID_CONTROLLER.err_23__N_3315 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n24789), .I0(motor_state[17]), 
            .I1(n1_adj_3521[17]), .CO(n24790));
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[14]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[15]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[16]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_3521[16]), .I3(n24788), .O(\PID_CONTROLLER.err_23__N_3315 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[17]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[18]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[19]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n24788), .I0(motor_state[16]), 
            .I1(n1_adj_3521[16]), .CO(n24789));
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_3521[15]), .I3(n24787), .O(\PID_CONTROLLER.err_23__N_3315 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[20]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[21]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n24787), .I0(motor_state[15]), 
            .I1(n1_adj_3521[15]), .CO(n24788));
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[22]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_3521[14]), .I3(n24786), .O(\PID_CONTROLLER.err_23__N_3315 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3521[23]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n24786), .I0(motor_state[14]), 
            .I1(n1_adj_3521[14]), .CO(n24787));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_3521[13]), .I3(n24785), .O(\PID_CONTROLLER.err_23__N_3315 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n24785), .I0(motor_state[13]), 
            .I1(n1_adj_3521[13]), .CO(n24786));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_3521[12]), .I3(n24784), .O(\PID_CONTROLLER.err_23__N_3315 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n24784), .I0(motor_state[12]), 
            .I1(n1_adj_3521[12]), .CO(n24785));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_3521[11]), .I3(n24783), .O(\PID_CONTROLLER.err_23__N_3315 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n24783), .I0(motor_state[11]), 
            .I1(n1_adj_3521[11]), .CO(n24784));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_3521[10]), .I3(n24782), .O(\PID_CONTROLLER.err_23__N_3315 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n24782), .I0(motor_state[10]), 
            .I1(n1_adj_3521[10]), .CO(n24783));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_3521[9]), .I3(n24781), .O(\PID_CONTROLLER.err_23__N_3315 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n24781), .I0(motor_state[9]), .I1(n1_adj_3521[9]), 
            .CO(n24782));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_3521[8]), .I3(n24780), .O(\PID_CONTROLLER.err_23__N_3315 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n24780), .I0(motor_state[8]), .I1(n1_adj_3521[8]), 
            .CO(n24781));
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_3521[7]), .I3(n24779), .O(\PID_CONTROLLER.err_23__N_3315 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n24779), .I0(motor_state[7]), .I1(n1_adj_3521[7]), 
            .CO(n24780));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_3521[6]), .I3(n24778), .O(\PID_CONTROLLER.err_23__N_3315 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n24778), .I0(motor_state[6]), .I1(n1_adj_3521[6]), 
            .CO(n24779));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_3521[5]), .I3(n24777), .O(\PID_CONTROLLER.err_23__N_3315 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n24777), .I0(motor_state[5]), .I1(n1_adj_3521[5]), 
            .CO(n24778));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_3521[4]), .I3(n24776), .O(\PID_CONTROLLER.err_23__N_3315 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_7_lut (.I0(GND_net), .I1(n31625), .I2(n490), .I3(n25888), 
            .O(n8561[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_6_lut (.I0(GND_net), .I1(n8569[3]), .I2(n417), .I3(n25887), 
            .O(n8561[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_6 (.CI(n25887), .I0(n8569[3]), .I1(n417), .CO(n25888));
    SB_LUT4 add_4444_5_lut (.I0(GND_net), .I1(n8569[2]), .I2(n344), .I3(n25886), 
            .O(n8561[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_5 (.CI(n25886), .I0(n8569[2]), .I1(n344), .CO(n25887));
    SB_LUT4 add_4444_4_lut (.I0(GND_net), .I1(n8569[1]), .I2(n271), .I3(n25885), 
            .O(n8561[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_4 (.CI(n25885), .I0(n8569[1]), .I1(n271), .CO(n25886));
    SB_LUT4 add_4444_3_lut (.I0(GND_net), .I1(n8569[0]), .I2(n198), .I3(n25884), 
            .O(n8561[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_3 (.CI(n25884), .I0(n8569[0]), .I1(n198), .CO(n25885));
    SB_LUT4 add_4444_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n8561[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n25884));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n24776), .I0(motor_state[4]), .I1(n1_adj_3521[4]), 
            .CO(n24777));
    SB_LUT4 add_4443_8_lut (.I0(GND_net), .I1(n8561[5]), .I2(n560), .I3(n25883), 
            .O(n8552[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4443_7_lut (.I0(GND_net), .I1(n8561[4]), .I2(n487), .I3(n25882), 
            .O(n8552[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_7 (.CI(n25882), .I0(n8561[4]), .I1(n487), .CO(n25883));
    SB_LUT4 add_4443_6_lut (.I0(GND_net), .I1(n8561[3]), .I2(n414), .I3(n25881), 
            .O(n8552[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_6 (.CI(n25881), .I0(n8561[3]), .I1(n414), .CO(n25882));
    SB_LUT4 add_4443_5_lut (.I0(GND_net), .I1(n8561[2]), .I2(n341), .I3(n25880), 
            .O(n8552[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_5 (.CI(n25880), .I0(n8561[2]), .I1(n341), .CO(n25881));
    SB_LUT4 add_4443_4_lut (.I0(GND_net), .I1(n8561[1]), .I2(n268), .I3(n25879), 
            .O(n8552[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_4 (.CI(n25879), .I0(n8561[1]), .I1(n268), .CO(n25880));
    SB_LUT4 add_4443_3_lut (.I0(GND_net), .I1(n8561[0]), .I2(n195), .I3(n25878), 
            .O(n8552[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_3 (.CI(n25878), .I0(n8561[0]), .I1(n195), .CO(n25879));
    SB_LUT4 add_4443_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n8552[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n25878));
    SB_LUT4 add_4442_9_lut (.I0(GND_net), .I1(n8552[6]), .I2(GND_net), 
            .I3(n25877), .O(n8542[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_8_lut (.I0(GND_net), .I1(n8552[5]), .I2(n557), .I3(n25876), 
            .O(n8542[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_8 (.CI(n25876), .I0(n8552[5]), .I1(n557), .CO(n25877));
    SB_LUT4 add_4442_7_lut (.I0(GND_net), .I1(n8552[4]), .I2(n484), .I3(n25875), 
            .O(n8542[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_7 (.CI(n25875), .I0(n8552[4]), .I1(n484), .CO(n25876));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_3521[3]), .I3(n24775), .O(\PID_CONTROLLER.err_23__N_3315 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n24775), .I0(motor_state[3]), .I1(n1_adj_3521[3]), 
            .CO(n24776));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_3521[2]), .I3(n24774), .O(\PID_CONTROLLER.err_23__N_3315 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n24774), .I0(motor_state[2]), .I1(n1_adj_3521[2]), 
            .CO(n24775));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_3521[1]), .I3(n24773), .O(\PID_CONTROLLER.err_23__N_3315 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_6_lut (.I0(GND_net), .I1(n8552[3]), .I2(n411), .I3(n25874), 
            .O(n8542[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_6 (.CI(n25874), .I0(n8552[3]), .I1(n411), .CO(n25875));
    SB_LUT4 add_4442_5_lut (.I0(GND_net), .I1(n8552[2]), .I2(n338), .I3(n25873), 
            .O(n8542[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_5 (.CI(n25873), .I0(n8552[2]), .I1(n338), .CO(n25874));
    SB_LUT4 add_4442_4_lut (.I0(GND_net), .I1(n8552[1]), .I2(n265), .I3(n25872), 
            .O(n8542[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_4 (.CI(n25872), .I0(n8552[1]), .I1(n265), .CO(n25873));
    SB_LUT4 add_4442_3_lut (.I0(GND_net), .I1(n8552[0]), .I2(n192), .I3(n25871), 
            .O(n8542[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n24773), .I0(motor_state[1]), .I1(n1_adj_3521[1]), 
            .CO(n24774));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_3521[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3315 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_3 (.CI(n25871), .I0(n8552[0]), .I1(n192), .CO(n25872));
    SB_LUT4 add_4442_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n8542[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n25871));
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_3521[0]), 
            .CO(n24773));
    SB_LUT4 unary_minus_8_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n24772), .O(n103[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_10_lut (.I0(GND_net), .I1(n8542[7]), .I2(GND_net), 
            .I3(n25870), .O(n8531[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_9_lut (.I0(GND_net), .I1(n8542[6]), .I2(GND_net), 
            .I3(n25869), .O(n8531[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_9 (.CI(n25869), .I0(n8542[6]), .I1(GND_net), .CO(n25870));
    SB_LUT4 add_4441_8_lut (.I0(GND_net), .I1(n8542[5]), .I2(n554), .I3(n25868), 
            .O(n8531[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_8 (.CI(n25868), .I0(n8542[5]), .I1(n554), .CO(n25869));
    SB_LUT4 add_4441_7_lut (.I0(GND_net), .I1(n8542[4]), .I2(n481), .I3(n25867), 
            .O(n8531[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_7 (.CI(n25867), .I0(n8542[4]), .I1(n481), .CO(n25868));
    SB_LUT4 add_4441_6_lut (.I0(GND_net), .I1(n8542[3]), .I2(n408), .I3(n25866), 
            .O(n8531[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_6 (.CI(n25866), .I0(n8542[3]), .I1(n408), .CO(n25867));
    SB_LUT4 add_4441_5_lut (.I0(GND_net), .I1(n8542[2]), .I2(n335), .I3(n25865), 
            .O(n8531[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_5 (.CI(n25865), .I0(n8542[2]), .I1(n335), .CO(n25866));
    SB_LUT4 add_4441_4_lut (.I0(GND_net), .I1(n8542[1]), .I2(n262), .I3(n25864), 
            .O(n8531[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n24771), .O(n103[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_24 (.CI(n24771), .I0(GND_net), .I1(n1[22]), 
            .CO(n24772));
    SB_LUT4 unary_minus_8_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n24770), .O(n103[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_23 (.CI(n24770), .I0(GND_net), .I1(n1[21]), 
            .CO(n24771));
    SB_LUT4 unary_minus_8_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n24769), .O(n103[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_22 (.CI(n24769), .I0(GND_net), .I1(n1[20]), 
            .CO(n24770));
    SB_LUT4 unary_minus_8_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n24768), .O(n103[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_21 (.CI(n24768), .I0(GND_net), .I1(n1[19]), 
            .CO(n24769));
    SB_CARRY add_4441_4 (.CI(n25864), .I0(n8542[1]), .I1(n262), .CO(n25865));
    SB_LUT4 add_4441_3_lut (.I0(GND_net), .I1(n8542[0]), .I2(n189), .I3(n25863), 
            .O(n8531[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_3 (.CI(n25863), .I0(n8542[0]), .I1(n189), .CO(n25864));
    SB_LUT4 add_4441_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n8531[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n25863));
    SB_LUT4 add_4440_11_lut (.I0(GND_net), .I1(n8531[8]), .I2(GND_net), 
            .I3(n25862), .O(n8519[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4440_10_lut (.I0(GND_net), .I1(n8531[7]), .I2(GND_net), 
            .I3(n25861), .O(n8519[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_10 (.CI(n25861), .I0(n8531[7]), .I1(GND_net), .CO(n25862));
    SB_LUT4 add_4440_9_lut (.I0(GND_net), .I1(n8531[6]), .I2(GND_net), 
            .I3(n25860), .O(n8519[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_9 (.CI(n25860), .I0(n8531[6]), .I1(GND_net), .CO(n25861));
    SB_LUT4 add_4440_8_lut (.I0(GND_net), .I1(n8531[5]), .I2(n551), .I3(n25859), 
            .O(n8519[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_8 (.CI(n25859), .I0(n8531[5]), .I1(n551), .CO(n25860));
    SB_LUT4 add_4440_7_lut (.I0(GND_net), .I1(n8531[4]), .I2(n478), .I3(n25858), 
            .O(n8519[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_7 (.CI(n25858), .I0(n8531[4]), .I1(n478), .CO(n25859));
    SB_LUT4 add_4440_6_lut (.I0(GND_net), .I1(n8531[3]), .I2(n405), .I3(n25857), 
            .O(n8519[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_6 (.CI(n25857), .I0(n8531[3]), .I1(n405), .CO(n25858));
    SB_LUT4 add_4440_5_lut (.I0(GND_net), .I1(n8531[2]), .I2(n332), .I3(n25856), 
            .O(n8519[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_5 (.CI(n25856), .I0(n8531[2]), .I1(n332), .CO(n25857));
    SB_LUT4 add_4440_4_lut (.I0(GND_net), .I1(n8531[1]), .I2(n259), .I3(n25855), 
            .O(n8519[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_4 (.CI(n25855), .I0(n8531[1]), .I1(n259), .CO(n25856));
    SB_LUT4 add_4440_3_lut (.I0(GND_net), .I1(n8531[0]), .I2(n186), .I3(n25854), 
            .O(n8519[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_3 (.CI(n25854), .I0(n8531[0]), .I1(n186), .CO(n25855));
    SB_LUT4 add_4440_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n8519[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n25854));
    SB_LUT4 add_4439_12_lut (.I0(GND_net), .I1(n8519[9]), .I2(GND_net), 
            .I3(n25853), .O(n8506[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_11_lut (.I0(GND_net), .I1(n8519[8]), .I2(GND_net), 
            .I3(n25852), .O(n8506[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n24767), .O(n103[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_11 (.CI(n25852), .I0(n8519[8]), .I1(GND_net), .CO(n25853));
    SB_LUT4 add_4439_10_lut (.I0(GND_net), .I1(n8519[7]), .I2(GND_net), 
            .I3(n25851), .O(n8506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_10 (.CI(n25851), .I0(n8519[7]), .I1(GND_net), .CO(n25852));
    SB_LUT4 add_4439_9_lut (.I0(GND_net), .I1(n8519[6]), .I2(GND_net), 
            .I3(n25850), .O(n8506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_20 (.CI(n24767), .I0(GND_net), .I1(n1[18]), 
            .CO(n24768));
    SB_CARRY add_4439_9 (.CI(n25850), .I0(n8519[6]), .I1(GND_net), .CO(n25851));
    SB_LUT4 add_4439_8_lut (.I0(GND_net), .I1(n8519[5]), .I2(n548), .I3(n25849), 
            .O(n8506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_8 (.CI(n25849), .I0(n8519[5]), .I1(n548), .CO(n25850));
    SB_LUT4 add_4439_7_lut (.I0(GND_net), .I1(n8519[4]), .I2(n475), .I3(n25848), 
            .O(n8506[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n24766), .O(n103[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_19 (.CI(n24766), .I0(GND_net), .I1(n1[17]), 
            .CO(n24767));
    SB_CARRY add_4439_7 (.CI(n25848), .I0(n8519[4]), .I1(n475), .CO(n25849));
    SB_LUT4 add_4439_6_lut (.I0(GND_net), .I1(n8519[3]), .I2(n402), .I3(n25847), 
            .O(n8506[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n24765), .O(n103[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_6 (.CI(n25847), .I0(n8519[3]), .I1(n402), .CO(n25848));
    SB_LUT4 add_4439_5_lut (.I0(GND_net), .I1(n8519[2]), .I2(n329), .I3(n25846), 
            .O(n8506[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_5 (.CI(n25846), .I0(n8519[2]), .I1(n329), .CO(n25847));
    SB_LUT4 add_4439_4_lut (.I0(GND_net), .I1(n8519[1]), .I2(n256), .I3(n25845), 
            .O(n8506[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_4 (.CI(n25845), .I0(n8519[1]), .I1(n256), .CO(n25846));
    SB_LUT4 add_4439_3_lut (.I0(GND_net), .I1(n8519[0]), .I2(n183), .I3(n25844), 
            .O(n8506[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_3 (.CI(n25844), .I0(n8519[0]), .I1(n183), .CO(n25845));
    SB_LUT4 add_4439_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n8506[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n25844));
    SB_LUT4 add_4438_13_lut (.I0(GND_net), .I1(n8506[10]), .I2(GND_net), 
            .I3(n25843), .O(n8492[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_12_lut (.I0(GND_net), .I1(n8506[9]), .I2(GND_net), 
            .I3(n25842), .O(n8492[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_12 (.CI(n25842), .I0(n8506[9]), .I1(GND_net), .CO(n25843));
    SB_LUT4 add_4438_11_lut (.I0(GND_net), .I1(n8506[8]), .I2(GND_net), 
            .I3(n25841), .O(n8492[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_11 (.CI(n25841), .I0(n8506[8]), .I1(GND_net), .CO(n25842));
    SB_LUT4 add_4438_10_lut (.I0(GND_net), .I1(n8506[7]), .I2(GND_net), 
            .I3(n25840), .O(n8492[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_10 (.CI(n25840), .I0(n8506[7]), .I1(GND_net), .CO(n25841));
    SB_LUT4 add_4438_9_lut (.I0(GND_net), .I1(n8506[6]), .I2(GND_net), 
            .I3(n25839), .O(n8492[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_9 (.CI(n25839), .I0(n8506[6]), .I1(GND_net), .CO(n25840));
    SB_LUT4 add_4438_8_lut (.I0(GND_net), .I1(n8506[5]), .I2(n545), .I3(n25838), 
            .O(n8492[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_8 (.CI(n25838), .I0(n8506[5]), .I1(n545), .CO(n25839));
    SB_LUT4 add_4438_7_lut (.I0(GND_net), .I1(n8506[4]), .I2(n472), .I3(n25837), 
            .O(n8492[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_7 (.CI(n25837), .I0(n8506[4]), .I1(n472), .CO(n25838));
    SB_LUT4 add_4438_6_lut (.I0(GND_net), .I1(n8506[3]), .I2(n399), .I3(n25836), 
            .O(n8492[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_6 (.CI(n25836), .I0(n8506[3]), .I1(n399), .CO(n25837));
    SB_LUT4 add_4438_5_lut (.I0(GND_net), .I1(n8506[2]), .I2(n326), .I3(n25835), 
            .O(n8492[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_5 (.CI(n25835), .I0(n8506[2]), .I1(n326), .CO(n25836));
    SB_LUT4 add_4438_4_lut (.I0(GND_net), .I1(n8506[1]), .I2(n253), .I3(n25834), 
            .O(n8492[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_4 (.CI(n25834), .I0(n8506[1]), .I1(n253), .CO(n25835));
    SB_LUT4 add_4438_3_lut (.I0(GND_net), .I1(n8506[0]), .I2(n180), .I3(n25833), 
            .O(n8492[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_3 (.CI(n25833), .I0(n8506[0]), .I1(n180), .CO(n25834));
    SB_LUT4 add_4438_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8492[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n25833));
    SB_LUT4 add_4437_14_lut (.I0(GND_net), .I1(n8492[11]), .I2(GND_net), 
            .I3(n25832), .O(n8477[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_13_lut (.I0(GND_net), .I1(n8492[10]), .I2(GND_net), 
            .I3(n25831), .O(n8477[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_13 (.CI(n25831), .I0(n8492[10]), .I1(GND_net), .CO(n25832));
    SB_LUT4 add_4437_12_lut (.I0(GND_net), .I1(n8492[9]), .I2(GND_net), 
            .I3(n25830), .O(n8477[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_12 (.CI(n25830), .I0(n8492[9]), .I1(GND_net), .CO(n25831));
    SB_LUT4 add_4437_11_lut (.I0(GND_net), .I1(n8492[8]), .I2(GND_net), 
            .I3(n25829), .O(n8477[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_11 (.CI(n25829), .I0(n8492[8]), .I1(GND_net), .CO(n25830));
    SB_LUT4 add_4437_10_lut (.I0(GND_net), .I1(n8492[7]), .I2(GND_net), 
            .I3(n25828), .O(n8477[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_18 (.CI(n24765), .I0(GND_net), .I1(n1[16]), 
            .CO(n24766));
    SB_CARRY add_4437_10 (.CI(n25828), .I0(n8492[7]), .I1(GND_net), .CO(n25829));
    SB_LUT4 add_4437_9_lut (.I0(GND_net), .I1(n8492[6]), .I2(GND_net), 
            .I3(n25827), .O(n8477[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_9 (.CI(n25827), .I0(n8492[6]), .I1(GND_net), .CO(n25828));
    SB_LUT4 add_4437_8_lut (.I0(GND_net), .I1(n8492[5]), .I2(n542), .I3(n25826), 
            .O(n8477[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_8 (.CI(n25826), .I0(n8492[5]), .I1(n542), .CO(n25827));
    SB_LUT4 add_4437_7_lut (.I0(GND_net), .I1(n8492[4]), .I2(n469), .I3(n25825), 
            .O(n8477[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_7 (.CI(n25825), .I0(n8492[4]), .I1(n469), .CO(n25826));
    SB_LUT4 add_4437_6_lut (.I0(GND_net), .I1(n8492[3]), .I2(n396), .I3(n25824), 
            .O(n8477[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_6 (.CI(n25824), .I0(n8492[3]), .I1(n396), .CO(n25825));
    SB_LUT4 unary_minus_8_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n24764), .O(n103[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_5_lut (.I0(GND_net), .I1(n8492[2]), .I2(n323), .I3(n25823), 
            .O(n8477[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_17 (.CI(n24764), .I0(GND_net), .I1(n1[15]), 
            .CO(n24765));
    SB_CARRY add_4437_5 (.CI(n25823), .I0(n8492[2]), .I1(n323), .CO(n25824));
    SB_LUT4 add_4437_4_lut (.I0(GND_net), .I1(n8492[1]), .I2(n250), .I3(n25822), 
            .O(n8477[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_4 (.CI(n25822), .I0(n8492[1]), .I1(n250), .CO(n25823));
    SB_LUT4 add_4437_3_lut (.I0(GND_net), .I1(n8492[0]), .I2(n177), .I3(n25821), 
            .O(n8477[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_3 (.CI(n25821), .I0(n8492[0]), .I1(n177), .CO(n25822));
    SB_LUT4 add_4437_2_lut (.I0(GND_net), .I1(n35_adj_3490), .I2(n104_adj_3491), 
            .I3(GND_net), .O(n8477[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_2 (.CI(GND_net), .I0(n35_adj_3490), .I1(n104_adj_3491), 
            .CO(n25821));
    SB_LUT4 add_4436_15_lut (.I0(GND_net), .I1(n8477[12]), .I2(GND_net), 
            .I3(n25820), .O(n8461[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_14_lut (.I0(GND_net), .I1(n8477[11]), .I2(GND_net), 
            .I3(n25819), .O(n8461[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n24763), .O(n103[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_14 (.CI(n25819), .I0(n8477[11]), .I1(GND_net), .CO(n25820));
    SB_LUT4 add_4436_13_lut (.I0(GND_net), .I1(n8477[10]), .I2(GND_net), 
            .I3(n25818), .O(n8461[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_13 (.CI(n25818), .I0(n8477[10]), .I1(GND_net), .CO(n25819));
    SB_LUT4 add_4436_12_lut (.I0(GND_net), .I1(n8477[9]), .I2(GND_net), 
            .I3(n25817), .O(n8461[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_12 (.CI(n25817), .I0(n8477[9]), .I1(GND_net), .CO(n25818));
    SB_LUT4 add_4436_11_lut (.I0(GND_net), .I1(n8477[8]), .I2(GND_net), 
            .I3(n25816), .O(n8461[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_11 (.CI(n25816), .I0(n8477[8]), .I1(GND_net), .CO(n25817));
    SB_LUT4 add_4436_10_lut (.I0(GND_net), .I1(n8477[7]), .I2(GND_net), 
            .I3(n25815), .O(n8461[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_10 (.CI(n25815), .I0(n8477[7]), .I1(GND_net), .CO(n25816));
    SB_LUT4 add_4436_9_lut (.I0(GND_net), .I1(n8477[6]), .I2(GND_net), 
            .I3(n25814), .O(n8461[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_9 (.CI(n25814), .I0(n8477[6]), .I1(GND_net), .CO(n25815));
    SB_CARRY unary_minus_8_add_3_16 (.CI(n24763), .I0(GND_net), .I1(n1[14]), 
            .CO(n24764));
    SB_LUT4 add_4436_8_lut (.I0(GND_net), .I1(n8477[5]), .I2(n539), .I3(n25813), 
            .O(n8461[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_8 (.CI(n25813), .I0(n8477[5]), .I1(n539), .CO(n25814));
    SB_LUT4 add_4436_7_lut (.I0(GND_net), .I1(n8477[4]), .I2(n466), .I3(n25812), 
            .O(n8461[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n24762), .O(n103[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_7 (.CI(n25812), .I0(n8477[4]), .I1(n466), .CO(n25813));
    SB_CARRY unary_minus_8_add_3_15 (.CI(n24762), .I0(GND_net), .I1(n1[13]), 
            .CO(n24763));
    SB_LUT4 add_4436_6_lut (.I0(GND_net), .I1(n8477[3]), .I2(n393), .I3(n25811), 
            .O(n8461[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_6 (.CI(n25811), .I0(n8477[3]), .I1(n393), .CO(n25812));
    SB_LUT4 unary_minus_8_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n24761), .O(n103[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_14 (.CI(n24761), .I0(GND_net), .I1(n1[12]), 
            .CO(n24762));
    SB_LUT4 add_4436_5_lut (.I0(GND_net), .I1(n8477[2]), .I2(n320), .I3(n25810), 
            .O(n8461[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n24760), .O(n103[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_13 (.CI(n24760), .I0(GND_net), .I1(n1[11]), 
            .CO(n24761));
    SB_LUT4 unary_minus_8_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n24759), .O(n103[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_12 (.CI(n24759), .I0(GND_net), .I1(n1[10]), 
            .CO(n24760));
    SB_CARRY add_4436_5 (.CI(n25810), .I0(n8477[2]), .I1(n320), .CO(n25811));
    SB_LUT4 unary_minus_8_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n24758), .O(n103[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_11 (.CI(n24758), .I0(GND_net), .I1(n1[9]), 
            .CO(n24759));
    SB_LUT4 unary_minus_8_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n24757), .O(n103[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_4_lut (.I0(GND_net), .I1(n8477[1]), .I2(n247), .I3(n25809), 
            .O(n8461[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_10 (.CI(n24757), .I0(GND_net), .I1(n1[8]), 
            .CO(n24758));
    SB_LUT4 unary_minus_8_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n24756), .O(n103[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_9 (.CI(n24756), .I0(GND_net), .I1(n1[7]), 
            .CO(n24757));
    SB_LUT4 unary_minus_8_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n24755), .O(n103[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_8 (.CI(n24755), .I0(GND_net), .I1(n1[6]), 
            .CO(n24756));
    SB_LUT4 unary_minus_8_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n24754), .O(n103[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_7 (.CI(n24754), .I0(GND_net), .I1(n1[5]), 
            .CO(n24755));
    SB_LUT4 unary_minus_8_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n24753), .O(n103[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_6 (.CI(n24753), .I0(GND_net), .I1(n1[4]), 
            .CO(n24754));
    SB_LUT4 unary_minus_8_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n24752), .O(n103[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_4 (.CI(n25809), .I0(n8477[1]), .I1(n247), .CO(n25810));
    SB_CARRY unary_minus_8_add_3_5 (.CI(n24752), .I0(GND_net), .I1(n1[3]), 
            .CO(n24753));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3291[1]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 unary_minus_8_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n24751), .O(n103[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_3_lut (.I0(GND_net), .I1(n8477[0]), .I2(n174), .I3(n25808), 
            .O(n8461[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_3 (.CI(n25808), .I0(n8477[0]), .I1(n174), .CO(n25809));
    SB_LUT4 add_4436_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8461[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n25808));
    SB_LUT4 add_4435_16_lut (.I0(GND_net), .I1(n8461[13]), .I2(GND_net), 
            .I3(n25807), .O(n8444[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_15_lut (.I0(GND_net), .I1(n8461[12]), .I2(GND_net), 
            .I3(n25806), .O(n8444[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_15 (.CI(n25806), .I0(n8461[12]), .I1(GND_net), .CO(n25807));
    SB_LUT4 add_4435_14_lut (.I0(GND_net), .I1(n8461[11]), .I2(GND_net), 
            .I3(n25805), .O(n8444[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_14 (.CI(n25805), .I0(n8461[11]), .I1(GND_net), .CO(n25806));
    SB_LUT4 add_4435_13_lut (.I0(GND_net), .I1(n8461[10]), .I2(GND_net), 
            .I3(n25804), .O(n8444[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_13 (.CI(n25804), .I0(n8461[10]), .I1(GND_net), .CO(n25805));
    SB_LUT4 add_4435_12_lut (.I0(GND_net), .I1(n8461[9]), .I2(GND_net), 
            .I3(n25803), .O(n8444[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_12 (.CI(n25803), .I0(n8461[9]), .I1(GND_net), .CO(n25804));
    SB_LUT4 add_4435_11_lut (.I0(GND_net), .I1(n8461[8]), .I2(GND_net), 
            .I3(n25802), .O(n8444[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_11 (.CI(n25802), .I0(n8461[8]), .I1(GND_net), .CO(n25803));
    SB_LUT4 add_4435_10_lut (.I0(GND_net), .I1(n8461[7]), .I2(GND_net), 
            .I3(n25801), .O(n8444[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_10 (.CI(n25801), .I0(n8461[7]), .I1(GND_net), .CO(n25802));
    SB_LUT4 add_4435_9_lut (.I0(GND_net), .I1(n8461[6]), .I2(GND_net), 
            .I3(n25800), .O(n8444[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_9 (.CI(n25800), .I0(n8461[6]), .I1(GND_net), .CO(n25801));
    SB_LUT4 add_4435_8_lut (.I0(GND_net), .I1(n8461[5]), .I2(n536), .I3(n25799), 
            .O(n8444[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_8 (.CI(n25799), .I0(n8461[5]), .I1(n536), .CO(n25800));
    SB_LUT4 add_4435_7_lut (.I0(GND_net), .I1(n8461[4]), .I2(n463), .I3(n25798), 
            .O(n8444[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_7 (.CI(n25798), .I0(n8461[4]), .I1(n463), .CO(n25799));
    SB_LUT4 add_4435_6_lut (.I0(GND_net), .I1(n8461[3]), .I2(n390), .I3(n25797), 
            .O(n8444[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_6 (.CI(n25797), .I0(n8461[3]), .I1(n390), .CO(n25798));
    SB_LUT4 add_4435_5_lut (.I0(GND_net), .I1(n8461[2]), .I2(n317), .I3(n25796), 
            .O(n8444[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_5 (.CI(n25796), .I0(n8461[2]), .I1(n317), .CO(n25797));
    SB_LUT4 add_4435_4_lut (.I0(GND_net), .I1(n8461[1]), .I2(n244), .I3(n25795), 
            .O(n8444[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_4 (.CI(n25795), .I0(n8461[1]), .I1(n244), .CO(n25796));
    SB_LUT4 add_4435_3_lut (.I0(GND_net), .I1(n8461[0]), .I2(n171), .I3(n25794), 
            .O(n8444[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_3 (.CI(n25794), .I0(n8461[0]), .I1(n171), .CO(n25795));
    SB_LUT4 add_4435_2_lut (.I0(GND_net), .I1(n29_adj_3506), .I2(n98), 
            .I3(GND_net), .O(n8444[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_2 (.CI(GND_net), .I0(n29_adj_3506), .I1(n98), .CO(n25794));
    SB_LUT4 add_4434_17_lut (.I0(GND_net), .I1(n8444[14]), .I2(GND_net), 
            .I3(n25793), .O(n8426[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_16_lut (.I0(GND_net), .I1(n8444[13]), .I2(GND_net), 
            .I3(n25792), .O(n8426[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_16 (.CI(n25792), .I0(n8444[13]), .I1(GND_net), .CO(n25793));
    SB_LUT4 add_4434_15_lut (.I0(GND_net), .I1(n8444[12]), .I2(GND_net), 
            .I3(n25791), .O(n8426[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_15 (.CI(n25791), .I0(n8444[12]), .I1(GND_net), .CO(n25792));
    SB_LUT4 add_4434_14_lut (.I0(GND_net), .I1(n8444[11]), .I2(GND_net), 
            .I3(n25790), .O(n8426[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_14 (.CI(n25790), .I0(n8444[11]), .I1(GND_net), .CO(n25791));
    SB_LUT4 add_4434_13_lut (.I0(GND_net), .I1(n8444[10]), .I2(GND_net), 
            .I3(n25789), .O(n8426[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_13 (.CI(n25789), .I0(n8444[10]), .I1(GND_net), .CO(n25790));
    SB_LUT4 add_4434_12_lut (.I0(GND_net), .I1(n8444[9]), .I2(GND_net), 
            .I3(n25788), .O(n8426[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_12 (.CI(n25788), .I0(n8444[9]), .I1(GND_net), .CO(n25789));
    SB_LUT4 add_4434_11_lut (.I0(GND_net), .I1(n8444[8]), .I2(GND_net), 
            .I3(n25787), .O(n8426[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_11 (.CI(n25787), .I0(n8444[8]), .I1(GND_net), .CO(n25788));
    SB_LUT4 add_4434_10_lut (.I0(GND_net), .I1(n8444[7]), .I2(GND_net), 
            .I3(n25786), .O(n8426[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_10 (.CI(n25786), .I0(n8444[7]), .I1(GND_net), .CO(n25787));
    SB_LUT4 add_4434_9_lut (.I0(GND_net), .I1(n8444[6]), .I2(GND_net), 
            .I3(n25785), .O(n8426[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_9 (.CI(n25785), .I0(n8444[6]), .I1(GND_net), .CO(n25786));
    SB_LUT4 add_4434_8_lut (.I0(GND_net), .I1(n8444[5]), .I2(n533), .I3(n25784), 
            .O(n8426[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_8 (.CI(n25784), .I0(n8444[5]), .I1(n533), .CO(n25785));
    SB_LUT4 add_4434_7_lut (.I0(GND_net), .I1(n8444[4]), .I2(n460), .I3(n25783), 
            .O(n8426[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_7 (.CI(n25783), .I0(n8444[4]), .I1(n460), .CO(n25784));
    SB_LUT4 add_4434_6_lut (.I0(GND_net), .I1(n8444[3]), .I2(n387), .I3(n25782), 
            .O(n8426[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_6 (.CI(n25782), .I0(n8444[3]), .I1(n387), .CO(n25783));
    SB_LUT4 add_4434_5_lut (.I0(GND_net), .I1(n8444[2]), .I2(n314), .I3(n25781), 
            .O(n8426[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_5 (.CI(n25781), .I0(n8444[2]), .I1(n314), .CO(n25782));
    SB_LUT4 add_4434_4_lut (.I0(GND_net), .I1(n8444[1]), .I2(n241), .I3(n25780), 
            .O(n8426[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_4 (.CI(n25780), .I0(n8444[1]), .I1(n241), .CO(n25781));
    SB_LUT4 add_4434_3_lut (.I0(GND_net), .I1(n8444[0]), .I2(n168), .I3(n25779), 
            .O(n8426[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_3 (.CI(n25779), .I0(n8444[0]), .I1(n168), .CO(n25780));
    SB_LUT4 add_4434_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n8426[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n25779));
    SB_LUT4 add_4433_18_lut (.I0(GND_net), .I1(n8426[15]), .I2(GND_net), 
            .I3(n25778), .O(n8407[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_17_lut (.I0(GND_net), .I1(n8426[14]), .I2(GND_net), 
            .I3(n25777), .O(n8407[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_17 (.CI(n25777), .I0(n8426[14]), .I1(GND_net), .CO(n25778));
    SB_LUT4 add_4433_16_lut (.I0(GND_net), .I1(n8426[13]), .I2(GND_net), 
            .I3(n25776), .O(n8407[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_16 (.CI(n25776), .I0(n8426[13]), .I1(GND_net), .CO(n25777));
    SB_LUT4 add_4433_15_lut (.I0(GND_net), .I1(n8426[12]), .I2(GND_net), 
            .I3(n25775), .O(n8407[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_15 (.CI(n25775), .I0(n8426[12]), .I1(GND_net), .CO(n25776));
    SB_LUT4 add_4433_14_lut (.I0(GND_net), .I1(n8426[11]), .I2(GND_net), 
            .I3(n25774), .O(n8407[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_14 (.CI(n25774), .I0(n8426[11]), .I1(GND_net), .CO(n25775));
    SB_LUT4 add_4433_13_lut (.I0(GND_net), .I1(n8426[10]), .I2(GND_net), 
            .I3(n25773), .O(n8407[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_13 (.CI(n25773), .I0(n8426[10]), .I1(GND_net), .CO(n25774));
    SB_LUT4 add_4433_12_lut (.I0(GND_net), .I1(n8426[9]), .I2(GND_net), 
            .I3(n25772), .O(n8407[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_12 (.CI(n25772), .I0(n8426[9]), .I1(GND_net), .CO(n25773));
    SB_LUT4 add_4433_11_lut (.I0(GND_net), .I1(n8426[8]), .I2(GND_net), 
            .I3(n25771), .O(n8407[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_11 (.CI(n25771), .I0(n8426[8]), .I1(GND_net), .CO(n25772));
    SB_LUT4 add_4433_10_lut (.I0(GND_net), .I1(n8426[7]), .I2(GND_net), 
            .I3(n25770), .O(n8407[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_10 (.CI(n25770), .I0(n8426[7]), .I1(GND_net), .CO(n25771));
    SB_LUT4 add_4433_9_lut (.I0(GND_net), .I1(n8426[6]), .I2(GND_net), 
            .I3(n25769), .O(n8407[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_9 (.CI(n25769), .I0(n8426[6]), .I1(GND_net), .CO(n25770));
    SB_LUT4 add_4433_8_lut (.I0(GND_net), .I1(n8426[5]), .I2(n530), .I3(n25768), 
            .O(n8407[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_8 (.CI(n25768), .I0(n8426[5]), .I1(n530), .CO(n25769));
    SB_LUT4 add_4433_7_lut (.I0(GND_net), .I1(n8426[4]), .I2(n457), .I3(n25767), 
            .O(n8407[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_7 (.CI(n25767), .I0(n8426[4]), .I1(n457), .CO(n25768));
    SB_LUT4 add_4433_6_lut (.I0(GND_net), .I1(n8426[3]), .I2(n384), .I3(n25766), 
            .O(n8407[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_6 (.CI(n25766), .I0(n8426[3]), .I1(n384), .CO(n25767));
    SB_LUT4 add_4433_5_lut (.I0(GND_net), .I1(n8426[2]), .I2(n311), .I3(n25765), 
            .O(n8407[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_5 (.CI(n25765), .I0(n8426[2]), .I1(n311), .CO(n25766));
    SB_LUT4 add_4433_4_lut (.I0(GND_net), .I1(n8426[1]), .I2(n238), .I3(n25764), 
            .O(n8407[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_4 (.CI(n25764), .I0(n8426[1]), .I1(n238), .CO(n25765));
    SB_LUT4 add_4433_3_lut (.I0(GND_net), .I1(n8426[0]), .I2(n165), .I3(n25763), 
            .O(n8407[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_3 (.CI(n25763), .I0(n8426[0]), .I1(n165), .CO(n25764));
    SB_LUT4 add_4433_2_lut (.I0(GND_net), .I1(n23_adj_3507), .I2(n92), 
            .I3(GND_net), .O(n8407[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_2 (.CI(GND_net), .I0(n23_adj_3507), .I1(n92), .CO(n25763));
    SB_LUT4 add_4432_19_lut (.I0(GND_net), .I1(n8407[16]), .I2(GND_net), 
            .I3(n25762), .O(n8387[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_18_lut (.I0(GND_net), .I1(n8407[15]), .I2(GND_net), 
            .I3(n25761), .O(n8387[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_18 (.CI(n25761), .I0(n8407[15]), .I1(GND_net), .CO(n25762));
    SB_LUT4 add_4432_17_lut (.I0(GND_net), .I1(n8407[14]), .I2(GND_net), 
            .I3(n25760), .O(n8387[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_17 (.CI(n25760), .I0(n8407[14]), .I1(GND_net), .CO(n25761));
    SB_LUT4 add_4432_16_lut (.I0(GND_net), .I1(n8407[13]), .I2(GND_net), 
            .I3(n25759), .O(n8387[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_16 (.CI(n25759), .I0(n8407[13]), .I1(GND_net), .CO(n25760));
    SB_LUT4 add_4432_15_lut (.I0(GND_net), .I1(n8407[12]), .I2(GND_net), 
            .I3(n25758), .O(n8387[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_15 (.CI(n25758), .I0(n8407[12]), .I1(GND_net), .CO(n25759));
    SB_LUT4 add_4432_14_lut (.I0(GND_net), .I1(n8407[11]), .I2(GND_net), 
            .I3(n25757), .O(n8387[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_14 (.CI(n25757), .I0(n8407[11]), .I1(GND_net), .CO(n25758));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3291[2]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 add_4432_13_lut (.I0(GND_net), .I1(n8407[10]), .I2(GND_net), 
            .I3(n25756), .O(n8387[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3291[3]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3291[4]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3291[5]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3291[6]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3291[7]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3291[8]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3291[9]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3291[10]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3291[11]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3291[12]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3291[13]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3291[14]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3291[15]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3291[16]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3291[17]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3291[18]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3291[19]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3291[20]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3291[21]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3291[22]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3291[23]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [1]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [2]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [3]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [4]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [5]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [6]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [7]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [8]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [9]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [10]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [11]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [12]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [13]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [14]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [15]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [16]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [17]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [18]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [19]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [20]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [21]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [22]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3315 [23]));   // verilog/motorControl.v(36[14] 55[8])
    SB_CARRY add_4432_13 (.CI(n25756), .I0(n8407[10]), .I1(GND_net), .CO(n25757));
    SB_LUT4 add_4432_12_lut (.I0(GND_net), .I1(n8407[9]), .I2(GND_net), 
            .I3(n25755), .O(n8387[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_12 (.CI(n25755), .I0(n8407[9]), .I1(GND_net), .CO(n25756));
    SB_LUT4 add_4432_11_lut (.I0(GND_net), .I1(n8407[8]), .I2(GND_net), 
            .I3(n25754), .O(n8387[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_11 (.CI(n25754), .I0(n8407[8]), .I1(GND_net), .CO(n25755));
    SB_LUT4 add_4432_10_lut (.I0(GND_net), .I1(n8407[7]), .I2(GND_net), 
            .I3(n25753), .O(n8387[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_10 (.CI(n25753), .I0(n8407[7]), .I1(GND_net), .CO(n25754));
    SB_LUT4 add_4432_9_lut (.I0(GND_net), .I1(n8407[6]), .I2(GND_net), 
            .I3(n25752), .O(n8387[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_9 (.CI(n25752), .I0(n8407[6]), .I1(GND_net), .CO(n25753));
    SB_LUT4 add_4432_8_lut (.I0(GND_net), .I1(n8407[5]), .I2(n527), .I3(n25751), 
            .O(n8387[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_8 (.CI(n25751), .I0(n8407[5]), .I1(n527), .CO(n25752));
    SB_LUT4 add_4432_7_lut (.I0(GND_net), .I1(n8407[4]), .I2(n454), .I3(n25750), 
            .O(n8387[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_7 (.CI(n25750), .I0(n8407[4]), .I1(n454), .CO(n25751));
    SB_LUT4 i29202_3_lut_4_lut (.I0(duty[3]), .I1(n103[3]), .I2(n103[2]), 
            .I3(duty[2]), .O(n34839));   // verilog/motorControl.v(45[19:35])
    defparam i29202_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_4432_6_lut (.I0(GND_net), .I1(n8407[3]), .I2(n381), .I3(n25749), 
            .O(n8387[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_6 (.CI(n25749), .I0(n8407[3]), .I1(n381), .CO(n25750));
    SB_LUT4 add_4432_5_lut (.I0(GND_net), .I1(n8407[2]), .I2(n308), .I3(n25748), 
            .O(n8387[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_5 (.CI(n25748), .I0(n8407[2]), .I1(n308), .CO(n25749));
    SB_LUT4 add_4432_4_lut (.I0(GND_net), .I1(n8407[1]), .I2(n235), .I3(n25747), 
            .O(n8387[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_4 (.CI(n25747), .I0(n8407[1]), .I1(n235), .CO(n25748));
    SB_LUT4 add_4432_3_lut (.I0(GND_net), .I1(n8407[0]), .I2(n162), .I3(n25746), 
            .O(n8387[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_3 (.CI(n25746), .I0(n8407[0]), .I1(n162), .CO(n25747));
    SB_LUT4 add_4432_2_lut (.I0(GND_net), .I1(n20_adj_3508), .I2(n89), 
            .I3(GND_net), .O(n8387[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_2 (.CI(GND_net), .I0(n20_adj_3508), .I1(n89), .CO(n25746));
    SB_LUT4 add_4431_20_lut (.I0(GND_net), .I1(n8387[17]), .I2(GND_net), 
            .I3(n25745), .O(n8366[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_19_lut (.I0(GND_net), .I1(n8387[16]), .I2(GND_net), 
            .I3(n25744), .O(n8366[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_19 (.CI(n25744), .I0(n8387[16]), .I1(GND_net), .CO(n25745));
    SB_LUT4 add_4431_18_lut (.I0(GND_net), .I1(n8387[15]), .I2(GND_net), 
            .I3(n25743), .O(n8366[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_4 (.CI(n24751), .I0(GND_net), .I1(n1[2]), 
            .CO(n24752));
    SB_CARRY add_4431_18 (.CI(n25743), .I0(n8387[15]), .I1(GND_net), .CO(n25744));
    SB_LUT4 add_4431_17_lut (.I0(GND_net), .I1(n8387[14]), .I2(GND_net), 
            .I3(n25742), .O(n8366[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_17 (.CI(n25742), .I0(n8387[14]), .I1(GND_net), .CO(n25743));
    SB_LUT4 add_4431_16_lut (.I0(GND_net), .I1(n8387[13]), .I2(GND_net), 
            .I3(n25741), .O(n8366[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_16 (.CI(n25741), .I0(n8387[13]), .I1(GND_net), .CO(n25742));
    SB_LUT4 add_4431_15_lut (.I0(GND_net), .I1(n8387[12]), .I2(GND_net), 
            .I3(n25740), .O(n8366[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_15 (.CI(n25740), .I0(n8387[12]), .I1(GND_net), .CO(n25741));
    SB_LUT4 add_4431_14_lut (.I0(GND_net), .I1(n8387[11]), .I2(GND_net), 
            .I3(n25739), .O(n8366[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_14 (.CI(n25739), .I0(n8387[11]), .I1(GND_net), .CO(n25740));
    SB_LUT4 add_4431_13_lut (.I0(GND_net), .I1(n8387[10]), .I2(GND_net), 
            .I3(n25738), .O(n8366[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_13 (.CI(n25738), .I0(n8387[10]), .I1(GND_net), .CO(n25739));
    SB_LUT4 add_4431_12_lut (.I0(GND_net), .I1(n8387[9]), .I2(GND_net), 
            .I3(n25737), .O(n8366[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_12 (.CI(n25737), .I0(n8387[9]), .I1(GND_net), .CO(n25738));
    SB_LUT4 add_4431_11_lut (.I0(GND_net), .I1(n8387[8]), .I2(GND_net), 
            .I3(n25736), .O(n8366[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_11 (.CI(n25736), .I0(n8387[8]), .I1(GND_net), .CO(n25737));
    SB_LUT4 add_4431_10_lut (.I0(GND_net), .I1(n8387[7]), .I2(GND_net), 
            .I3(n25735), .O(n8366[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_10 (.CI(n25735), .I0(n8387[7]), .I1(GND_net), .CO(n25736));
    SB_LUT4 add_4431_9_lut (.I0(GND_net), .I1(n8387[6]), .I2(GND_net), 
            .I3(n25734), .O(n8366[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_9 (.CI(n25734), .I0(n8387[6]), .I1(GND_net), .CO(n25735));
    SB_LUT4 add_4431_8_lut (.I0(GND_net), .I1(n8387[5]), .I2(n524), .I3(n25733), 
            .O(n8366[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_8 (.CI(n25733), .I0(n8387[5]), .I1(n524), .CO(n25734));
    SB_LUT4 add_4431_7_lut (.I0(GND_net), .I1(n8387[4]), .I2(n451), .I3(n25732), 
            .O(n8366[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_7 (.CI(n25732), .I0(n8387[4]), .I1(n451), .CO(n25733));
    SB_LUT4 add_4431_6_lut (.I0(GND_net), .I1(n8387[3]), .I2(n378), .I3(n25731), 
            .O(n8366[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_6 (.CI(n25731), .I0(n8387[3]), .I1(n378), .CO(n25732));
    SB_LUT4 add_4431_5_lut (.I0(GND_net), .I1(n8387[2]), .I2(n305), .I3(n25730), 
            .O(n8366[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_5 (.CI(n25730), .I0(n8387[2]), .I1(n305), .CO(n25731));
    SB_LUT4 add_4431_4_lut (.I0(GND_net), .I1(n8387[1]), .I2(n232), .I3(n25729), 
            .O(n8366[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_4 (.CI(n25729), .I0(n8387[1]), .I1(n232), .CO(n25730));
    SB_LUT4 LessThan_7_i6_3_lut_3_lut (.I0(duty[3]), .I1(n103[3]), .I2(n103[2]), 
            .I3(GND_net), .O(n6_adj_3469));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_4431_3_lut (.I0(GND_net), .I1(n8387[0]), .I2(n159), .I3(n25728), 
            .O(n8366[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_3 (.CI(n25728), .I0(n8387[0]), .I1(n159), .CO(n25729));
    SB_LUT4 add_4431_2_lut (.I0(GND_net), .I1(n17_adj_3509), .I2(n86), 
            .I3(GND_net), .O(n8366[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20162_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_3510), .I3(n8576[1]), .O(n6_adj_3430));   // verilog/motorControl.v(41[17:23])
    defparam i20162_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_4431_2 (.CI(GND_net), .I0(n17_adj_3509), .I1(n86), .CO(n25728));
    SB_LUT4 add_4430_21_lut (.I0(GND_net), .I1(n8366[18]), .I2(GND_net), 
            .I3(n25727), .O(n8344[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_20_lut (.I0(GND_net), .I1(n8366[17]), .I2(GND_net), 
            .I3(n25726), .O(n8344[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_20 (.CI(n25726), .I0(n8366[17]), .I1(GND_net), .CO(n25727));
    SB_LUT4 add_4430_19_lut (.I0(GND_net), .I1(n8366[16]), .I2(GND_net), 
            .I3(n25725), .O(n8344[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_19 (.CI(n25725), .I0(n8366[16]), .I1(GND_net), .CO(n25726));
    SB_LUT4 add_4430_18_lut (.I0(GND_net), .I1(n8366[15]), .I2(GND_net), 
            .I3(n25724), .O(n8344[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_18 (.CI(n25724), .I0(n8366[15]), .I1(GND_net), .CO(n25725));
    SB_LUT4 add_4430_17_lut (.I0(GND_net), .I1(n8366[14]), .I2(GND_net), 
            .I3(n25723), .O(n8344[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_17 (.CI(n25723), .I0(n8366[14]), .I1(GND_net), .CO(n25724));
    SB_LUT4 add_4430_16_lut (.I0(GND_net), .I1(n8366[13]), .I2(GND_net), 
            .I3(n25722), .O(n8344[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_16 (.CI(n25722), .I0(n8366[13]), .I1(GND_net), .CO(n25723));
    SB_LUT4 add_4430_15_lut (.I0(GND_net), .I1(n8366[12]), .I2(GND_net), 
            .I3(n25721), .O(n8344[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_15 (.CI(n25721), .I0(n8366[12]), .I1(GND_net), .CO(n25722));
    SB_LUT4 add_4430_14_lut (.I0(GND_net), .I1(n8366[11]), .I2(GND_net), 
            .I3(n25720), .O(n8344[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_14 (.CI(n25720), .I0(n8366[11]), .I1(GND_net), .CO(n25721));
    SB_LUT4 add_4430_13_lut (.I0(GND_net), .I1(n8366[10]), .I2(GND_net), 
            .I3(n25719), .O(n8344[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_13 (.CI(n25719), .I0(n8366[10]), .I1(GND_net), .CO(n25720));
    SB_LUT4 add_4430_12_lut (.I0(GND_net), .I1(n8366[9]), .I2(GND_net), 
            .I3(n25718), .O(n8344[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_12 (.CI(n25718), .I0(n8366[9]), .I1(GND_net), .CO(n25719));
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8576[1]), .I3(n4_adj_3510), .O(n8569[2]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 add_4430_11_lut (.I0(GND_net), .I1(n8366[8]), .I2(GND_net), 
            .I3(n25717), .O(n8344[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_11 (.CI(n25717), .I0(n8366[8]), .I1(GND_net), .CO(n25718));
    SB_LUT4 add_4430_10_lut (.I0(GND_net), .I1(n8366[7]), .I2(GND_net), 
            .I3(n25716), .O(n8344[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_10 (.CI(n25716), .I0(n8366[7]), .I1(GND_net), .CO(n25717));
    SB_LUT4 add_4430_9_lut (.I0(GND_net), .I1(n8366[6]), .I2(GND_net), 
            .I3(n25715), .O(n8344[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_9 (.CI(n25715), .I0(n8366[6]), .I1(GND_net), .CO(n25716));
    SB_LUT4 add_4430_8_lut (.I0(GND_net), .I1(n8366[5]), .I2(n521), .I3(n25714), 
            .O(n8344[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_8 (.CI(n25714), .I0(n8366[5]), .I1(n521), .CO(n25715));
    SB_LUT4 add_4430_7_lut (.I0(GND_net), .I1(n8366[4]), .I2(n448), .I3(n25713), 
            .O(n8344[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_7 (.CI(n25713), .I0(n8366[4]), .I1(n448), .CO(n25714));
    SB_LUT4 add_4430_6_lut (.I0(GND_net), .I1(n8366[3]), .I2(n375), .I3(n25712), 
            .O(n8344[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_6 (.CI(n25712), .I0(n8366[3]), .I1(n375), .CO(n25713));
    SB_LUT4 add_4430_5_lut (.I0(GND_net), .I1(n8366[2]), .I2(n302), .I3(n25711), 
            .O(n8344[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_5 (.CI(n25711), .I0(n8366[2]), .I1(n302), .CO(n25712));
    SB_LUT4 add_4430_4_lut (.I0(GND_net), .I1(n8366[1]), .I2(n229), .I3(n25710), 
            .O(n8344[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_4 (.CI(n25710), .I0(n8366[1]), .I1(n229), .CO(n25711));
    SB_LUT4 add_4430_3_lut (.I0(GND_net), .I1(n8366[0]), .I2(n156), .I3(n25709), 
            .O(n8344[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_3 (.CI(n25709), .I0(n8366[0]), .I1(n156), .CO(n25710));
    SB_LUT4 add_4430_2_lut (.I0(GND_net), .I1(n14_adj_3511), .I2(n83), 
            .I3(GND_net), .O(n8344[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_2 (.CI(GND_net), .I0(n14_adj_3511), .I1(n83), .CO(n25709));
    SB_LUT4 add_4429_22_lut (.I0(GND_net), .I1(n8344[19]), .I2(GND_net), 
            .I3(n25708), .O(n8321[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_21_lut (.I0(GND_net), .I1(n8344[18]), .I2(GND_net), 
            .I3(n25707), .O(n8321[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_21 (.CI(n25707), .I0(n8344[18]), .I1(GND_net), .CO(n25708));
    SB_LUT4 add_4429_20_lut (.I0(GND_net), .I1(n8344[17]), .I2(GND_net), 
            .I3(n25706), .O(n8321[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_20 (.CI(n25706), .I0(n8344[17]), .I1(GND_net), .CO(n25707));
    SB_LUT4 add_4429_19_lut (.I0(GND_net), .I1(n8344[16]), .I2(GND_net), 
            .I3(n25705), .O(n8321[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_19 (.CI(n25705), .I0(n8344[16]), .I1(GND_net), .CO(n25706));
    SB_LUT4 add_4429_18_lut (.I0(GND_net), .I1(n8344[15]), .I2(GND_net), 
            .I3(n25704), .O(n8321[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_18 (.CI(n25704), .I0(n8344[15]), .I1(GND_net), .CO(n25705));
    SB_LUT4 add_4429_17_lut (.I0(GND_net), .I1(n8344[14]), .I2(GND_net), 
            .I3(n25703), .O(n8321[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_17 (.CI(n25703), .I0(n8344[14]), .I1(GND_net), .CO(n25704));
    SB_LUT4 add_4429_16_lut (.I0(GND_net), .I1(n8344[13]), .I2(GND_net), 
            .I3(n25702), .O(n8321[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_16 (.CI(n25702), .I0(n8344[13]), .I1(GND_net), .CO(n25703));
    SB_LUT4 add_4429_15_lut (.I0(GND_net), .I1(n8344[12]), .I2(GND_net), 
            .I3(n25701), .O(n8321[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_15 (.CI(n25701), .I0(n8344[12]), .I1(GND_net), .CO(n25702));
    SB_LUT4 add_4429_14_lut (.I0(GND_net), .I1(n8344[11]), .I2(GND_net), 
            .I3(n25700), .O(n8321[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_14 (.CI(n25700), .I0(n8344[11]), .I1(GND_net), .CO(n25701));
    SB_LUT4 add_4429_13_lut (.I0(GND_net), .I1(n8344[10]), .I2(GND_net), 
            .I3(n25699), .O(n8321[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_13 (.CI(n25699), .I0(n8344[10]), .I1(GND_net), .CO(n25700));
    SB_LUT4 add_4429_12_lut (.I0(GND_net), .I1(n8344[9]), .I2(GND_net), 
            .I3(n25698), .O(n8321[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_12 (.CI(n25698), .I0(n8344[9]), .I1(GND_net), .CO(n25699));
    SB_LUT4 add_4429_11_lut (.I0(GND_net), .I1(n8344[8]), .I2(GND_net), 
            .I3(n25697), .O(n8321[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_11 (.CI(n25697), .I0(n8344[8]), .I1(GND_net), .CO(n25698));
    SB_LUT4 add_4429_10_lut (.I0(GND_net), .I1(n8344[7]), .I2(GND_net), 
            .I3(n25696), .O(n8321[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_10 (.CI(n25696), .I0(n8344[7]), .I1(GND_net), .CO(n25697));
    SB_LUT4 add_4429_9_lut (.I0(GND_net), .I1(n8344[6]), .I2(GND_net), 
            .I3(n25695), .O(n8321[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_9 (.CI(n25695), .I0(n8344[6]), .I1(GND_net), .CO(n25696));
    SB_LUT4 add_4429_8_lut (.I0(GND_net), .I1(n8344[5]), .I2(n518), .I3(n25694), 
            .O(n8321[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_8 (.CI(n25694), .I0(n8344[5]), .I1(n518), .CO(n25695));
    SB_LUT4 add_4429_7_lut (.I0(GND_net), .I1(n8344[4]), .I2(n445), .I3(n25693), 
            .O(n8321[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_7 (.CI(n25693), .I0(n8344[4]), .I1(n445), .CO(n25694));
    SB_LUT4 i2_3_lut_4_lut_adj_842 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8576[0]), .I3(n24463), .O(n8569[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut_adj_842.LUT_INIT = 16'h8778;
    SB_LUT4 add_4429_6_lut (.I0(GND_net), .I1(n8344[3]), .I2(n372), .I3(n25692), 
            .O(n8321[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_6 (.CI(n25692), .I0(n8344[3]), .I1(n372), .CO(n25693));
    SB_LUT4 add_4429_5_lut (.I0(GND_net), .I1(n8344[2]), .I2(n299), .I3(n25691), 
            .O(n8321[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_5 (.CI(n25691), .I0(n8344[2]), .I1(n299), .CO(n25692));
    SB_LUT4 add_4429_4_lut (.I0(GND_net), .I1(n8344[1]), .I2(n226), .I3(n25690), 
            .O(n8321[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_4 (.CI(n25690), .I0(n8344[1]), .I1(n226), .CO(n25691));
    SB_LUT4 add_4429_3_lut (.I0(GND_net), .I1(n8344[0]), .I2(n153), .I3(n25689), 
            .O(n8321[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_3 (.CI(n25689), .I0(n8344[0]), .I1(n153), .CO(n25690));
    SB_LUT4 add_4429_2_lut (.I0(GND_net), .I1(n11_adj_3512), .I2(n80), 
            .I3(GND_net), .O(n8321[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_2 (.CI(GND_net), .I0(n11_adj_3512), .I1(n80), .CO(n25689));
    SB_LUT4 mult_4_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n8297[21]), 
            .I2(GND_net), .I3(n25688), .O(n34262)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_4_add_1225_23_lut (.I0(GND_net), .I1(n8297[20]), .I2(GND_net), 
            .I3(n25687), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_23 (.CI(n25687), .I0(n8297[20]), .I1(GND_net), 
            .CO(n25688));
    SB_LUT4 mult_4_add_1225_22_lut (.I0(GND_net), .I1(n8297[19]), .I2(GND_net), 
            .I3(n25686), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_22 (.CI(n25686), .I0(n8297[19]), .I1(GND_net), 
            .CO(n25687));
    SB_LUT4 mult_4_add_1225_21_lut (.I0(GND_net), .I1(n8297[18]), .I2(GND_net), 
            .I3(n25685), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_21 (.CI(n25685), .I0(n8297[18]), .I1(GND_net), 
            .CO(n25686));
    SB_LUT4 mult_4_add_1225_20_lut (.I0(GND_net), .I1(n8297[17]), .I2(GND_net), 
            .I3(n25684), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_20 (.CI(n25684), .I0(n8297[17]), .I1(GND_net), 
            .CO(n25685));
    SB_LUT4 mult_4_add_1225_19_lut (.I0(GND_net), .I1(n8297[16]), .I2(GND_net), 
            .I3(n25683), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_19 (.CI(n25683), .I0(n8297[16]), .I1(GND_net), 
            .CO(n25684));
    SB_LUT4 mult_4_add_1225_18_lut (.I0(GND_net), .I1(n8297[15]), .I2(GND_net), 
            .I3(n25682), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_18 (.CI(n25682), .I0(n8297[15]), .I1(GND_net), 
            .CO(n25683));
    SB_LUT4 mult_4_add_1225_17_lut (.I0(GND_net), .I1(n8297[14]), .I2(GND_net), 
            .I3(n25681), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_17 (.CI(n25681), .I0(n8297[14]), .I1(GND_net), 
            .CO(n25682));
    SB_LUT4 mult_4_add_1225_16_lut (.I0(GND_net), .I1(n8297[13]), .I2(GND_net), 
            .I3(n25680), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_16 (.CI(n25680), .I0(n8297[13]), .I1(GND_net), 
            .CO(n25681));
    SB_LUT4 mult_4_add_1225_15_lut (.I0(GND_net), .I1(n8297[12]), .I2(GND_net), 
            .I3(n25679), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_15 (.CI(n25679), .I0(n8297[12]), .I1(GND_net), 
            .CO(n25680));
    SB_LUT4 mult_4_add_1225_14_lut (.I0(GND_net), .I1(n8297[11]), .I2(GND_net), 
            .I3(n25678), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_14 (.CI(n25678), .I0(n8297[11]), .I1(GND_net), 
            .CO(n25679));
    SB_LUT4 mult_4_add_1225_13_lut (.I0(GND_net), .I1(n8297[10]), .I2(GND_net), 
            .I3(n25677), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_13 (.CI(n25677), .I0(n8297[10]), .I1(GND_net), 
            .CO(n25678));
    SB_LUT4 mult_4_add_1225_12_lut (.I0(GND_net), .I1(n8297[9]), .I2(GND_net), 
            .I3(n25676), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n24750), .O(n103[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_12 (.CI(n25676), .I0(n8297[9]), .I1(GND_net), 
            .CO(n25677));
    SB_LUT4 mult_4_add_1225_11_lut (.I0(GND_net), .I1(n8297[8]), .I2(GND_net), 
            .I3(n25675), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_11 (.CI(n25675), .I0(n8297[8]), .I1(GND_net), 
            .CO(n25676));
    SB_LUT4 mult_4_add_1225_10_lut (.I0(GND_net), .I1(n8297[7]), .I2(GND_net), 
            .I3(n25674), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_10 (.CI(n25674), .I0(n8297[7]), .I1(GND_net), 
            .CO(n25675));
    SB_LUT4 mult_4_add_1225_9_lut (.I0(GND_net), .I1(n8297[6]), .I2(GND_net), 
            .I3(n25673), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_9 (.CI(n25673), .I0(n8297[6]), .I1(GND_net), 
            .CO(n25674));
    SB_LUT4 mult_4_add_1225_8_lut (.I0(GND_net), .I1(n8297[5]), .I2(n512), 
            .I3(n25672), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_8 (.CI(n25672), .I0(n8297[5]), .I1(n512), 
            .CO(n25673));
    SB_LUT4 mult_4_add_1225_7_lut (.I0(GND_net), .I1(n8297[4]), .I2(n439), 
            .I3(n25671), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_7 (.CI(n25671), .I0(n8297[4]), .I1(n439), 
            .CO(n25672));
    SB_LUT4 mult_4_add_1225_6_lut (.I0(GND_net), .I1(n8297[3]), .I2(n366), 
            .I3(n25670), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_6 (.CI(n25670), .I0(n8297[3]), .I1(n366), 
            .CO(n25671));
    SB_LUT4 mult_4_add_1225_5_lut (.I0(GND_net), .I1(n8297[2]), .I2(n293), 
            .I3(n25669), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31221_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36858));   // verilog/motorControl.v(36[14] 55[8])
    defparam i31221_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_4_add_1225_5 (.CI(n25669), .I0(n8297[2]), .I1(n293), 
            .CO(n25670));
    SB_LUT4 mult_4_add_1225_4_lut (.I0(GND_net), .I1(n8297[1]), .I2(n220), 
            .I3(n25668), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_4 (.CI(n25668), .I0(n8297[1]), .I1(n220), 
            .CO(n25669));
    SB_LUT4 mult_4_add_1225_3_lut (.I0(GND_net), .I1(n8297[0]), .I2(n147), 
            .I3(n25667), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_3 (.CI(n25667), .I0(n8297[0]), .I1(n147), 
            .CO(n25668));
    SB_LUT4 mult_4_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3517), .I2(n74_adj_3518), 
            .I3(GND_net), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_2 (.CI(GND_net), .I0(n5_adj_3517), .I1(n74_adj_3518), 
            .CO(n25667));
    SB_LUT4 add_4428_23_lut (.I0(GND_net), .I1(n8321[20]), .I2(GND_net), 
            .I3(n25666), .O(n8297[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_22_lut (.I0(GND_net), .I1(n8321[19]), .I2(GND_net), 
            .I3(n25665), .O(n8297[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_22 (.CI(n25665), .I0(n8321[19]), .I1(GND_net), .CO(n25666));
    SB_LUT4 add_4428_21_lut (.I0(GND_net), .I1(n8321[18]), .I2(GND_net), 
            .I3(n25664), .O(n8297[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_21 (.CI(n25664), .I0(n8321[18]), .I1(GND_net), .CO(n25665));
    SB_LUT4 add_4428_20_lut (.I0(GND_net), .I1(n8321[17]), .I2(GND_net), 
            .I3(n25663), .O(n8297[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_20 (.CI(n25663), .I0(n8321[17]), .I1(GND_net), .CO(n25664));
    SB_LUT4 add_4428_19_lut (.I0(GND_net), .I1(n8321[16]), .I2(GND_net), 
            .I3(n25662), .O(n8297[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_19 (.CI(n25662), .I0(n8321[16]), .I1(GND_net), .CO(n25663));
    SB_LUT4 add_4428_18_lut (.I0(GND_net), .I1(n8321[15]), .I2(GND_net), 
            .I3(n25661), .O(n8297[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_18 (.CI(n25661), .I0(n8321[15]), .I1(GND_net), .CO(n25662));
    SB_LUT4 add_4428_17_lut (.I0(GND_net), .I1(n8321[14]), .I2(GND_net), 
            .I3(n25660), .O(n8297[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_17 (.CI(n25660), .I0(n8321[14]), .I1(GND_net), .CO(n25661));
    SB_LUT4 add_4428_16_lut (.I0(GND_net), .I1(n8321[13]), .I2(GND_net), 
            .I3(n25659), .O(n8297[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_16 (.CI(n25659), .I0(n8321[13]), .I1(GND_net), .CO(n25660));
    SB_LUT4 add_4428_15_lut (.I0(GND_net), .I1(n8321[12]), .I2(GND_net), 
            .I3(n25658), .O(n8297[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20154_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n24463), .I3(n8576[0]), .O(n4_adj_3510));   // verilog/motorControl.v(41[17:23])
    defparam i20154_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_4428_15 (.CI(n25658), .I0(n8321[12]), .I1(GND_net), .CO(n25659));
    SB_LUT4 add_4428_14_lut (.I0(GND_net), .I1(n8321[11]), .I2(GND_net), 
            .I3(n25657), .O(n8297[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_14 (.CI(n25657), .I0(n8321[11]), .I1(GND_net), .CO(n25658));
    SB_LUT4 add_4428_13_lut (.I0(GND_net), .I1(n8321[10]), .I2(GND_net), 
            .I3(n25656), .O(n8297[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_13 (.CI(n25656), .I0(n8321[10]), .I1(GND_net), .CO(n25657));
    SB_LUT4 add_4428_12_lut (.I0(GND_net), .I1(n8321[9]), .I2(GND_net), 
            .I3(n25655), .O(n8297[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_12 (.CI(n25655), .I0(n8321[9]), .I1(GND_net), .CO(n25656));
    SB_LUT4 add_4428_11_lut (.I0(GND_net), .I1(n8321[8]), .I2(GND_net), 
            .I3(n25654), .O(n8297[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_11 (.CI(n25654), .I0(n8321[8]), .I1(GND_net), .CO(n25655));
    SB_LUT4 add_4428_10_lut (.I0(GND_net), .I1(n8321[7]), .I2(GND_net), 
            .I3(n25653), .O(n8297[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_10 (.CI(n25653), .I0(n8321[7]), .I1(GND_net), .CO(n25654));
    SB_LUT4 add_4428_9_lut (.I0(GND_net), .I1(n8321[6]), .I2(GND_net), 
            .I3(n25652), .O(n8297[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_9 (.CI(n25652), .I0(n8321[6]), .I1(GND_net), .CO(n25653));
    SB_LUT4 add_4428_8_lut (.I0(GND_net), .I1(n8321[5]), .I2(n515), .I3(n25651), 
            .O(n8297[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_8 (.CI(n25651), .I0(n8321[5]), .I1(n515), .CO(n25652));
    SB_LUT4 add_4428_7_lut (.I0(GND_net), .I1(n8321[4]), .I2(n442), .I3(n25650), 
            .O(n8297[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_7 (.CI(n25650), .I0(n8321[4]), .I1(n442), .CO(n25651));
    SB_LUT4 add_4428_6_lut (.I0(GND_net), .I1(n8321[3]), .I2(n369), .I3(n25649), 
            .O(n8297[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_6 (.CI(n25649), .I0(n8321[3]), .I1(n369), .CO(n25650));
    SB_LUT4 add_4428_5_lut (.I0(GND_net), .I1(n8321[2]), .I2(n296), .I3(n25648), 
            .O(n8297[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_5 (.CI(n25648), .I0(n8321[2]), .I1(n296), .CO(n25649));
    SB_LUT4 add_4428_4_lut (.I0(GND_net), .I1(n8321[1]), .I2(n223), .I3(n25647), 
            .O(n8297[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_4 (.CI(n25647), .I0(n8321[1]), .I1(n223), .CO(n25648));
    SB_LUT4 add_4428_3_lut (.I0(GND_net), .I1(n8321[0]), .I2(n150), .I3(n25646), 
            .O(n8297[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_3 (.CI(n25646), .I0(n8321[0]), .I1(n150), .CO(n25647));
    SB_LUT4 add_4428_2_lut (.I0(GND_net), .I1(n8_adj_3519), .I2(n77), 
            .I3(GND_net), .O(n8297[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_2 (.CI(GND_net), .I0(n8_adj_3519), .I1(n77), .CO(n25646));
    SB_CARRY unary_minus_8_add_3_3 (.CI(n24750), .I0(GND_net), .I1(n1[1]), 
            .CO(n24751));
    SB_LUT4 unary_minus_8_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n103[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20143_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n24463));   // verilog/motorControl.v(41[17:23])
    defparam i20143_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20141_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8569[0]));   // verilog/motorControl.v(41[17:23])
    defparam i20141_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY unary_minus_8_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n24750));
    SB_LUT4 i20224_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n24540), .I3(n8587[0]), .O(n4_adj_3455));   // verilog/motorControl.v(41[17:23])
    defparam i20224_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_843 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8587[0]), .I3(n24540), .O(n8582[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut_adj_843.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_844 (.I0(n62), .I1(n131), .I2(n8582[0]), 
            .I3(n204), .O(n8576[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut_adj_844.LUT_INIT = 16'h8778;
    SB_LUT4 i20193_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n8582[0]), 
            .O(n4_adj_3432));   // verilog/motorControl.v(41[17:23])
    defparam i20193_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20213_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n24540));   // verilog/motorControl.v(41[17:23])
    defparam i20213_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20211_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8582[0]));   // verilog/motorControl.v(41[17:23])
    defparam i20211_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_8_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3519));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3518));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3517));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3512));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3511));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3509));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3508));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_9_i24_3_lut (.I0(n34262), .I1(n103[23]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[23]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i24_3_lut (.I0(duty_23__N_3339[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[23]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i23_3_lut (.I0(n28[22]), .I1(n103[22]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[22]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i23_3_lut (.I0(duty_23__N_3339[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[22]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i22_3_lut (.I0(n28[21]), .I1(n103[21]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[21]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i22_3_lut (.I0(duty_23__N_3339[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[21]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i21_3_lut (.I0(n28[20]), .I1(n103[20]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[20]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i21_3_lut (.I0(duty_23__N_3339[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[20]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i20_3_lut (.I0(n28[19]), .I1(n103[19]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[19]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i20_3_lut (.I0(duty_23__N_3339[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[19]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i19_3_lut (.I0(n28[18]), .I1(n103[18]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[18]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i19_3_lut (.I0(duty_23__N_3339[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[18]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i18_3_lut (.I0(n28[17]), .I1(n103[17]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[17]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i18_3_lut (.I0(duty_23__N_3339[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[17]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i17_3_lut (.I0(n28[16]), .I1(n103[16]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[16]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i17_3_lut (.I0(duty_23__N_3339[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[16]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i16_3_lut (.I0(n28[15]), .I1(n103[15]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[15]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i16_3_lut (.I0(duty_23__N_3339[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[15]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i15_3_lut (.I0(n28[14]), .I1(n103[14]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[14]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i15_3_lut (.I0(duty_23__N_3339[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[14]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i14_3_lut (.I0(n28[13]), .I1(n103[13]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[13]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i14_3_lut (.I0(duty_23__N_3339[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[13]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i13_3_lut (.I0(n28[12]), .I1(n103[12]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[12]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i13_3_lut (.I0(duty_23__N_3339[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[12]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i12_3_lut (.I0(n28[11]), .I1(n103[11]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[11]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i12_3_lut (.I0(duty_23__N_3339[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[11]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i11_3_lut (.I0(n28[10]), .I1(n103[10]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[10]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i11_3_lut (.I0(duty_23__N_3339[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[10]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i10_3_lut (.I0(n28[9]), .I1(n103[9]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[9]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i10_3_lut (.I0(duty_23__N_3339[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[9]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i9_3_lut (.I0(n28[8]), .I1(n103[8]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[8]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i9_3_lut (.I0(duty_23__N_3339[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[8]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i8_3_lut (.I0(n28[7]), .I1(n103[7]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[7]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i8_3_lut (.I0(duty_23__N_3339[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[7]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i7_3_lut (.I0(n28[6]), .I1(n103[6]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[6]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i7_3_lut (.I0(duty_23__N_3339[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[6]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i6_3_lut (.I0(n28[5]), .I1(n103[5]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[5]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i6_3_lut (.I0(duty_23__N_3339[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[5]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i5_3_lut (.I0(n28[4]), .I1(n103[4]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[4]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i5_3_lut (.I0(duty_23__N_3339[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[4]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i4_3_lut (.I0(n28[3]), .I1(n103[3]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[3]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i4_3_lut (.I0(duty_23__N_3339[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[3]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i3_3_lut (.I0(n28[2]), .I1(n103[2]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[2]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i3_3_lut (.I0(duty_23__N_3339[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[2]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3507));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3506));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28754_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n34391));   // verilog/motorControl.v(43[10:25])
    defparam i28754_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_4_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_9_i2_3_lut (.I0(n28[1]), .I1(n103[1]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3339[1]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i2_3_lut (.I0(duty_23__N_3339[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3363), .I3(GND_net), .O(duty_23__N_3291[1]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3426));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i29153_2_lut_4_lut (.I0(duty[21]), .I1(n103[21]), .I2(duty[9]), 
            .I3(n103[9]), .O(n34790));
    defparam i29153_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i29163_2_lut_4_lut (.I0(duty[16]), .I1(n103[16]), .I2(duty[7]), 
            .I3(n103[7]), .O(n34800));
    defparam i29163_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i20180_2_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\Kp[1] ), .I3(\PID_CONTROLLER.err [19]), .O(n8576[0]));   // verilog/motorControl.v(41[17:23])
    defparam i20180_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3428));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29217_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n34855));
    defparam i29217_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29229_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n34867));
    defparam i29229_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_8_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3491));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3490));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i365_2_lut.LUT_INIT = 16'h8888;
    
endmodule
