// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jan 19 18:25:30 2022
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, n20154, LED_c, ENCODER0_A_N, ENCODER0_B_N, 
        ENCODER1_A_N, ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, 
        CS_c, CS_MISO_c, INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, 
        INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    
    wire n1767;
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(353[11:24])
    
    wire n59830;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(361[15:20])
    
    wire pwm_setpoint_23__N_207, n11456, n11458, n11460, n11462, n11464, 
        n11466, n11468, n11470, n11472, n11474, n11476, n11478, 
        n11480, n11482, n11484, n11486, n59913, n69708, n260, 
        n11494, n11492, n294, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n10;
    wire [23:0]pwm_setpoint_23__N_3;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    
    wire n31954, n1769, n1771, n1773;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n69765, GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, 
        GLC_N_400, dti_N_404, n31953, n31950, RX_N_2, n1765, n1763, 
        n1761, n1759, n68413, n1757, n1755;
    wire [44:0]encoder1_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
        read_N_409, n7, n1331, n68395, n24903, n20153, n62, n25, 
        n1805;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n31947;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    
    wire n59924;
    wire [5:0]color_bit_N_502;
    
    wire n59829, n41376, n41374, n59828, n59925, n41430, n24, 
        n23, n22, n21, n20, n19, n18, n17, n31945, n31942, 
        n41880, n31939, n2836, n16, n15, n14, n13;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n4, n2, n31936, n31933, n31930, n59827, n14_adj_5704, 
        n15_adj_5705, n16_adj_5706, n17_adj_5707, n18_adj_5708, n19_adj_5709, 
        n20_adj_5710, n21_adj_5711, n22_adj_5712, n23_adj_5713, n24_adj_5714, 
        n25_adj_5715, n24_adj_5716, n14992, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n27497, n4945, n4944, n4943, 
        n4923, n4922, n4924, n4925, n4926, n4927, n4928, n4929, 
        n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, 
        n4938, n4939, n4940, n4941, n4942, n20152, n3491, n2889, 
        n161, n41559, n69702, n69810, n10_adj_5717, n41590, n41584, 
        n69690, n41480, n1, n59770, n4_adj_5718, n52554, n59826, 
        n52537, n52553, n52552, n53886, n53885, n53884, n53332, 
        n53331, n53883, n53882, n53330, n53881, n53329, n53880, 
        n53879, n53328, n53878, n53327, n53326, n53877, n53876, 
        n53875, n53874, n14_adj_5719, n53873, n13_adj_5720, n53872, 
        n53871, n53870, n53869, n53868, n60434, n53867, n53866, 
        n53865, n13530, n52551, n53864, n53863, n53862, n53861, 
        n53860, n53859, n53858, n53857, n53856, n53855, n53854, 
        n53853, n53852, n53851, n53850, n52536, n53849, n53848, 
        n53847, n53846, n53845, n53844, n53843, n53842, n53841, 
        n14_adj_5721, n53840, n10_adj_5722, n70405, n53839, n53838, 
        n53837, n53836, n53835, n62592, n31927, n20159, n53834, 
        n53833, n53832, n27643, \FRAME_MATCHER.i_31__N_2509 , n53831, 
        n53830, n53829, n31908, n31897, n31893, n31890, n31887, 
        n31881, n31878, n31875, n59688, n31847, n31844, n31841, 
        n31836, n31833, n31830, n31827, n31824, n31797, n31794, 
        n31791, n31788, n31785, n31782, n31779, n31776, n31773, 
        n31770, n31767, n31755, n31745, n31742, n31739, n31736, 
        n31733, n53828, n11907, n31702, n31687, n31686, n31685, 
        n31684, n31683, n31682, n31681, n31680, n31679, n31678, 
        n31646, n31645, n31644, n31643, n31642, n31641, n31640, 
        n31639, n31638, n31637, n31636, n31635, n31634, n31633, 
        n31632, n31631, n31630, n31629, n31628, n31593, n31592, 
        n31591, n31590, n31589, n31582, n31579, n31566, n31557, 
        n53827, n53826, n53825, n61652, n53824, n26, n19_adj_5723, 
        n17_adj_5724, n16_adj_5725, n15_adj_5726, n13_adj_5727, n11, 
        n9, n8, n7_adj_5728, n6, n5, n4_adj_5729, n53823, n30, 
        n23_adj_5730, n21_adj_5731, n19_adj_5732, n17_adj_5733, n16_adj_5734, 
        n15_adj_5735, n13_adj_5736, n12, n11_adj_5737, n10_adj_5738, 
        n9_adj_5739, n8_adj_5740, n7_adj_5741, n6_adj_5742, n4_adj_5743, 
        n30_adj_5744, n23_adj_5745, n22_adj_5746, n21_adj_5747, n19_adj_5748, 
        n17_adj_5749, n16_adj_5750, n15_adj_5751, n13_adj_5752, n11_adj_5753, 
        n10_adj_5754, n9_adj_5755, n8_adj_5756, n7_adj_5757, n6_adj_5758, 
        n4_adj_5759, n17468, n53822, n59825, n31262, n59935, n59771, 
        n59824, n59823, n59919, n59822, n59920, n15_adj_5760, n59927, 
        n31257, n59922, n59821, n59946, n32706, n59820, n4_adj_5761, 
        n4_adj_5762, n32691, n4_adj_5763, n32669, n4_adj_5764, n27680, 
        n53821, n53820, n53819, n53818, n53817, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n25001, n52550, n11454, n336, n337, n338, n339, n340, 
        n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, 
        n359, n70725, n53816, n5235, n5232, n53815, n27501, n53814, 
        n3180;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, position_31__N_3836, n53813, 
        n69798, n21377, n70651, n69768, n32396, n32395, n32394, 
        n53812, n32393, n32392, n32391, n32390, n32389, n31503;
    wire [1:0]a_new_adj_5891;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5892;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5767, b_prev_adj_5768, n32388, debounce_cnt_N_3833_adj_5769, 
        n32387, n32386, n32385, n32384, position_31__N_3836_adj_5770, 
        n17_adj_5771, n13_adj_5772, n53811, n20158, n64800, n12_adj_5773, 
        n11_adj_5774, n10_adj_5775, n4_adj_5776, n3, n2_adj_5777, 
        n20151;
    wire [7:0]data_adj_5904;   // verilog/eeprom.v(23[12:16])
    wire [7:0]state_7__N_3918;
    
    wire n62593, n31500, n53810, n53809, n59921, n53808, n53807, 
        n32362, n5_adj_5778, n32360, n59062, n41527, n32356, n59819, 
        n11_adj_5779, n9_adj_5780, n32350, n53806, n53805, n6917, 
        n27667;
    wire [15:0]data_adj_5911;   // verilog/tli4970.v(27[14:18])
    
    wire n53804, n53803, n53802, n31491, n32339, n32338, n32337, 
        n32335, n32332, n32331, n32330, n32329, n32328, n32327, 
        n32326, n32325, n32324, n9_adj_5789, n8_adj_5790, n32323, 
        n32322, n32321, n32320, n32319, n32318, n32317, n32316, 
        n32315, n32314, n32313, n32312, n32311, n32308, n53801, 
        n53800, n53799, n53798, n11488, n31488, n11490, state_7__N_4319, 
        n7_adj_5791, n6_adj_5792, n5_adj_5793, n20160, n53797, n27494, 
        r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n71949;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n31482, n31481;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n31480, n53796;
    wire [2:0]r_SM_Main_adj_5927;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5928;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5929;   // verilog/uart_tx.v(34[16:27])
    
    wire n64335, n27538;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n53795, n27632, n32231, n32229, n32228, n32227, n32226, 
        n32225, n32222, n32221, n32220, n32218;
    wire [7:0]state_adj_5937;   // verilog/i2c_controller.v(33[12:17])
    
    wire n32217, n32216, n32215, n32214, n5_adj_5806, n32213, n32212, 
        n32211, n32210, n32209, n32208, n32207, n32206, enable_slow_N_4213, 
        n32203, n32202, n32201, n32200, n32199, n32197, n32196, 
        n32195, n32193, n32192, n32191, n32190;
    wire [7:0]state_7__N_4110;
    
    wire n32189, n32188, n32187, n32186, n32185, n21360, n6722;
    wire [7:0]state_7__N_4126;
    
    wire n53794, n53793, n53792, n31471, n52549, n53791, n53790, 
        n71425, n52548, n53789, n70677, n27624, n59818, n59931, 
        n59817, n31251, n59939, n53788, n29976, n59938, n53787, 
        n59937, n59816, n59815, n59941, n59814, n59940, n53786, 
        n59915, n59942, n59813, n29957, n59812, n32118, n59831, 
        n59811, n59810, n59809, n59808, n59807, n59806, n28, n53785, 
        n30_adj_5807, n31, n45, n70398, n71422, n59805, n59914, 
        n53784, n32115, n31237, n59804, n59803, n59802, n59836, 
        n59929, n59801, n53783, n8_adj_5808, n10012, n21370, n20161, 
        n152, n53782, n70835, n53781, n53780, n17462, n21376, 
        n17469, n53779, n53778, n14986, n13524, n11901, n53777, 
        n53776, n53775, n53774, n59800, n59799, n14993, n64878, 
        n13531, n11908, n52535, n21371, n17463, n71401, n1_adj_5809, 
        n53767, n59928, n53766, n53765, n53764, n52534, n144, 
        n53763, n67818, n59916, n59798, n53762, n53761, n17470, 
        n11902, n13525, n14987, n53760, n21372, n32112, n53759, 
        n71398, n20162, n53758, n59797, n14994, n13532, n11909, 
        n52547, n53757, n53756, n31269, n53755, n53754, n53753, 
        n53752, n53751, n53750, n53749, n53748, n17464, n21373, 
        n11903, n53747, n53746, n14988, n52788, n13526, n17471, 
        n14995, n69050, n52787, n53745, n20163, n13533, n52786, 
        n11910, n52785, n52784, n71395, n70900, n52783, n17465, 
        n11904, n13527, n52782, n14989, n69027, n167, n17472, 
        n52781, n27161, n52780, n52779, n14996, n52778, n13534, 
        n11911, n17466, n20164, n52777, n52776, n11905, n13528, 
        n14990, n59796, n163, n60241, n24553, n21368, n59832, 
        n59795, n14997, n13535, n11912, n59794, n53717, n59793, 
        n53716, n59792, n32108, n17467, n59791, n59947, n28963, 
        n59790, n51206, n21369, n53715, n53714, n52546, n53713, 
        n29874, n53712, n53711, n53710, n21357, n53709, n20157, 
        n20156, n20155, n53708, n53707, n53706, n20165, n53705, 
        n53704, n53703, n53702, n53701, n59789, n59945, n59788, 
        n4_adj_5810, n6_adj_5811, n8_adj_5812, n9_adj_5813, n11_adj_5814, 
        n13_adj_5815, n14_adj_5816, n15_adj_5817, n4_adj_5818, n6_adj_5819, 
        n8_adj_5820, n9_adj_5821, n29830, n71392, n29824, n29821, 
        n71389, n53700, n32101, n29817, n69433, n53699, n59787, 
        n17452, n38, n39, n40, n41, n42, n43, n44, n45_adj_5822, 
        n31463, n31462, n29799, n11914, n53698, n59786, n59944, 
        n53697, n21358, n29776, n59785, n59784, n32092, n29752, 
        n59934, n59783, n59782, n59936, n59781, n32088, n59780, 
        n32087, n59837, n59933, n59932, n68934, n69822, n55561, 
        n55706, n59779, n59910, n59778, n59909, n59777, n59908, 
        n59776, n59907, n59775, n59906, n59774, n59834, n59773, 
        n59905, n59833, n59904, n59772, n59903, n59902, n59901, 
        n59900, n59899, n59898, n59897, n59896, n59895, n59894, 
        n59893, n59892, n59891, n59890, n59889, n59888, n59887, 
        n59886, n59885, n59884, n59883, n59882, n59881, n59880, 
        n31321, n59879, n59878, n59877, n59876, n59875, n59874, 
        n59873, n59872, n59871, n59870, n59869, n59868, n59867, 
        n59866, n59865, n59864, n59863, n59862, n59861, n31159, 
        n59835, n59860, n69964, n31299, n59859, n59858, n59857, 
        n59856, n31294, n59855, n59854, n59853, n59852, n59851, 
        n59850, n59849, n59848, n55737, n60431, n59847, n31284, 
        n59846, n59845, n59844, n59843, n31109, n59842, n59841, 
        n31277, n59840, n59839, n59838, n6_adj_5823, n30452, n30449, 
        n30447, n60038, n60042, n60044, n30423, n60039, n30416, 
        n30414, n30382, n30865, n30370, n30368, n30366, n30362, 
        n28303, n28330, n59917, n20166, n59911, n59912, n68918, 
        n27629, n21359, n59930, n20167, n52533, n9949, n9947, 
        n13514, n11891, n14976, n20168, n17454, n13515, n14977, 
        n11892, n17453, n11893, n13516, n14978, n11894, n13517, 
        n52545, n14979, n24877, n17455, n14980, n17456, n54181, 
        n32083, n32078, n32074, n32066, n32065, n59136, n11896, 
        n13519, n14981, n17457, n29728, n11895, n13518, n71386, 
        n27672, n14982, n17458, n59138, n11897, n52544, n13520, 
        n31455, n52543, n32021, n32020, n59140, n17459, n11898, 
        n14983, n13521, n31452, n31449, n31446, n59142, n11899, 
        n13522, n14984, n21361, n21374, n17460, n61872, n59144, 
        n31996, n59146, n31990, n59148, n59150, n31977, n31974, 
        n31971, n21375, n17461, n52532, n31443, n31440, n31436, 
        n31968, n31965, n11900, n13523, n14985, n31961, n59943, 
        n52542, n20169, n21362, n11913, n13536, n21363, n59923, 
        n21364, n21365, n21366, n53618, n53617, n53616, n53615, 
        n21367, n52541, n53614, n68829, n53613, n53612, n53611, 
        n53610, n53609, n53608, n53607, n53606, n53605, n14991, 
        n53604, n53603, n53602, n53601, n53600, n10_adj_5824, n53599, 
        n52540, n64457, n11452, n64702, n64890, n62898, n54982, 
        n64614, n13508, n11885, n52706, n52705, n52704, n14971, 
        n52703, n13509, n27099, n11886, n62445, n13529, n52702, 
        n14972, n13510, n52701, n52700, n11887, n52699, n17449, 
        n52698, n52539, n14973, n13511, n11888, n52697, n55814, 
        n17450, n6_adj_5825, n52696, n52695, n52694, n14974, n71638, 
        n13512, n59660, n64459, n11889, n52693, n71632, n52692, 
        n11906, n71626, n17451, n28021, n71620, n14975, n27661, 
        n54699, n13513, n71614, n11890, n71608, n64693, n54679, 
        n52691, n52690, n52689, n52688, n52531, n52687, n52686, 
        n68812, n23767, n54659, n52685, n52684, n68795, n59926, 
        n20170, n20171, n20172, n52538, n71602, n52652, n62537, 
        n52651, n52650, n52649, n52648, n52647, n52560, n52646, 
        n52645, n52644, n52643, n52559, n52642, n52641, n30156, 
        n64701, n54578, n52640, n8_adj_5826, n7_adj_5827, n52639, 
        n52558, n70414, n52638, n52637, n64692, n52636, n52530, 
        n52635, n52634, n71596, n62228, n52633, n52557, n52632, 
        n52631, n52630, n52556, n59918, n52555, n70290, n12_adj_5828, 
        n71590, n70300, n70749, n70899, n68632, n4_adj_5829, n68610, 
        n69970, n6_adj_5830, n71584, n68582, n64469, n15_adj_5831, 
        n71578, n63595, n14_adj_5832, n17_adj_5833, n25_adj_5834, 
        n58068, n24_adj_5835, n63577, n63571, n70390, n63565, n4_adj_5836, 
        n70391, n15_adj_5837, n14_adj_5838, n63559, n58154, n63557, 
        n63551, n71572, n71705, n63545, n63537, n63531, n63525, 
        n6_adj_5839, n71566, n63519, n63513, n63507, n60846, n63501, 
        n60834, n63495, n60832, n71560, n67768, n63489, n63483, 
        n63477, n63471, n67759, n63465, n60355, n61989, n71554, 
        n25_adj_5840, n24_adj_5841, n23_adj_5842, n63459, n67750, 
        n63453, n60391, n63447, n67748, n63441, n67737, n67734, 
        n63435, n60741, n29, n27, n60669, n23_adj_5843, n62047, 
        n64287, n70724, n64615, n71341, n64891, n71548, n64880, 
        n64879, n67643, n70842, n70836, n71542, n58944, n71536, 
        n70736, n64291, n58986, n71530, n7_adj_5844, n64283, n22_adj_5845, 
        n71338, n70658, n71524, n71521, n70657, n59110, n59114, 
        n60470, n59122, n59126, n63199, n63193, n6_adj_5846, n63187, 
        n8_adj_5847, n63181, n63177, n63175, n67594, n37, n35, 
        n62670, n34, n70622, n32, n31_adj_5848, n25_adj_5849, n6_adj_5850, 
        n70565, n67837, n59686, n4_adj_5851, n67830, n70404, n63043, 
        n60254, n63019, n60592, n70653, n70088, n70403, n70417, 
        n64806, n64804, n64803, n70301, n7_adj_5852;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13), .I3(n52695), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n29728), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n52695), .I0(encoder0_position_scaled[12]), 
            .I1(n13), .CO(n52696));
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.n29957(n29957), .bit_ctr({bit_ctr[4], 
            Open_0, Open_1, bit_ctr[1], Open_2}), .clk16MHz(clk16MHz), 
            .GND_net(GND_net), .state({state}), .\neopxl_color[5] (neopxl_color[5]), 
            .\neopxl_color[4] (neopxl_color[4]), .\color_bit_N_502[1] (color_bit_N_502[1]), 
            .n31755(n31755), .VCC_net(VCC_net), .n58944(n58944), .n31687(n31687), 
            .t0({t0}), .n31686(n31686), .n31685(n31685), .timer({timer}), 
            .n31684(n31684), .n31683(n31683), .n31682(n31682), .\bit_ctr[3] (bit_ctr[3]), 
            .n31681(n31681), .n31680(n31680), .n31679(n31679), .n31678(n31678), 
            .\bit_ctr[0] (bit_ctr[0]), .NEOPXL_c(NEOPXL_c), .n31481(n31481), 
            .n27099(n27099), .LED_c(LED_c), .n41559(n41559), .n54699(n54699), 
            .\color_bit_N_502[2] (color_bit_N_502[2]), .n3180(n3180), .\neopxl_color[14] (neopxl_color[14]), 
            .\neopxl_color[15] (neopxl_color[15]), .\neopxl_color[12] (neopxl_color[12]), 
            .\neopxl_color[13] (neopxl_color[13]), .n71341(n71341), .n54679(n54679), 
            .n71425(n71425), .n71395(n71395), .\neopxl_color[6] (neopxl_color[6]), 
            .\neopxl_color[7] (neopxl_color[7])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 mux_245_i10_4_lut (.I0(displacement[9]), .I1(encoder0_position_scaled[9]), 
            .I2(n54181), .I3(n51206), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n52694), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n52694), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n52695));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15), .I3(n52693), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n52693), .I0(encoder0_position_scaled[10]), 
            .I1(n15), .CO(n52694));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16), .I3(n52692), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52112 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[0]), .O(n71398));
    defparam byte_transmit_counter_1__bdd_4_lut_52112.LUT_INIT = 16'he4aa;
    SB_LUT4 n71398_bdd_4_lut (.I0(n71398), .I1(\data_out_frame[26] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[0]), 
            .O(n71401));
    defparam n71398_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n71392_bdd_4_lut (.I0(n71392), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n71395));
    defparam n71392_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n60241));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut (.I0(n144), .I1(n10_adj_5717), .I2(reset), .I3(GND_net), 
            .O(n30423));
    defparam i2_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[6] [0]), .I1(n30382), .I2(n30423), 
            .I3(rx_data[0]), .O(n59122));
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i48560_3_lut_4_lut (.I0(r_Clock_Count_adj_5928[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5928[2]), .O(n67830));   // verilog/uart_tx.v(117[17:57])
    defparam i48560_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1183_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5928[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5811));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n52692), .I0(encoder0_position_scaled[9]), 
            .I1(n16), .CO(n52693));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17), .I3(n52691), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n52691), .I0(encoder0_position_scaled[8]), 
            .I1(n17), .CO(n52692));
    SB_LUT4 add_5391_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(encoder1_position[21]), 
            .I3(n53618), .O(n21357)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13683_3_lut (.I0(current[11]), .I1(data_adj_5911[11]), .I2(n29799), 
            .I3(GND_net), .O(n31628));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18), .I3(n52690), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n52690), .I0(encoder0_position_scaled[7]), 
            .I1(n18), .CO(n52691));
    SB_LUT4 i13684_3_lut (.I0(current[10]), .I1(data_adj_5911[10]), .I2(n29799), 
            .I3(GND_net), .O(n31629));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13685_3_lut (.I0(current[9]), .I1(data_adj_5911[9]), .I2(n29799), 
            .I3(GND_net), .O(n31630));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13686_3_lut (.I0(current[8]), .I1(data_adj_5911[8]), .I2(n29799), 
            .I3(GND_net), .O(n31631));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13687_3_lut (.I0(current[7]), .I1(data_adj_5911[7]), .I2(n29799), 
            .I3(GND_net), .O(n31632));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13688_3_lut (.I0(current[6]), .I1(data_adj_5911[6]), .I2(n29799), 
            .I3(GND_net), .O(n31633));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[16] [4]), .I1(n28330), .I2(n54659), 
            .I3(n4_adj_5836), .O(n27161));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\data_out_frame[23] [7]), .I1(n60741), .I2(\data_out_frame[24] [7]), 
            .I3(n60470), .O(n34));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n25_adj_5840), .I1(n60391), .I2(n23_adj_5842), 
            .I3(n24_adj_5841), .O(n25_adj_5849));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13689_3_lut (.I0(current[5]), .I1(data_adj_5911[5]), .I2(n29799), 
            .I3(GND_net), .O(n31634));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1789 (.I0(n60669), .I1(\data_out_frame[24] [2]), 
            .I2(n60431), .I3(\data_out_frame[25] [1]), .O(n32));
    defparam i12_4_lut_adj_1789.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_out_frame[25] [4]), .I1(n60434), .I2(\data_out_frame[23] [5]), 
            .I3(n61872), .O(n31_adj_5848));
    defparam i11_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[23] [1]), 
            .I2(n55706), .I3(\data_out_frame[24] [3]), .O(n35));
    defparam i15_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut (.I0(n25_adj_5849), .I1(n34), .I2(\data_out_frame[23] [4]), 
            .I3(n60592), .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13690_3_lut (.I0(current[4]), .I1(data_adj_5911[4]), .I2(n29799), 
            .I3(GND_net), .O(n31635));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n52689), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31_adj_5848), .I3(n32), 
            .O(n55737));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13691_3_lut (.I0(current[3]), .I1(data_adj_5911[3]), .I2(n29799), 
            .I3(GND_net), .O(n31636));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5391_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(encoder1_position[20]), 
            .I3(n53617), .O(n21358)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13692_3_lut (.I0(current[2]), .I1(data_adj_5911[2]), .I2(n29799), 
            .I3(GND_net), .O(n31637));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13693_3_lut (.I0(current[1]), .I1(data_adj_5911[1]), .I2(n29799), 
            .I3(GND_net), .O(n31638));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13693_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5391_21 (.CI(n53617), .I0(encoder1_position[19]), .I1(encoder1_position[20]), 
            .CO(n53618));
    SB_LUT4 add_5391_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(encoder1_position[19]), 
            .I3(n53616), .O(n21359)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n52689), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n52690));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n52688), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n52688), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n52689));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n52687), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n52687), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n52688));
    SB_CARRY add_5391_20 (.CI(n53616), .I0(encoder1_position[18]), .I1(encoder1_position[19]), 
            .CO(n53617));
    SB_LUT4 add_5391_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(encoder1_position[18]), 
            .I3(n53615), .O(n21360)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(n30), .I1(current_limit[15]), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5745));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13694_3_lut (.I0(baudrate[31]), .I1(data_adj_5904[7]), .I2(n29874), 
            .I3(GND_net), .O(n31639));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5757));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5755));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52092 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n71386));
    defparam byte_transmit_counter_0__bdd_4_lut_52092.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5748));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5747));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n52532), .O(n1248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5753));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5752));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13695_3_lut (.I0(baudrate[30]), .I1(data_adj_5904[6]), .I2(n29874), 
            .I3(GND_net), .O(n31640));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n52686), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n71386_bdd_4_lut (.I0(n71386), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n71389));
    defparam n71386_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5751));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n52686), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n52687));
    SB_LUT4 LessThan_14_i23_2_lut (.I0(current[11]), .I1(current_limit[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5730));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5733));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5732));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13696_3_lut (.I0(baudrate[29]), .I1(data_adj_5904[5]), .I2(n29874), 
            .I3(GND_net), .O(n31641));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13696_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5391_19 (.CI(n53615), .I0(encoder1_position[17]), .I1(encoder1_position[18]), 
            .CO(n53616));
    SB_LUT4 LessThan_14_i21_2_lut (.I0(current[10]), .I1(current_limit[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5731));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5737));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5736));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5735));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5391_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(encoder1_position[17]), 
            .I3(n53614), .O(n21361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n52685), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5391_18 (.CI(n53614), .I0(encoder1_position[16]), .I1(encoder1_position[17]), 
            .CO(n53615));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n52685), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n52686));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n52684), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5391_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(encoder1_position[16]), 
            .I3(n53613), .O(n21362)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5741));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5739));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n52684), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n52685));
    SB_LUT4 i50163_4_lut (.I0(n9_adj_5739), .I1(n7_adj_5741), .I2(current_limit[2]), 
            .I3(current[2]), .O(n69433));
    defparam i50163_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i13697_3_lut (.I0(baudrate[28]), .I1(data_adj_5904[4]), .I2(n29874), 
            .I3(GND_net), .O(n31642));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13697_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5391_17 (.CI(n53613), .I0(encoder1_position[15]), .I1(encoder1_position[16]), 
            .CO(n53614));
    SB_LUT4 add_5391_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(encoder1_position[15]), 
            .I3(n53612), .O(n21363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50700_4_lut (.I0(n15_adj_5735), .I1(n13_adj_5736), .I2(n11_adj_5737), 
            .I3(n69433), .O(n69970));
    defparam i50700_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50694_4_lut (.I0(n21_adj_5731), .I1(n19_adj_5732), .I2(n17_adj_5733), 
            .I3(n69970), .O(n69964));
    defparam i50694_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5743));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 LessThan_14_i12_3_lut (.I0(n10_adj_5738), .I1(current_limit[7]), 
            .I2(n15_adj_5735), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25), .CO(n52684));
    SB_LUT4 n9949_bdd_4_lut (.I0(n9949), .I1(current[15]), .I2(duty[22]), 
            .I3(n9947), .O(n71638));
    defparam n9949_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_CARRY add_5391_16 (.CI(n53612), .I0(encoder1_position[14]), .I1(encoder1_position[15]), 
            .CO(n53613));
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i13698_3_lut (.I0(baudrate[27]), .I1(data_adj_5904[3]), .I2(n29874), 
            .I3(GND_net), .O(n31643));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13822_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n60042), 
            .I3(GND_net), .O(n31767));   // verilog/coms.v(130[12] 305[6])
    defparam i13822_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5740), .I1(current_limit[9]), 
            .I2(n19_adj_5732), .I3(GND_net), .O(n16_adj_5734));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i51387_4_lut (.I0(n16_adj_5734), .I1(n6_adj_5742), .I2(n19_adj_5732), 
            .I3(n68395), .O(n70657));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51387_4_lut.LUT_INIT = 16'haaac;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i51388_3_lut (.I0(n70657), .I1(current_limit[10]), .I2(n21_adj_5731), 
            .I3(GND_net), .O(n70658));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51128_3_lut (.I0(n70658), .I1(current_limit[11]), .I2(n23_adj_5730), 
            .I3(GND_net), .O(n70398));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5391_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(encoder1_position[14]), 
            .I3(n53611), .O(n21364)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51295_4_lut (.I0(current[15]), .I1(n23_adj_5730), .I2(current_limit[12]), 
            .I3(n69964), .O(n70565));
    defparam i51295_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51147_4_lut (.I0(n12), .I1(n4_adj_5743), .I2(n15_adj_5735), 
            .I3(n68413), .O(n70417));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51147_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50495_3_lut (.I0(n70398), .I1(current_limit[12]), .I2(current[15]), 
            .I3(GND_net), .O(n69765));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50495_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51381_3_lut (.I0(n69765), .I1(n70417), .I2(n70565), .I3(GND_net), 
            .O(n70651));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51381_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5391_15 (.CI(n53611), .I0(encoder1_position[13]), .I1(encoder1_position[14]), 
            .CO(n53612));
    SB_LUT4 add_5391_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(encoder1_position[13]), 
            .I3(n53610), .O(n21365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51156_4_lut (.I0(n70651), .I1(current_limit[14]), .I2(current[15]), 
            .I3(current_limit[13]), .O(n30));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51156_4_lut.LUT_INIT = 16'h8f0e;
    SB_CARRY add_5391_14 (.CI(n53610), .I0(encoder1_position[12]), .I1(encoder1_position[13]), 
            .CO(n53611));
    SB_LUT4 n71638_bdd_4_lut (.I0(n71638), .I1(duty[19]), .I2(n4926), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[19]));
    defparam n71638_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13699_3_lut (.I0(baudrate[26]), .I1(data_adj_5904[2]), .I2(n29874), 
            .I3(GND_net), .O(n31644));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5391_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(encoder1_position[12]), 
            .I3(n53609), .O(n21366)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19282_3_lut (.I0(n30), .I1(current_limit[15]), .I2(current[15]), 
            .I3(GND_net), .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i19282_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i13825_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n60042), 
            .I3(GND_net), .O(n31770));   // verilog/coms.v(130[12] 305[6])
    defparam i13825_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13700_3_lut (.I0(baudrate[25]), .I1(data_adj_5904[1]), .I2(n29874), 
            .I3(GND_net), .O(n31645));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13700_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5391_13 (.CI(n53609), .I0(encoder1_position[11]), .I1(encoder1_position[12]), 
            .CO(n53610));
    SB_LUT4 add_5391_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(encoder1_position[11]), 
            .I3(n53608), .O(n21367)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13828_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n60042), 
            .I3(GND_net), .O(n31773));   // verilog/coms.v(130[12] 305[6])
    defparam i13828_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5391_12 (.CI(n53608), .I0(encoder1_position[10]), .I1(encoder1_position[11]), 
            .CO(n53609));
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5723));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5391_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(encoder1_position[10]), 
            .I3(n53607), .O(n21368)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13831_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n60039), .I3(GND_net), .O(n31776));   // verilog/coms.v(130[12] 305[6])
    defparam i13831_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5391_11 (.CI(n53607), .I0(encoder1_position[9]), .I1(encoder1_position[10]), 
            .CO(n53608));
    SB_LUT4 add_5391_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(encoder1_position[9]), 
            .I3(n53606), .O(n21369)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5391_10 (.CI(n53606), .I0(encoder1_position[8]), .I1(encoder1_position[9]), 
            .CO(n53607));
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5728));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5726));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5724));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13834_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n60039), .I3(GND_net), .O(n31779));   // verilog/coms.v(130[12] 305[6])
    defparam i13834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5727));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n67594), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5729));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51030_3_lut (.I0(n4_adj_5729), .I1(n305), .I2(n11), .I3(GND_net), 
            .O(n70300));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13701_3_lut (.I0(baudrate[24]), .I1(data_adj_5904[0]), .I2(n29874), 
            .I3(GND_net), .O(n31646));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51031_3_lut (.I0(n70300), .I1(n304), .I2(n13_adj_5727), .I3(GND_net), 
            .O(n70301));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13837_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n60039), .I3(GND_net), .O(n31782));   // verilog/coms.v(130[12] 305[6])
    defparam i13837_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17_adj_5724), 
            .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7_adj_5728), 
            .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13840_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n60039), .I3(GND_net), .O(n31785));   // verilog/coms.v(130[12] 305[6])
    defparam i13840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8), .I1(n301), .I2(n19_adj_5723), 
            .I3(GND_net), .O(n16_adj_5725));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13843_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n60039), .I3(GND_net), .O(n31788));   // verilog/coms.v(130[12] 305[6])
    defparam i13843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_5391_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(encoder1_position[8]), 
            .I3(n53605), .O(n21370)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13846_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n60039), .I3(GND_net), .O(n31791));   // verilog/coms.v(130[12] 305[6])
    defparam i13846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13849_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n60039), .I3(GND_net), .O(n31794));   // verilog/coms.v(130[12] 305[6])
    defparam i13849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49362_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5728), .I3(n5), 
            .O(n68632));
    defparam i49362_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49340_4_lut (.I0(n17_adj_5724), .I1(n15_adj_5726), .I2(n13_adj_5727), 
            .I3(n68632), .O(n68610));
    defparam i49340_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13852_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n60039), .I3(GND_net), .O(n31797));   // verilog/coms.v(130[12] 305[6])
    defparam i13852_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i51383_4_lut (.I0(n16_adj_5725), .I1(n6), .I2(n19_adj_5723), 
            .I3(n68582), .O(n70653));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51383_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49648_3_lut (.I0(n70301), .I1(n303), .I2(n15_adj_5726), .I3(GND_net), 
            .O(n68918));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i49648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51565_4_lut (.I0(n68918), .I1(n70653), .I2(n19_adj_5723), 
            .I3(n68610), .O(n70835));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51565_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51566_3_lut (.I0(n70835), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n70836));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51566_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51479_3_lut (.I0(n70836), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n70749));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51479_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n9949_bdd_4_lut_52285 (.I0(n9949), .I1(current[15]), .I2(duty[21]), 
            .I3(n9947), .O(n71632));
    defparam n9949_bdd_4_lut_52285.LUT_INIT = 16'he4aa;
    SB_LUT4 i45032_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n294), .I3(GND_net), 
            .O(n64287));
    defparam i45032_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i26_3_lut (.I0(n70749), .I1(n298), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45036_3_lut (.I0(duty[13]), .I1(duty[21]), .I2(n294), .I3(GND_net), 
            .O(n64291));
    defparam i45036_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i45198_4_lut (.I0(duty[15]), .I1(n64287), .I2(duty[20]), .I3(n294), 
            .O(n64459));
    defparam i45198_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i45028_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n64283));
    defparam i45028_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i10_4_lut (.I0(n294), .I1(n64459), .I2(n64291), .I3(n26), 
            .O(n22_adj_5845));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i45196_4_lut (.I0(duty[19]), .I1(n64283), .I2(duty[16]), .I3(n294), 
            .O(n64457));
    defparam i45196_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i13991_3_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(n62228), .I3(GND_net), .O(n31936));   // verilog/coms.v(130[12] 305[6])
    defparam i13991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49757_3_lut (.I0(n15_adj_5751), .I1(n13_adj_5752), .I2(n11_adj_5753), 
            .I3(GND_net), .O(n69027));
    defparam i49757_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_5391_9 (.CI(n53605), .I0(encoder1_position[7]), .I1(encoder1_position[8]), 
            .CO(n53606));
    SB_LUT4 add_5391_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(encoder1_position[7]), 
            .I3(n53604), .O(n21371)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5391_8 (.CI(n53604), .I0(encoder1_position[6]), .I1(encoder1_position[7]), 
            .CO(n53605));
    SB_LUT4 i50432_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n69027), .O(n69702));
    defparam i50432_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i48567_4_lut (.I0(n21_adj_5747), .I1(n19_adj_5748), .I2(n17_adj_5749), 
            .I3(n9_adj_5755), .O(n67837));
    defparam i48567_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n71632_bdd_4_lut (.I0(n71632), .I1(duty[18]), .I2(n4927), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[18]));
    defparam n71632_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49780_4_lut (.I0(n9_adj_5755), .I1(n7_adj_5757), .I2(current[2]), 
            .I3(duty[2]), .O(n69050));
    defparam i49780_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 add_5391_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(encoder1_position[6]), 
            .I3(n53603), .O(n21372)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50540_4_lut (.I0(n15_adj_5751), .I1(n13_adj_5752), .I2(n11_adj_5753), 
            .I3(n69050), .O(n69810));
    defparam i50540_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50528_4_lut (.I0(n21_adj_5747), .I1(n19_adj_5748), .I2(n17_adj_5749), 
            .I3(n69810), .O(n69798));
    defparam i50528_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51135_4_lut (.I0(current[15]), .I1(n23_adj_5745), .I2(duty[12]), 
            .I3(n69798), .O(n70405));
    defparam i51135_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i49542_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n70405), .O(n68812));
    defparam i49542_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5759));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i51020_3_lut (.I0(n4_adj_5759), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n70290));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51020_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n9949_bdd_4_lut_52280 (.I0(n9949), .I1(current[15]), .I2(duty[20]), 
            .I3(n9947), .O(n71626));
    defparam n9949_bdd_4_lut_52280.LUT_INIT = 16'he4aa;
    SB_LUT4 i50420_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5751), .O(n69690));
    defparam i50420_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5744));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i49525_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n69702), .O(n68795));
    defparam i49525_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_11_i35_rep_238_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n71949));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_238_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51466_3_lut (.I0(n30_adj_5744), .I1(n10_adj_5754), .I2(n69690), 
            .I3(GND_net), .O(n70736));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49664_4_lut (.I0(n70290), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n68934));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i49664_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 n71626_bdd_4_lut (.I0(n71626), .I1(duty[17]), .I2(n4928), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[17]));
    defparam n71626_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51133_3_lut (.I0(n6_adj_5758), .I1(duty[10]), .I2(n21_adj_5747), 
            .I3(GND_net), .O(n70403));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51134_3_lut (.I0(n70403), .I1(duty[11]), .I2(n23_adj_5745), 
            .I3(GND_net), .O(n70404));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50438_4_lut (.I0(current[15]), .I1(n23_adj_5745), .I2(duty[12]), 
            .I3(n67837), .O(n69708));
    defparam i50438_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5756), .I1(duty[9]), .I2(n19_adj_5748), 
            .I3(GND_net), .O(n16_adj_5750));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50848_3_lut (.I0(n70404), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n22_adj_5746));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50848_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50818_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n68812), .O(n70088));
    defparam i50818_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i13994_3_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(n62228), .I3(GND_net), .O(n31939));   // verilog/coms.v(130[12] 305[6])
    defparam i13994_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_14 (.CI(n52541), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n52542));
    SB_LUT4 i51572_4_lut (.I0(n68934), .I1(n70736), .I2(n71949), .I3(n68795), 
            .O(n70842));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51572_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50498_3_lut (.I0(n22_adj_5746), .I1(n16_adj_5750), .I2(n69708), 
            .I3(GND_net), .O(n69768));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51629_4_lut (.I0(n69768), .I1(n70842), .I2(n71949), .I3(n70088), 
            .O(n70899));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51629_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51630_3_lut (.I0(n70899), .I1(duty[18]), .I2(current[15]), 
            .I3(GND_net), .O(n70900));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51630_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5391_7 (.CI(n53603), .I0(encoder1_position[5]), .I1(encoder1_position[6]), 
            .CO(n53604));
    SB_LUT4 i51144_4_lut (.I0(n70900), .I1(duty[20]), .I2(current[15]), 
            .I3(duty[19]), .O(n70414));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51144_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 add_5391_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(encoder1_position[5]), 
            .I3(n53602), .O(n21373)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1790 (.I0(n70414), .I1(n7), .I2(duty[21]), .I3(current[15]), 
            .O(n6_adj_5823));
    defparam i2_4_lut_adj_1790.LUT_INIT = 16'hecfe;
    SB_LUT4 i7_4_lut (.I0(duty[22]), .I1(duty[23]), .I2(n6_adj_5823), 
            .I3(current[15]), .O(n9949));
    defparam i7_4_lut.LUT_INIT = 16'h3332;
    SB_CARRY add_5391_6 (.CI(n53602), .I0(encoder1_position[4]), .I1(encoder1_position[5]), 
            .CO(n53603));
    SB_LUT4 add_5391_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[4]), 
            .I3(n53601), .O(n21374)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9949_bdd_4_lut_52275 (.I0(n9949), .I1(current[15]), .I2(duty[19]), 
            .I3(n9947), .O(n71620));
    defparam n9949_bdd_4_lut_52275.LUT_INIT = 16'he4aa;
    SB_CARRY add_5391_5 (.CI(n53601), .I0(encoder1_position[3]), .I1(encoder1_position[4]), 
            .CO(n53602));
    SB_LUT4 add_5391_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[3]), 
            .I3(n53600), .O(n21375)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13879_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n60038), .I3(GND_net), .O(n31824));   // verilog/coms.v(130[12] 305[6])
    defparam i13879_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_5391_4 (.CI(n53600), .I0(encoder1_position[2]), .I1(encoder1_position[3]), 
            .CO(n53601));
    SB_LUT4 i13882_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n60038), .I3(GND_net), .O(n31827));   // verilog/coms.v(130[12] 305[6])
    defparam i13882_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_5391_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n53599), .O(n21376)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13885_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n60038), .I3(GND_net), .O(n31830));   // verilog/coms.v(130[12] 305[6])
    defparam i13885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71620_bdd_4_lut (.I0(n71620), .I1(duty[16]), .I2(n4929), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[16]));
    defparam n71620_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_5391_3 (.CI(n53599), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n53600));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5391_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n21377)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5391_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5391_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n53599));
    SB_LUT4 n9949_bdd_4_lut_52270 (.I0(n9949), .I1(current[15]), .I2(duty[18]), 
            .I3(n9947), .O(n71614));
    defparam n9949_bdd_4_lut_52270.LUT_INIT = 16'he4aa;
    SB_LUT4 n71614_bdd_4_lut (.I0(n71614), .I1(duty[15]), .I2(n4930), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[15]));
    defparam n71614_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52265 (.I0(n9949), .I1(current[15]), .I2(duty[17]), 
            .I3(n9947), .O(n71608));
    defparam n9949_bdd_4_lut_52265.LUT_INIT = 16'he4aa;
    SB_LUT4 n71608_bdd_4_lut (.I0(n71608), .I1(duty[14]), .I2(n4931), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[14]));
    defparam n71608_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52260 (.I0(n9949), .I1(current[15]), .I2(duty[16]), 
            .I3(n9947), .O(n71602));
    defparam n9949_bdd_4_lut_52260.LUT_INIT = 16'he4aa;
    SB_LUT4 n71602_bdd_4_lut (.I0(n71602), .I1(duty[13]), .I2(n4932), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[13]));
    defparam n71602_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52255 (.I0(n9949), .I1(current[15]), .I2(duty[15]), 
            .I3(n9947), .O(n71596));
    defparam n9949_bdd_4_lut_52255.LUT_INIT = 16'he4aa;
    SB_LUT4 n71596_bdd_4_lut (.I0(n71596), .I1(duty[12]), .I2(n4933), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[12]));
    defparam n71596_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52250 (.I0(n9949), .I1(current[11]), .I2(duty[14]), 
            .I3(n9947), .O(n71590));
    defparam n9949_bdd_4_lut_52250.LUT_INIT = 16'he4aa;
    SB_LUT4 n71590_bdd_4_lut (.I0(n71590), .I1(duty[11]), .I2(n4934), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[11]));
    defparam n71590_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52245 (.I0(n9949), .I1(current[10]), .I2(duty[13]), 
            .I3(n9947), .O(n71584));
    defparam n9949_bdd_4_lut_52245.LUT_INIT = 16'he4aa;
    SB_LUT4 n71584_bdd_4_lut (.I0(n71584), .I1(duty[10]), .I2(n4935), 
            .I3(n9947), .O(pwm_setpoint_23__N_3[10]));
    defparam n71584_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52240 (.I0(n9949), .I1(current[9]), .I2(duty[12]), 
            .I3(n9947), .O(n71578));
    defparam n9949_bdd_4_lut_52240.LUT_INIT = 16'he4aa;
    SB_LUT4 n71578_bdd_4_lut (.I0(n71578), .I1(duty[9]), .I2(n4936), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n71578_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52235 (.I0(n9949), .I1(current[8]), .I2(duty[11]), 
            .I3(n9947), .O(n71572));
    defparam n9949_bdd_4_lut_52235.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1791 (.I0(\data_out_frame[24] [2]), .I1(n62047), 
            .I2(GND_net), .I3(GND_net), .O(n60254));
    defparam i1_2_lut_adj_1791.LUT_INIT = 16'h9999;
    SB_LUT4 i13997_3_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(n62228), .I3(GND_net), .O(n31942));   // verilog/coms.v(130[12] 305[6])
    defparam i13997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13888_3_lut (.I0(\data_in_frame[12] [3]), .I1(rx_data[3]), 
            .I2(n60038), .I3(GND_net), .O(n31833));   // verilog/coms.v(130[12] 305[6])
    defparam i13888_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n71572_bdd_4_lut (.I0(n71572), .I1(duty[8]), .I2(n4937), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n71572_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13891_3_lut (.I0(\data_in_frame[12] [4]), .I1(rx_data[4]), 
            .I2(n60038), .I3(GND_net), .O(n31836));   // verilog/coms.v(130[12] 305[6])
    defparam i13891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9949_bdd_4_lut_52230 (.I0(n9949), .I1(current[7]), .I2(duty[10]), 
            .I3(n9947), .O(n71566));
    defparam n9949_bdd_4_lut_52230.LUT_INIT = 16'he4aa;
    SB_LUT4 i13896_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n60038), .I3(GND_net), .O(n31841));   // verilog/coms.v(130[12] 305[6])
    defparam i13896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71566_bdd_4_lut (.I0(n71566), .I1(duty[7]), .I2(n4938), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n71566_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_245_i4_4_lut (.I0(displacement[3]), .I1(encoder0_position_scaled[3]), 
            .I2(n54181), .I3(n51206), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i13899_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n60038), .I3(GND_net), .O(n31844));   // verilog/coms.v(130[12] 305[6])
    defparam i13899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i5_4_lut (.I0(displacement[4]), .I1(encoder0_position_scaled[4]), 
            .I2(n54181), .I3(n51206), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 n9949_bdd_4_lut_52225 (.I0(n9949), .I1(current[6]), .I2(duty[9]), 
            .I3(n9947), .O(n71560));
    defparam n9949_bdd_4_lut_52225.LUT_INIT = 16'he4aa;
    SB_LUT4 n71560_bdd_4_lut (.I0(n71560), .I1(duty[6]), .I2(n4939), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n71560_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52220 (.I0(n9949), .I1(current[5]), .I2(duty[8]), 
            .I3(n9947), .O(n71554));
    defparam n9949_bdd_4_lut_52220.LUT_INIT = 16'he4aa;
    SB_LUT4 n71554_bdd_4_lut (.I0(n71554), .I1(duty[5]), .I2(n4940), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n71554_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52215 (.I0(n9949), .I1(current[4]), .I2(duty[7]), 
            .I3(n9947), .O(n71548));
    defparam n9949_bdd_4_lut_52215.LUT_INIT = 16'he4aa;
    SB_LUT4 n71548_bdd_4_lut (.I0(n71548), .I1(duty[4]), .I2(n4941), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n71548_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5833));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 n9949_bdd_4_lut_52210 (.I0(n9949), .I1(current[3]), .I2(duty[6]), 
            .I3(n9947), .O(n71542));
    defparam n9949_bdd_4_lut_52210.LUT_INIT = 16'he4aa;
    SB_LUT4 i13733_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3180), .I3(GND_net), 
            .O(n31678));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n52540), .O(n1240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71542_bdd_4_lut (.I0(n71542), .I1(duty[3]), .I2(n4942), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n71542_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13734_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3180), .I3(GND_net), 
            .O(n31679));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9949_bdd_4_lut_52205 (.I0(n9949), .I1(current[2]), .I2(duty[5]), 
            .I3(n9947), .O(n71536));
    defparam n9949_bdd_4_lut_52205.LUT_INIT = 16'he4aa;
    SB_DFFESR dti_counter_2039__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n29976), 
            .D(n45_adj_5822), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_151_5 (.CI(n52532), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n52533));
    SB_LUT4 n71536_bdd_4_lut (.I0(n71536), .I1(duty[2]), .I2(n4943), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n71536_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13735_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3180), .I3(GND_net), 
            .O(n31680));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_52107 (.I0(color_bit_N_502[1]), .I1(n64692), 
            .I2(n64693), .I3(color_bit_N_502[2]), .O(n71338));
    defparam color_bit_N_502_1__bdd_4_lut_52107.LUT_INIT = 16'he4aa;
    SB_CARRY add_151_13 (.CI(n52540), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n52541));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n52560), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71338_bdd_4_lut (.I0(n71338), .I1(n64702), .I2(n64701), .I3(color_bit_N_502[2]), 
            .O(n71341));
    defparam n71338_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9949_bdd_4_lut_52200 (.I0(n9949), .I1(current[1]), .I2(duty[4]), 
            .I3(n9947), .O(n71530));
    defparam n9949_bdd_4_lut_52200.LUT_INIT = 16'he4aa;
    SB_LUT4 i13736_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3180), .I3(GND_net), 
            .O(n31681));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13736_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n52559), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 n71530_bdd_4_lut (.I0(n71530), .I1(duty[1]), .I2(n4944), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n71530_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_151_32 (.CI(n52559), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n52560));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n52558), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n52652), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_24_lut (.I0(GND_net), .I1(GND_net), .I2(n11452), 
            .I3(n52651), .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dti_counter_2039__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n29976), 
            .D(n38), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n29976), 
            .D(n39), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n29976), 
            .D(n40), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n29976), 
            .D(n41), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n29976), 
            .D(n42), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n29976), 
            .D(n43), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2039__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n29976), 
            .D(n44), .R(n31159));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n62898));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n60846));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY add_1192_24 (.CI(n52651), .I0(GND_net), .I1(n11452), .CO(n52652));
    SB_LUT4 n9949_bdd_4_lut_52195 (.I0(n9949), .I1(current[0]), .I2(duty[3]), 
            .I3(n9947), .O(n71524));
    defparam n9949_bdd_4_lut_52195.LUT_INIT = 16'he4aa;
    SB_LUT4 n71524_bdd_4_lut (.I0(n71524), .I1(duty[0]), .I2(n4945), .I3(n9947), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n71524_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 add_1192_23_lut (.I0(GND_net), .I1(GND_net), .I2(n11454), 
            .I3(n52650), .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n52558), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n52559));
    SB_CARRY add_1192_23 (.CI(n52650), .I0(GND_net), .I1(n11454), .CO(n52651));
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n52539), .O(n1241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_12 (.CI(n52539), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n52540));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n52557), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_22_lut (.I0(GND_net), .I1(GND_net), .I2(n11456), 
            .I3(n52649), .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_22 (.CI(n52649), .I0(GND_net), .I1(n11456), .CO(n52650));
    SB_LUT4 add_1192_21_lut (.I0(GND_net), .I1(GND_net), .I2(n11458), 
            .I3(n52648), .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_30 (.CI(n52557), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n52558));
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n52538), .O(n1242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_21 (.CI(n52648), .I0(GND_net), .I1(n11458), .CO(n52649));
    SB_LUT4 add_1192_20_lut (.I0(GND_net), .I1(GND_net), .I2(n11460), 
            .I3(n52647), .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_20 (.CI(n52647), .I0(GND_net), .I1(n11460), .CO(n52648));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n52556), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_29 (.CI(n52556), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n52557));
    SB_LUT4 add_1192_19_lut (.I0(GND_net), .I1(GND_net), .I2(n11462), 
            .I3(n52646), .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n52531), .O(n1249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_19 (.CI(n52646), .I0(GND_net), .I1(n11462), .CO(n52647));
    SB_LUT4 add_1192_18_lut (.I0(GND_net), .I1(GND_net), .I2(n11464), 
            .I3(n52645), .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_18 (.CI(n52645), .I0(GND_net), .I1(n11464), .CO(n52646));
    SB_LUT4 i13902_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n60038), .I3(GND_net), .O(n31847));   // verilog/coms.v(130[12] 305[6])
    defparam i13902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1192_17_lut (.I0(GND_net), .I1(GND_net), .I2(n11466), 
            .I3(n52644), .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_17 (.CI(n52644), .I0(GND_net), .I1(n11466), .CO(n52645));
    SB_LUT4 add_1192_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11468), 
            .I3(n52643), .O(n4931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_16 (.CI(n52643), .I0(GND_net), .I1(n11468), .CO(n52644));
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n29830), 
            .D(n1251), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_CARRY add_151_11 (.CI(n52538), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n52539));
    SB_LUT4 add_1192_15_lut (.I0(GND_net), .I1(GND_net), .I2(n11470), 
            .I3(n52642), .O(n4932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_15 (.CI(n52642), .I0(GND_net), .I1(n11470), .CO(n52643));
    SB_LUT4 add_1192_14_lut (.I0(GND_net), .I1(GND_net), .I2(n11472), 
            .I3(n52641), .O(n4933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n52537), .O(n1243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n52555), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_28 (.CI(n52555), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n52556));
    SB_CARRY add_1192_14 (.CI(n52641), .I0(GND_net), .I1(n11472), .CO(n52642));
    SB_LUT4 add_1192_13_lut (.I0(GND_net), .I1(GND_net), .I2(n11474), 
            .I3(n52640), .O(n4934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n52554), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1679_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n11452));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i23_3_lut.LUT_INIT = 16'h3535;
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n29752), .D(GHC_N_391), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_1192_13 (.CI(n52640), .I0(GND_net), .I1(n11474), .CO(n52641));
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n29752), .D(GHB_N_377), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n29752), .D(GHA_N_355), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5852), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n29752), .D(GLA_N_372), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n29752), .D(GLB_N_386), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_151_27 (.CI(n52554), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n52555));
    SB_LUT4 add_1192_12_lut (.I0(GND_net), .I1(GND_net), .I2(n11476), 
            .I3(n52639), .O(n4935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_12 (.CI(n52639), .I0(GND_net), .I1(n11476), .CO(n52640));
    SB_LUT4 add_1192_11_lut (.I0(GND_net), .I1(GND_net), .I2(n11478), 
            .I3(n52638), .O(n4936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_11 (.CI(n52638), .I0(GND_net), .I1(n11478), .CO(n52639));
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n29752), .D(GLC_N_400), 
            .R(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_151_4 (.CI(n52531), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n52532));
    SB_CARRY add_151_10 (.CI(n52537), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n52538));
    SB_LUT4 encoder1_position_31__I_0_add_2126_32_lut (.I0(encoder1_position[31]), 
            .I1(n11885), .I2(GND_net), .I3(n53886), .O(encoder1_position_scaled_23__N_43[31])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder1_position_31__I_0_add_2126_31_lut (.I0(GND_net), .I1(n11886), 
            .I2(encoder1_position[30]), .I3(n53885), .O(encoder1_position_scaled_23__N_43[30])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_31 (.CI(n53885), .I0(n11886), 
            .I1(encoder1_position[30]), .CO(n53886));
    SB_LUT4 encoder1_position_31__I_0_add_2126_30_lut (.I0(GND_net), .I1(n11887), 
            .I2(encoder1_position[29]), .I3(n53884), .O(encoder1_position_scaled_23__N_43[29])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_30_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n52553), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13737_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3180), .I3(GND_net), 
            .O(n31682));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13738_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3180), .I3(GND_net), 
            .O(n31683));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13738_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_151_26 (.CI(n52553), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n52554));
    SB_LUT4 mux_245_i6_4_lut (.I0(displacement[5]), .I1(encoder0_position_scaled[5]), 
            .I2(n54181), .I3(n51206), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'hf353;
    SB_CARRY encoder1_position_31__I_0_add_2126_30 (.CI(n53884), .I0(n11887), 
            .I1(encoder1_position[29]), .CO(n53885));
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n52536), .O(n1244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13739_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3180), .I3(GND_net), 
            .O(n31684));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45536_3_lut (.I0(n4925), .I1(duty[20]), .I2(n9949), .I3(GND_net), 
            .O(n64806));
    defparam i45536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_29_lut (.I0(GND_net), .I1(n11888), 
            .I2(encoder1_position[28]), .I3(n53883), .O(encoder1_position_scaled_23__N_43[28])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_29 (.CI(n53883), .I0(n11888), 
            .I1(encoder1_position[28]), .CO(n53884));
    SB_LUT4 add_1192_10_lut (.I0(GND_net), .I1(GND_net), .I2(n11480), 
            .I3(n52637), .O(n4937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_10 (.CI(n52637), .I0(GND_net), .I1(n11480), .CO(n52638));
    SB_LUT4 encoder1_position_31__I_0_add_2126_28_lut (.I0(GND_net), .I1(n11889), 
            .I2(encoder1_position[27]), .I3(n53882), .O(encoder1_position_scaled_23__N_43[27])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n52552), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_25 (.CI(n52552), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n52553));
    SB_LUT4 add_1192_9_lut (.I0(GND_net), .I1(GND_net), .I2(n11482), .I3(n52636), 
            .O(n4938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_28 (.CI(n53882), .I0(n11889), 
            .I1(encoder1_position[27]), .CO(n53883));
    SB_LUT4 encoder1_position_31__I_0_add_2126_27_lut (.I0(GND_net), .I1(n11890), 
            .I2(encoder1_position[26]), .I3(n53881), .O(encoder1_position_scaled_23__N_43[26])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_9 (.CI(n52536), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n52537));
    SB_CARRY add_1192_9 (.CI(n52636), .I0(GND_net), .I1(n11482), .CO(n52637));
    SB_CARRY encoder1_position_31__I_0_add_2126_27 (.CI(n53881), .I0(n11890), 
            .I1(encoder1_position[26]), .CO(n53882));
    SB_LUT4 encoder1_position_31__I_0_add_2126_26_lut (.I0(GND_net), .I1(n11891), 
            .I2(encoder1_position[25]), .I3(n53880), .O(encoder1_position_scaled_23__N_43[25])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_26 (.CI(n53880), .I0(n11891), 
            .I1(encoder1_position[25]), .CO(n53881));
    SB_LUT4 encoder1_position_31__I_0_add_2126_25_lut (.I0(GND_net), .I1(n11892), 
            .I2(encoder1_position[24]), .I3(n53879), .O(encoder1_position_scaled_23__N_43[24])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_25 (.CI(n53879), .I0(n11892), 
            .I1(encoder1_position[24]), .CO(n53880));
    SB_LUT4 encoder1_position_31__I_0_add_2126_24_lut (.I0(GND_net), .I1(n11893), 
            .I2(encoder1_position[23]), .I3(n53878), .O(encoder1_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_24 (.CI(n53878), .I0(n11893), 
            .I1(encoder1_position[23]), .CO(n53879));
    SB_LUT4 encoder1_position_31__I_0_add_2126_23_lut (.I0(GND_net), .I1(n11894), 
            .I2(encoder1_position[22]), .I3(n53877), .O(encoder1_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_23 (.CI(n53877), .I0(n11894), 
            .I1(encoder1_position[22]), .CO(n53878));
    SB_LUT4 encoder1_position_31__I_0_add_2126_22_lut (.I0(GND_net), .I1(n11895), 
            .I2(encoder1_position[21]), .I3(n53876), .O(encoder1_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_22 (.CI(n53876), .I0(n11895), 
            .I1(encoder1_position[21]), .CO(n53877));
    SB_LUT4 encoder1_position_31__I_0_add_2126_21_lut (.I0(GND_net), .I1(n11896), 
            .I2(encoder1_position[20]), .I3(n53875), .O(encoder1_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_21 (.CI(n53875), .I0(n11896), 
            .I1(encoder1_position[20]), .CO(n53876));
    SB_LUT4 add_1192_8_lut (.I0(GND_net), .I1(GND_net), .I2(n11484), .I3(n52635), 
            .O(n4939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_31__I_0_add_2126_20_lut (.I0(GND_net), .I1(n11897), 
            .I2(encoder1_position[19]), .I3(n53874), .O(encoder1_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_20 (.CI(n53874), .I0(n11897), 
            .I1(encoder1_position[19]), .CO(n53875));
    SB_LUT4 i45538_3_lut (.I0(n64806), .I1(n64804), .I2(n9947), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i45538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45533_3_lut (.I0(n4924), .I1(duty[21]), .I2(n9949), .I3(GND_net), 
            .O(n64803));
    defparam i45533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_19_lut (.I0(GND_net), .I1(n11898), 
            .I2(encoder1_position[18]), .I3(n53873), .O(encoder1_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45535_3_lut (.I0(n64803), .I1(n64804), .I2(n9947), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i45535_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_31__I_0_add_2126_19 (.CI(n53873), .I0(n11898), 
            .I1(encoder1_position[18]), .CO(n53874));
    SB_LUT4 encoder1_position_31__I_0_add_2126_18_lut (.I0(GND_net), .I1(n11899), 
            .I2(encoder1_position[17]), .I3(n53872), .O(encoder1_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_18 (.CI(n53872), .I0(n11899), 
            .I1(encoder1_position[17]), .CO(n53873));
    SB_LUT4 i45534_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n9949), 
            .I3(GND_net), .O(n64804));
    defparam i45534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_17_lut (.I0(GND_net), .I1(n11900), 
            .I2(encoder1_position[16]), .I3(n53871), .O(encoder1_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_17 (.CI(n53871), .I0(n11900), 
            .I1(encoder1_position[16]), .CO(n53872));
    SB_LUT4 encoder1_position_31__I_0_add_2126_16_lut (.I0(GND_net), .I1(n11901), 
            .I2(encoder1_position[15]), .I3(n53870), .O(encoder1_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_16 (.CI(n53870), .I0(n11901), 
            .I1(encoder1_position[15]), .CO(n53871));
    SB_LUT4 encoder1_position_31__I_0_add_2126_15_lut (.I0(GND_net), .I1(n11902), 
            .I2(encoder1_position[14]), .I3(n53869), .O(encoder1_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_15 (.CI(n53869), .I0(n11902), 
            .I1(encoder1_position[14]), .CO(n53870));
    SB_LUT4 i45530_3_lut (.I0(n4923), .I1(duty[22]), .I2(n9949), .I3(GND_net), 
            .O(n64800));
    defparam i45530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_14_lut (.I0(GND_net), .I1(n11903), 
            .I2(encoder1_position[13]), .I3(n53868), .O(encoder1_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_14 (.CI(n53868), .I0(n11903), 
            .I1(encoder1_position[13]), .CO(n53869));
    SB_LUT4 encoder1_position_31__I_0_add_2126_13_lut (.I0(GND_net), .I1(n11904), 
            .I2(encoder1_position[12]), .I3(n53867), .O(encoder1_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_13 (.CI(n53867), .I0(n11904), 
            .I1(encoder1_position[12]), .CO(n53868));
    SB_LUT4 i45532_3_lut (.I0(n64800), .I1(n64804), .I2(n9947), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i45532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_12_lut (.I0(GND_net), .I1(n11905), 
            .I2(encoder1_position[11]), .I3(n53866), .O(encoder1_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_12 (.CI(n53866), .I0(n11905), 
            .I1(encoder1_position[11]), .CO(n53867));
    SB_LUT4 encoder1_position_31__I_0_add_2126_11_lut (.I0(GND_net), .I1(n11906), 
            .I2(encoder1_position[10]), .I3(n53865), .O(encoder1_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_11 (.CI(n53865), .I0(n11906), 
            .I1(encoder1_position[10]), .CO(n53866));
    SB_LUT4 i6170_3_lut (.I0(n4922), .I1(current[15]), .I2(n9947), .I3(GND_net), 
            .O(n23767));
    defparam i6170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_10_lut (.I0(GND_net), .I1(n11907), 
            .I2(encoder1_position[9]), .I3(n53864), .O(encoder1_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_10 (.CI(n53864), .I0(n11907), 
            .I1(encoder1_position[9]), .CO(n53865));
    SB_LUT4 i6171_3_lut (.I0(n23767), .I1(duty[23]), .I2(n9949), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i6171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_31__I_0_add_2126_9_lut (.I0(GND_net), .I1(n11908), 
            .I2(encoder1_position[8]), .I3(n53863), .O(encoder1_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_9 (.CI(n53863), .I0(n11908), 
            .I1(encoder1_position[8]), .CO(n53864));
    SB_CARRY encoder1_position_31__I_0_add_2126_8 (.CI(n53862), .I0(n11909), 
            .I1(encoder1_position[7]), .CO(n53863));
    SB_CARRY encoder1_position_31__I_0_add_2126_7 (.CI(n53861), .I0(n11910), 
            .I1(encoder1_position[6]), .CO(n53862));
    SB_CARRY encoder1_position_31__I_0_add_2126_6 (.CI(n53860), .I0(n11911), 
            .I1(encoder1_position[5]), .CO(n53861));
    SB_CARRY encoder1_position_31__I_0_add_2126_5 (.CI(n53859), .I0(n11912), 
            .I1(encoder1_position[4]), .CO(n53860));
    SB_CARRY encoder1_position_31__I_0_add_2126_4 (.CI(n53858), .I0(n11913), 
            .I1(encoder1_position[3]), .CO(n53859));
    SB_CARRY encoder1_position_31__I_0_add_2126_3 (.CI(n53857), .I0(n11914), 
            .I1(encoder1_position[2]), .CO(n53858));
    SB_CARRY encoder1_position_31__I_0_add_2126_2 (.CI(GND_net), .I0(encoder1_position[0]), 
            .I1(encoder1_position[1]), .CO(n53857));
    SB_LUT4 add_4946_31_lut (.I0(GND_net), .I1(n13508), .I2(encoder1_position[30]), 
            .I3(n53856), .O(n11885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4946_30_lut (.I0(GND_net), .I1(n13509), .I2(encoder1_position[29]), 
            .I3(n53855), .O(n11886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_30 (.CI(n53855), .I0(n13509), .I1(encoder1_position[29]), 
            .CO(n53856));
    SB_LUT4 add_4946_29_lut (.I0(GND_net), .I1(n13510), .I2(encoder1_position[28]), 
            .I3(n53854), .O(n11887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_29 (.CI(n53854), .I0(n13510), .I1(encoder1_position[28]), 
            .CO(n53855));
    SB_LUT4 add_4946_28_lut (.I0(GND_net), .I1(n13511), .I2(encoder1_position[27]), 
            .I3(n53853), .O(n11888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14746_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n32691));   // verilog/coms.v(130[12] 305[6])
    defparam i14746_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4946_28 (.CI(n53853), .I0(n13511), .I1(encoder1_position[27]), 
            .CO(n53854));
    SB_LUT4 add_4946_27_lut (.I0(GND_net), .I1(n13512), .I2(encoder1_position[26]), 
            .I3(n53852), .O(n11889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_27 (.CI(n53852), .I0(n13512), .I1(encoder1_position[26]), 
            .CO(n53853));
    SB_LUT4 i13740_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3180), .I3(GND_net), 
            .O(n31685));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4946_26_lut (.I0(GND_net), .I1(n13513), .I2(encoder1_position[25]), 
            .I3(n53851), .O(n11890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_26 (.CI(n53851), .I0(n13513), .I1(encoder1_position[25]), 
            .CO(n53852));
    SB_LUT4 add_4946_25_lut (.I0(GND_net), .I1(n13514), .I2(encoder1_position[24]), 
            .I3(n53850), .O(n11891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_25 (.CI(n53850), .I0(n13514), .I1(encoder1_position[24]), 
            .CO(n53851));
    SB_LUT4 add_4946_24_lut (.I0(GND_net), .I1(n13515), .I2(encoder1_position[23]), 
            .I3(n53849), .O(n11892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_24 (.CI(n53849), .I0(n13515), .I1(encoder1_position[23]), 
            .CO(n53850));
    SB_LUT4 add_4946_23_lut (.I0(GND_net), .I1(n13516), .I2(encoder1_position[22]), 
            .I3(n53848), .O(n11893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_23 (.CI(n53848), .I0(n13516), .I1(encoder1_position[22]), 
            .CO(n53849));
    SB_LUT4 add_4946_22_lut (.I0(GND_net), .I1(n13517), .I2(encoder1_position[21]), 
            .I3(n53847), .O(n11894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_22 (.CI(n53847), .I0(n13517), .I1(encoder1_position[21]), 
            .CO(n53848));
    SB_LUT4 add_4946_21_lut (.I0(GND_net), .I1(n13518), .I2(encoder1_position[20]), 
            .I3(n53846), .O(n11895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_21 (.CI(n53846), .I0(n13518), .I1(encoder1_position[20]), 
            .CO(n53847));
    SB_LUT4 add_4946_20_lut (.I0(GND_net), .I1(n13519), .I2(encoder1_position[19]), 
            .I3(n53845), .O(n11896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_20 (.CI(n53845), .I0(n13519), .I1(encoder1_position[19]), 
            .CO(n53846));
    SB_LUT4 add_4946_19_lut (.I0(GND_net), .I1(n13520), .I2(encoder1_position[18]), 
            .I3(n53844), .O(n11897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_19 (.CI(n53844), .I0(n13520), .I1(encoder1_position[18]), 
            .CO(n53845));
    SB_LUT4 add_4946_18_lut (.I0(GND_net), .I1(n13521), .I2(encoder1_position[17]), 
            .I3(n53843), .O(n11898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_18 (.CI(n53843), .I0(n13521), .I1(encoder1_position[17]), 
            .CO(n53844));
    SB_LUT4 add_4946_17_lut (.I0(GND_net), .I1(n13522), .I2(encoder1_position[16]), 
            .I3(n53842), .O(n11899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_17 (.CI(n53842), .I0(n13522), .I1(encoder1_position[16]), 
            .CO(n53843));
    SB_LUT4 add_4946_16_lut (.I0(GND_net), .I1(n13523), .I2(encoder1_position[15]), 
            .I3(n53841), .O(n11900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_16 (.CI(n53841), .I0(n13523), .I1(encoder1_position[15]), 
            .CO(n53842));
    SB_LUT4 add_4946_15_lut (.I0(GND_net), .I1(n13524), .I2(encoder1_position[14]), 
            .I3(n53840), .O(n11901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_15 (.CI(n53840), .I0(n13524), .I1(encoder1_position[14]), 
            .CO(n53841));
    SB_LUT4 add_4946_14_lut (.I0(GND_net), .I1(n13525), .I2(encoder1_position[13]), 
            .I3(n53839), .O(n11902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_14 (.CI(n53839), .I0(n13525), .I1(encoder1_position[13]), 
            .CO(n53840));
    SB_LUT4 add_4946_13_lut (.I0(GND_net), .I1(n13526), .I2(encoder1_position[12]), 
            .I3(n53838), .O(n11903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_13 (.CI(n53838), .I0(n13526), .I1(encoder1_position[12]), 
            .CO(n53839));
    SB_LUT4 add_4946_12_lut (.I0(GND_net), .I1(n13527), .I2(encoder1_position[11]), 
            .I3(n53837), .O(n11904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_12 (.CI(n53837), .I0(n13527), .I1(encoder1_position[11]), 
            .CO(n53838));
    SB_LUT4 add_4946_11_lut (.I0(GND_net), .I1(n13528), .I2(encoder1_position[10]), 
            .I3(n53836), .O(n11905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_11 (.CI(n53836), .I0(n13528), .I1(encoder1_position[10]), 
            .CO(n53837));
    SB_LUT4 add_4946_10_lut (.I0(GND_net), .I1(n13529), .I2(encoder1_position[9]), 
            .I3(n53835), .O(n11906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13741_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3180), .I3(GND_net), 
            .O(n31686));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13741_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4946_10 (.CI(n53835), .I0(n13529), .I1(encoder1_position[9]), 
            .CO(n53836));
    SB_LUT4 add_4946_9_lut (.I0(GND_net), .I1(n13530), .I2(encoder1_position[8]), 
            .I3(n53834), .O(n11907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_9 (.CI(n53834), .I0(n13530), .I1(encoder1_position[8]), 
            .CO(n53835));
    SB_LUT4 add_4946_8_lut (.I0(GND_net), .I1(n13531), .I2(encoder1_position[7]), 
            .I3(n53833), .O(n11908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_8 (.CI(n53833), .I0(n13531), .I1(encoder1_position[7]), 
            .CO(n53834));
    SB_LUT4 add_4946_7_lut (.I0(GND_net), .I1(n13532), .I2(encoder1_position[6]), 
            .I3(n53832), .O(n11909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_7 (.CI(n53832), .I0(n13532), .I1(encoder1_position[6]), 
            .CO(n53833));
    SB_LUT4 add_4946_6_lut (.I0(GND_net), .I1(n13533), .I2(encoder1_position[5]), 
            .I3(n53831), .O(n11910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_6 (.CI(n53831), .I0(n13533), .I1(encoder1_position[5]), 
            .CO(n53832));
    SB_LUT4 add_4946_5_lut (.I0(GND_net), .I1(n13534), .I2(encoder1_position[4]), 
            .I3(n53830), .O(n11911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_5 (.CI(n53830), .I0(n13534), .I1(encoder1_position[4]), 
            .CO(n53831));
    SB_LUT4 add_4946_4_lut (.I0(GND_net), .I1(n13535), .I2(encoder1_position[3]), 
            .I3(n53829), .O(n11912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_4 (.CI(n53829), .I0(n13535), .I1(encoder1_position[3]), 
            .CO(n53830));
    SB_LUT4 add_4946_3_lut (.I0(GND_net), .I1(n13536), .I2(encoder1_position[2]), 
            .I3(n53828), .O(n11913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_3 (.CI(n53828), .I0(n13536), .I1(encoder1_position[2]), 
            .CO(n53829));
    SB_LUT4 add_4946_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n11914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4946_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4946_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n53828));
    SB_LUT4 i1_3_lut (.I0(n23_adj_5843), .I1(o_Rx_DV_N_3488[12]), .I2(n5235), 
            .I3(GND_net), .O(n63019));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), .I3(n63019), 
            .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_1183_i15_2_lut (.I0(r_Clock_Count_adj_5928[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5817));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1183_i9_2_lut (.I0(r_Clock_Count_adj_5928[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5813));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1183_i11_2_lut (.I0(r_Clock_Count_adj_5928[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5814));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1183_i13_2_lut (.I0(r_Clock_Count_adj_5928[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5815));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5012_30_lut (.I0(GND_net), .I1(n14971), .I2(encoder1_position[29]), 
            .I3(n53827), .O(n13508)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5012_29_lut (.I0(GND_net), .I1(n14972), .I2(encoder1_position[28]), 
            .I3(n53826), .O(n13509)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_29 (.CI(n53826), .I0(n14972), .I1(encoder1_position[28]), 
            .CO(n53827));
    SB_LUT4 add_5012_28_lut (.I0(GND_net), .I1(n14973), .I2(encoder1_position[27]), 
            .I3(n53825), .O(n13510)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_28 (.CI(n53825), .I0(n14973), .I1(encoder1_position[27]), 
            .CO(n53826));
    SB_LUT4 add_5012_27_lut (.I0(GND_net), .I1(n14974), .I2(encoder1_position[26]), 
            .I3(n53824), .O(n13511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_27 (.CI(n53824), .I0(n14974), .I1(encoder1_position[26]), 
            .CO(n53825));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 LessThan_1183_i4_4_lut (.I0(r_Clock_Count_adj_5928[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5928[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5810));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 add_5012_26_lut (.I0(GND_net), .I1(n14975), .I2(encoder1_position[25]), 
            .I3(n53823), .O(n13512)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_26 (.CI(n53823), .I0(n14975), .I1(encoder1_position[25]), 
            .CO(n53824));
    SB_CARRY add_1192_8 (.CI(n52635), .I0(GND_net), .I1(n11484), .CO(n52636));
    SB_LUT4 add_5012_25_lut (.I0(GND_net), .I1(n14976), .I2(encoder1_position[24]), 
            .I3(n53822), .O(n13513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51120_3_lut (.I0(n4_adj_5810), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5814), 
            .I3(GND_net), .O(n70390));   // verilog/uart_tx.v(117[17:57])
    defparam i51120_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5012_25 (.CI(n53822), .I0(n14976), .I1(encoder1_position[24]), 
            .CO(n53823));
    SB_LUT4 add_5012_24_lut (.I0(GND_net), .I1(n14977), .I2(encoder1_position[23]), 
            .I3(n53821), .O(n13514)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_24 (.CI(n53821), .I0(n14977), .I1(encoder1_position[23]), 
            .CO(n53822));
    SB_LUT4 add_5012_23_lut (.I0(GND_net), .I1(n14978), .I2(encoder1_position[22]), 
            .I3(n53820), .O(n13515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_7_lut (.I0(GND_net), .I1(GND_net), .I2(n11486), .I3(n52634), 
            .O(n4940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[31]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[30]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[29]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[28]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[27]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[26]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[25]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[24]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_CARRY add_5012_23 (.CI(n53820), .I0(n14978), .I1(encoder1_position[22]), 
            .CO(n53821));
    SB_LUT4 i51121_3_lut (.I0(n70390), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5815), 
            .I3(GND_net), .O(n70391));   // verilog/uart_tx.v(117[17:57])
    defparam i51121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49559_4_lut (.I0(n13_adj_5815), .I1(n11_adj_5814), .I2(n9_adj_5813), 
            .I3(n67830), .O(n68829));
    defparam i49559_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1183_i8_3_lut (.I0(n6_adj_5811), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5813), .I3(GND_net), .O(n8_adj_5812));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1183_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5012_22_lut (.I0(GND_net), .I1(n14979), .I2(encoder1_position[21]), 
            .I3(n53819), .O(n13516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_22 (.CI(n53819), .I0(n14979), .I1(encoder1_position[21]), 
            .CO(n53820));
    SB_LUT4 add_5012_21_lut (.I0(GND_net), .I1(n14980), .I2(encoder1_position[20]), 
            .I3(n53818), .O(n13517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_21 (.CI(n53818), .I0(n14980), .I1(encoder1_position[20]), 
            .CO(n53819));
    SB_LUT4 add_5012_20_lut (.I0(GND_net), .I1(n14981), .I2(encoder1_position[19]), 
            .I3(n53817), .O(n13518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_20 (.CI(n53817), .I0(n14981), .I1(encoder1_position[19]), 
            .CO(n53818));
    SB_LUT4 add_5012_19_lut (.I0(GND_net), .I1(n14982), .I2(encoder1_position[18]), 
            .I3(n53816), .O(n13519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_19 (.CI(n53816), .I0(n14982), .I1(encoder1_position[18]), 
            .CO(n53817));
    SB_LUT4 i50916_3_lut (.I0(n70391), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5817), 
            .I3(GND_net), .O(n14_adj_5816));   // verilog/uart_tx.v(117[17:57])
    defparam i50916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5012_18_lut (.I0(GND_net), .I1(n14983), .I2(encoder1_position[17]), 
            .I3(n53815), .O(n13520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_18 (.CI(n53815), .I0(n14983), .I1(encoder1_position[17]), 
            .CO(n53816));
    SB_LUT4 add_5012_17_lut (.I0(GND_net), .I1(n14984), .I2(encoder1_position[16]), 
            .I3(n53814), .O(n13521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_17 (.CI(n53814), .I0(n14984), .I1(encoder1_position[16]), 
            .CO(n53815));
    SB_LUT4 add_5012_16_lut (.I0(GND_net), .I1(n14985), .I2(encoder1_position[15]), 
            .I3(n53813), .O(n13522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_16 (.CI(n53813), .I0(n14985), .I1(encoder1_position[15]), 
            .CO(n53814));
    SB_LUT4 i50552_4_lut (.I0(n14_adj_5816), .I1(n8_adj_5812), .I2(n15_adj_5817), 
            .I3(n68829), .O(n69822));   // verilog/uart_tx.v(117[17:57])
    defparam i50552_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50553_3_lut (.I0(n69822), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5928[8]), 
            .I3(GND_net), .O(n5235));   // verilog/uart_tx.v(117[17:57])
    defparam i50553_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5012_15_lut (.I0(GND_net), .I1(n14986), .I2(encoder1_position[14]), 
            .I3(n53812), .O(n13523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_15 (.CI(n53812), .I0(n14986), .I1(encoder1_position[14]), 
            .CO(n53813));
    SB_CARRY add_1192_7 (.CI(n52634), .I0(GND_net), .I1(n11486), .CO(n52635));
    SB_LUT4 i1_3_lut_adj_1792 (.I0(o_Rx_DV_N_3488[12]), .I1(n5235), .I2(n59688), 
            .I3(GND_net), .O(n63181));
    defparam i1_3_lut_adj_1792.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63181), .O(n63187));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5012_14_lut (.I0(GND_net), .I1(n14987), .I2(encoder1_position[13]), 
            .I3(n53811), .O(n13524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_14 (.CI(n53811), .I0(n14987), .I1(encoder1_position[13]), 
            .CO(n53812));
    SB_LUT4 add_5012_13_lut (.I0(GND_net), .I1(n14988), .I2(encoder1_position[12]), 
            .I3(n53810), .O(n13525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_13 (.CI(n53810), .I0(n14988), .I1(encoder1_position[12]), 
            .CO(n53811));
    SB_LUT4 add_5012_12_lut (.I0(GND_net), .I1(n14989), .I2(encoder1_position[11]), 
            .I3(n53809), .O(n13526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_12 (.CI(n53809), .I0(n14989), .I1(encoder1_position[11]), 
            .CO(n53810));
    SB_LUT4 add_5012_11_lut (.I0(GND_net), .I1(n14990), .I2(encoder1_position[10]), 
            .I3(n53808), .O(n13527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_11 (.CI(n53808), .I0(n14990), .I1(encoder1_position[10]), 
            .CO(n53809));
    SB_LUT4 add_5012_10_lut (.I0(GND_net), .I1(n14991), .I2(encoder1_position[9]), 
            .I3(n53807), .O(n13528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_10 (.CI(n53807), .I0(n14991), .I1(encoder1_position[9]), 
            .CO(n53808));
    SB_LUT4 add_5012_9_lut (.I0(GND_net), .I1(n14992), .I2(encoder1_position[8]), 
            .I3(n53806), .O(n13529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_9 (.CI(n53806), .I0(n14992), .I1(encoder1_position[8]), 
            .CO(n53807));
    SB_LUT4 add_5012_8_lut (.I0(GND_net), .I1(n14993), .I2(encoder1_position[7]), 
            .I3(n53805), .O(n13530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_8 (.CI(n53805), .I0(n14993), .I1(encoder1_position[7]), 
            .CO(n53806));
    SB_LUT4 add_5012_7_lut (.I0(GND_net), .I1(n14994), .I2(encoder1_position[6]), 
            .I3(n53804), .O(n13531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_7 (.CI(n53804), .I0(n14994), .I1(encoder1_position[6]), 
            .CO(n53805));
    SB_LUT4 add_5012_6_lut (.I0(GND_net), .I1(n14995), .I2(encoder1_position[5]), 
            .I3(n53803), .O(n13532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_6 (.CI(n53803), .I0(n14995), .I1(encoder1_position[5]), 
            .CO(n53804));
    SB_LUT4 add_5012_5_lut (.I0(GND_net), .I1(n14996), .I2(encoder1_position[4]), 
            .I3(n53802), .O(n13533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_5 (.CI(n53802), .I0(n14996), .I1(encoder1_position[4]), 
            .CO(n53803));
    SB_LUT4 add_5012_4_lut (.I0(GND_net), .I1(n14997), .I2(encoder1_position[3]), 
            .I3(n53801), .O(n13534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_4 (.CI(n53801), .I0(n14997), .I1(encoder1_position[3]), 
            .CO(n53802));
    SB_LUT4 i45431_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64701));
    defparam i45431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45432_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64702));
    defparam i45432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i2_4_lut (.I0(displacement[1]), .I1(encoder0_position_scaled[1]), 
            .I2(n54181), .I3(n51206), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_2_lut_adj_1794 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60741));
    defparam i1_2_lut_adj_1794.LUT_INIT = 16'h6666;
    SB_LUT4 i45423_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64693));
    defparam i45423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45422_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64692));
    defparam i45422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1192_6_lut (.I0(GND_net), .I1(GND_net), .I2(n11488), .I3(n52633), 
            .O(n4941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n52551), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_6 (.CI(n52633), .I0(GND_net), .I1(n11488), .CO(n52634));
    SB_LUT4 add_5012_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n53800), .O(n13535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n58068));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_CARRY add_5012_3 (.CI(n53800), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n53801));
    SB_LUT4 add_5012_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n13536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_5_lut (.I0(GND_net), .I1(GND_net), .I2(n11490), .I3(n52632), 
            .O(n4942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1192_5 (.CI(n52632), .I0(GND_net), .I1(n11490), .CO(n52633));
    SB_CARRY add_5012_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n53800));
    SB_LUT4 add_5185_28_lut (.I0(GND_net), .I1(n17449), .I2(encoder1_position[28]), 
            .I3(n53799), .O(n14971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_27_lut (.I0(GND_net), .I1(n17450), .I2(encoder1_position[27]), 
            .I3(n53798), .O(n14972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_27 (.CI(n53798), .I0(n17450), .I1(encoder1_position[27]), 
            .CO(n53799));
    SB_LUT4 add_5185_26_lut (.I0(GND_net), .I1(n17451), .I2(encoder1_position[26]), 
            .I3(n53797), .O(n14973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_26 (.CI(n53797), .I0(n17451), .I1(encoder1_position[26]), 
            .CO(n53798));
    SB_LUT4 add_5185_25_lut (.I0(GND_net), .I1(n17452), .I2(encoder1_position[25]), 
            .I3(n53796), .O(n14974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_25 (.CI(n53796), .I0(n17452), .I1(encoder1_position[25]), 
            .CO(n53797));
    SB_LUT4 add_5185_24_lut (.I0(GND_net), .I1(n17453), .I2(encoder1_position[24]), 
            .I3(n53795), .O(n14975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1192_4_lut (.I0(GND_net), .I1(GND_net), .I2(n11492), .I3(n52631), 
            .O(n4943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n52551), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n52552));
    SB_CARRY add_1192_4 (.CI(n52631), .I0(GND_net), .I1(n11492), .CO(n52632));
    SB_LUT4 mux_245_i7_4_lut (.I0(displacement[6]), .I1(encoder0_position_scaled[6]), 
            .I2(n54181), .I3(n51206), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 add_1192_3_lut (.I0(GND_net), .I1(GND_net), .I2(n11494), .I3(n52630), 
            .O(n4944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_24 (.CI(n53795), .I0(n17453), .I1(encoder1_position[24]), 
            .CO(n53796));
    SB_CARRY add_1192_3 (.CI(n52630), .I0(GND_net), .I1(n11494), .CO(n52631));
    SB_LUT4 add_1192_2_lut (.I0(GND_net), .I1(GND_net), .I2(n10012), .I3(VCC_net), 
            .O(n4945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1192_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_23_lut (.I0(GND_net), .I1(n17454), .I2(encoder1_position[23]), 
            .I3(n53794), .O(n14976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_23 (.CI(n53794), .I0(n17454), .I1(encoder1_position[23]), 
            .CO(n53795));
    SB_LUT4 add_5185_22_lut (.I0(GND_net), .I1(n17455), .I2(encoder1_position[22]), 
            .I3(n53793), .O(n14977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_22 (.CI(n53793), .I0(n17455), .I1(encoder1_position[22]), 
            .CO(n53794));
    SB_LUT4 mux_245_i3_4_lut (.I0(displacement[2]), .I1(encoder0_position_scaled[2]), 
            .I2(n54181), .I3(n51206), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 add_5185_21_lut (.I0(GND_net), .I1(n17456), .I2(encoder1_position[21]), 
            .I3(n53792), .O(n14978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_21 (.CI(n53792), .I0(n17456), .I1(encoder1_position[21]), 
            .CO(n53793));
    SB_LUT4 add_5185_20_lut (.I0(GND_net), .I1(n17457), .I2(encoder1_position[20]), 
            .I3(n53791), .O(n14979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_20 (.CI(n53791), .I0(n17457), .I1(encoder1_position[20]), 
            .CO(n53792));
    SB_CARRY add_1192_2 (.CI(VCC_net), .I0(GND_net), .I1(n10012), .CO(n52630));
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n29830), 
            .D(n1250), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n29830), 
            .D(n1249), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n29830), 
            .D(n1248), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 add_5185_19_lut (.I0(GND_net), .I1(n17458), .I2(encoder1_position[19]), 
            .I3(n53790), .O(n14980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_19 (.CI(n53790), .I0(n17458), .I1(encoder1_position[19]), 
            .CO(n53791));
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n29830), 
            .D(n1247), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n29830), 
            .D(n1246), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 add_5185_18_lut (.I0(GND_net), .I1(n17459), .I2(encoder1_position[18]), 
            .I3(n53789), .O(n14981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_18 (.CI(n53789), .I0(n17459), .I1(encoder1_position[18]), 
            .CO(n53790));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n52550), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_17_lut (.I0(GND_net), .I1(n17460), .I2(encoder1_position[17]), 
            .I3(n53788), .O(n14982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_17 (.CI(n53788), .I0(n17460), .I1(encoder1_position[17]), 
            .CO(n53789));
    SB_LUT4 i7_2_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28330));   // verilog/coms.v(100[12:26])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5185_16_lut (.I0(GND_net), .I1(n17461), .I2(encoder1_position[16]), 
            .I3(n53787), .O(n14983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_16 (.CI(n53787), .I0(n17461), .I1(encoder1_position[16]), 
            .CO(n53788));
    SB_LUT4 add_5185_15_lut (.I0(GND_net), .I1(n17462), .I2(encoder1_position[15]), 
            .I3(n53786), .O(n14984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n29830), 
            .D(n1245), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n29830), 
            .D(n1244), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n29830), 
            .D(n1243), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n29830), 
            .D(n1242), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n29830), 
            .D(n1241), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n29830), 
            .D(n1240), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n29830), 
            .D(n1239), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n29830), 
            .D(n1238), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n29830), 
            .D(n1237), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n29830), 
            .D(n1236), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n29830), 
            .D(n1235), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n29830), 
            .D(n1234), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n29830), 
            .D(n1233), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n29830), 
            .D(n1232), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n29830), 
            .D(n1231), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n29830), 
            .D(n1230), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n29830), 
            .D(n1229), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n29830), 
            .D(n1228), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n29830), 
            .D(n1227), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n29830), 
            .D(n1226), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n29830), 
            .D(n1225), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n29830), 
            .D(n1224), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n29830), 
            .D(n1223), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n29830), 
            .D(n1222), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n29830), 
            .D(n1221), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n29830), 
            .D(n1220), .R(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_CARRY add_151_23 (.CI(n52550), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n52551));
    SB_CARRY add_5185_15 (.CI(n53786), .I0(n17462), .I1(encoder1_position[15]), 
            .CO(n53787));
    SB_LUT4 add_5185_14_lut (.I0(GND_net), .I1(n17463), .I2(encoder1_position[14]), 
            .I3(n53785), .O(n14985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_14 (.CI(n53785), .I0(n17463), .I1(encoder1_position[14]), 
            .CO(n53786));
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n58154));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 add_5185_13_lut (.I0(GND_net), .I1(n17464), .I2(encoder1_position[13]), 
            .I3(n53784), .O(n14986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_5185_13 (.CI(n53784), .I0(n17464), .I1(encoder1_position[13]), 
            .CO(n53785));
    SB_LUT4 add_5185_12_lut (.I0(GND_net), .I1(n17465), .I2(encoder1_position[12]), 
            .I3(n53783), .O(n14987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_12 (.CI(n53783), .I0(n17465), .I1(encoder1_position[12]), 
            .CO(n53784));
    SB_LUT4 add_5185_11_lut (.I0(GND_net), .I1(n17466), .I2(encoder1_position[11]), 
            .I3(n53782), .O(n14988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_11 (.CI(n53782), .I0(n17466), .I1(encoder1_position[11]), 
            .CO(n53783));
    SB_LUT4 add_5185_10_lut (.I0(GND_net), .I1(n17467), .I2(encoder1_position[10]), 
            .I3(n53781), .O(n14989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_10 (.CI(n53781), .I0(n17467), .I1(encoder1_position[10]), 
            .CO(n53782));
    SB_LUT4 add_5185_9_lut (.I0(GND_net), .I1(n17468), .I2(encoder1_position[9]), 
            .I3(n53780), .O(n14990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_9 (.CI(n53780), .I0(n17468), .I1(encoder1_position[9]), 
            .CO(n53781));
    SB_LUT4 add_5185_8_lut (.I0(GND_net), .I1(n17469), .I2(encoder1_position[8]), 
            .I3(n53779), .O(n14991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_8 (.CI(n53779), .I0(n17469), .I1(encoder1_position[8]), 
            .CO(n53780));
    SB_LUT4 add_5185_7_lut (.I0(GND_net), .I1(n17470), .I2(encoder1_position[7]), 
            .I3(n53778), .O(n14992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_7 (.CI(n53778), .I0(n17470), .I1(encoder1_position[7]), 
            .CO(n53779));
    SB_LUT4 add_5185_6_lut (.I0(GND_net), .I1(n17471), .I2(encoder1_position[6]), 
            .I3(n53777), .O(n14993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_6 (.CI(n53777), .I0(n17471), .I1(encoder1_position[6]), 
            .CO(n53778));
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n52530), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_5_lut (.I0(GND_net), .I1(n17472), .I2(encoder1_position[5]), 
            .I3(n53776), .O(n14994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_5 (.CI(n53776), .I0(n17472), .I1(encoder1_position[5]), 
            .CO(n53777));
    SB_LUT4 add_5185_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[4]), 
            .I3(n53775), .O(n14995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_4 (.CI(n53775), .I0(encoder1_position[2]), .I1(encoder1_position[4]), 
            .CO(n53776));
    SB_LUT4 add_5185_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[3]), 
            .I3(n53774), .O(n14996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_3 (.CI(n53774), .I0(encoder1_position[1]), .I1(encoder1_position[3]), 
            .CO(n53775));
    SB_LUT4 add_5185_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n14997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n53774));
    SB_LUT4 add_5360_25_lut (.I0(GND_net), .I1(n20151), .I2(encoder1_position[26]), 
            .I3(n53767), .O(n17449)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_24_lut (.I0(GND_net), .I1(n20152), .I2(encoder1_position[25]), 
            .I3(n53766), .O(n17450)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_24 (.CI(n53766), .I0(n20152), .I1(encoder1_position[25]), 
            .CO(n53767));
    SB_LUT4 add_5360_23_lut (.I0(GND_net), .I1(n20153), .I2(encoder1_position[24]), 
            .I3(n53765), .O(n17451)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_23 (.CI(n53765), .I0(n20153), .I1(encoder1_position[24]), 
            .CO(n53766));
    SB_LUT4 add_5360_22_lut (.I0(GND_net), .I1(n20154), .I2(encoder1_position[23]), 
            .I3(n53764), .O(n17452)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_22 (.CI(n53764), .I0(n20154), .I1(encoder1_position[23]), 
            .CO(n53765));
    SB_LUT4 add_5360_21_lut (.I0(GND_net), .I1(n20155), .I2(encoder1_position[22]), 
            .I3(n53763), .O(n17453)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_21 (.CI(n53763), .I0(n20155), .I1(encoder1_position[22]), 
            .CO(n53764));
    SB_LUT4 add_5360_20_lut (.I0(GND_net), .I1(n20156), .I2(encoder1_position[21]), 
            .I3(n53762), .O(n17454)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_20 (.CI(n53762), .I0(n20156), .I1(encoder1_position[21]), 
            .CO(n53763));
    SB_LUT4 dti_counter_2039_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n53332), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n52549), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_22 (.CI(n52549), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n52550));
    SB_LUT4 dti_counter_2039_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n53331), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5360_19_lut (.I0(GND_net), .I1(n20157), .I2(encoder1_position[20]), 
            .I3(n53761), .O(n17455)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_19 (.CI(n53761), .I0(n20157), .I1(encoder1_position[20]), 
            .CO(n53762));
    SB_LUT4 add_5360_18_lut (.I0(GND_net), .I1(n20158), .I2(encoder1_position[19]), 
            .I3(n53760), .O(n17456)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_8 (.CI(n53331), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n53332));
    SB_LUT4 dti_counter_2039_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n53330), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_18 (.CI(n53760), .I0(n20158), .I1(encoder1_position[19]), 
            .CO(n53761));
    SB_LUT4 add_5360_17_lut (.I0(GND_net), .I1(n20159), .I2(encoder1_position[18]), 
            .I3(n53759), .O(n17457)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_7 (.CI(n53330), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n53331));
    SB_LUT4 dti_counter_2039_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n53329), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n52535), .O(n1245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_6 (.CI(n53329), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n53330));
    SB_CARRY add_5360_17 (.CI(n53759), .I0(n20159), .I1(encoder1_position[18]), 
            .CO(n53760));
    SB_LUT4 add_5360_16_lut (.I0(GND_net), .I1(n20160), .I2(encoder1_position[17]), 
            .I3(n53758), .O(n17458)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2039_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n53328), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_16 (.CI(n53758), .I0(n20160), .I1(encoder1_position[17]), 
            .CO(n53759));
    SB_CARRY dti_counter_2039_add_4_5 (.CI(n53328), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n53329));
    SB_LUT4 add_5360_15_lut (.I0(GND_net), .I1(n20161), .I2(encoder1_position[16]), 
            .I3(n53757), .O(n17459)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_15 (.CI(n53757), .I0(n20161), .I1(encoder1_position[16]), 
            .CO(n53758));
    SB_LUT4 dti_counter_2039_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n53327), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_4 (.CI(n53327), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n53328));
    SB_LUT4 add_5360_14_lut (.I0(GND_net), .I1(n20162), .I2(encoder1_position[15]), 
            .I3(n53756), .O(n17460)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_14 (.CI(n53756), .I0(n20162), .I1(encoder1_position[15]), 
            .CO(n53757));
    SB_LUT4 dti_counter_2039_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n53326), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_3 (.CI(n53326), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n53327));
    SB_LUT4 add_5360_13_lut (.I0(GND_net), .I1(n20163), .I2(encoder1_position[14]), 
            .I3(n53755), .O(n17461)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_13 (.CI(n53755), .I0(n20163), .I1(encoder1_position[14]), 
            .CO(n53756));
    SB_LUT4 dti_counter_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45_adj_5822)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n53326));
    SB_LUT4 add_5360_12_lut (.I0(GND_net), .I1(n20164), .I2(encoder1_position[13]), 
            .I3(n53754), .O(n17462)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_12 (.CI(n53754), .I0(n20164), .I1(encoder1_position[13]), 
            .CO(n53755));
    SB_LUT4 add_5360_11_lut (.I0(GND_net), .I1(n20165), .I2(encoder1_position[12]), 
            .I3(n53753), .O(n17463)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_11 (.CI(n53753), .I0(n20165), .I1(encoder1_position[12]), 
            .CO(n53754));
    SB_LUT4 add_5360_10_lut (.I0(GND_net), .I1(n20166), .I2(encoder1_position[11]), 
            .I3(n53752), .O(n17464)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_10 (.CI(n53752), .I0(n20166), .I1(encoder1_position[11]), 
            .CO(n53753));
    SB_LUT4 add_5360_9_lut (.I0(GND_net), .I1(n20167), .I2(encoder1_position[10]), 
            .I3(n53751), .O(n17465)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_9 (.CI(n53751), .I0(n20167), .I1(encoder1_position[10]), 
            .CO(n53752));
    SB_LUT4 add_5360_8_lut (.I0(GND_net), .I1(n20168), .I2(encoder1_position[9]), 
            .I3(n53750), .O(n17466)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_8 (.CI(n53750), .I0(n20168), .I1(encoder1_position[9]), 
            .CO(n53751));
    SB_LUT4 add_5360_7_lut (.I0(GND_net), .I1(n20169), .I2(encoder1_position[8]), 
            .I3(n53749), .O(n17467)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_7 (.CI(n53749), .I0(n20169), .I1(encoder1_position[8]), 
            .CO(n53750));
    SB_LUT4 add_5360_6_lut (.I0(GND_net), .I1(n20170), .I2(encoder1_position[7]), 
            .I3(n53748), .O(n17468)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_6 (.CI(n53748), .I0(n20170), .I1(encoder1_position[7]), 
            .CO(n53749));
    SB_LUT4 add_5360_5_lut (.I0(GND_net), .I1(n20171), .I2(encoder1_position[6]), 
            .I3(n53747), .O(n17469)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_5 (.CI(n53747), .I0(n20171), .I1(encoder1_position[6]), 
            .CO(n53748));
    SB_LUT4 add_5360_4_lut (.I0(GND_net), .I1(n20172), .I2(encoder1_position[5]), 
            .I3(n53746), .O(n17470)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_4 (.CI(n53746), .I0(n20172), .I1(encoder1_position[5]), 
            .CO(n53747));
    SB_LUT4 add_5360_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[4]), 
            .I3(n53745), .O(n17471)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_3 (.CI(n53745), .I0(encoder1_position[1]), .I1(encoder1_position[4]), 
            .CO(n53746));
    SB_LUT4 add_5360_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[3]), 
            .I3(GND_net), .O(n17472)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5360_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5360_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[3]), 
            .CO(n53745));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n52548), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_21 (.CI(n52548), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n52549));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n52547), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_3 (.CI(n52530), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n52531));
    SB_CARRY add_151_8 (.CI(n52535), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n52536));
    SB_CARRY add_151_20 (.CI(n52547), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n52548));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n52546), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n52788), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n52787), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n52787), .I0(GND_net), .I1(n2), 
            .CO(n52788));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5704), 
            .I3(n52786), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5393_23_lut (.I0(GND_net), .I1(n21357), .I2(encoder1_position[23]), 
            .I3(n53717), .O(n20151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5393_22_lut (.I0(GND_net), .I1(n21358), .I2(encoder1_position[22]), 
            .I3(n53716), .O(n20152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_22 (.CI(n53716), .I0(n21358), .I1(encoder1_position[22]), 
            .CO(n53717));
    SB_LUT4 add_5393_21_lut (.I0(GND_net), .I1(n21359), .I2(encoder1_position[21]), 
            .I3(n53715), .O(n20153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_21 (.CI(n53715), .I0(n21359), .I1(encoder1_position[21]), 
            .CO(n53716));
    SB_LUT4 add_5393_20_lut (.I0(GND_net), .I1(n21360), .I2(encoder1_position[20]), 
            .I3(n53714), .O(n20154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_20 (.CI(n53714), .I0(n21360), .I1(encoder1_position[20]), 
            .CO(n53715));
    SB_LUT4 add_5393_19_lut (.I0(GND_net), .I1(n21361), .I2(encoder1_position[19]), 
            .I3(n53713), .O(n20155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_19 (.CI(n53713), .I0(n21361), .I1(encoder1_position[19]), 
            .CO(n53714));
    SB_LUT4 add_5393_18_lut (.I0(GND_net), .I1(n21362), .I2(encoder1_position[18]), 
            .I3(n53712), .O(n20156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_18 (.CI(n53712), .I0(n21362), .I1(encoder1_position[18]), 
            .CO(n53713));
    SB_LUT4 add_5393_17_lut (.I0(GND_net), .I1(n21363), .I2(encoder1_position[17]), 
            .I3(n53711), .O(n20157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_17 (.CI(n53711), .I0(n21363), .I1(encoder1_position[17]), 
            .CO(n53712));
    SB_LUT4 add_5393_16_lut (.I0(GND_net), .I1(n21364), .I2(encoder1_position[16]), 
            .I3(n53710), .O(n20158)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_16 (.CI(n53710), .I0(n21364), .I1(encoder1_position[16]), 
            .CO(n53711));
    SB_LUT4 add_5393_15_lut (.I0(GND_net), .I1(n21365), .I2(encoder1_position[15]), 
            .I3(n53709), .O(n20159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_15 (.CI(n53709), .I0(n21365), .I1(encoder1_position[15]), 
            .CO(n53710));
    SB_LUT4 add_5393_14_lut (.I0(GND_net), .I1(n21366), .I2(encoder1_position[14]), 
            .I3(n53708), .O(n20160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n52786), .I0(GND_net), .I1(n14_adj_5704), 
            .CO(n52787));
    SB_CARRY add_5393_14 (.CI(n53708), .I0(n21366), .I1(encoder1_position[14]), 
            .CO(n53709));
    SB_LUT4 add_5393_13_lut (.I0(GND_net), .I1(n21367), .I2(encoder1_position[13]), 
            .I3(n53707), .O(n20161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_13 (.CI(n53707), .I0(n21367), .I1(encoder1_position[13]), 
            .CO(n53708));
    SB_LUT4 add_5393_12_lut (.I0(GND_net), .I1(n21368), .I2(encoder1_position[12]), 
            .I3(n53706), .O(n20162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_12 (.CI(n53706), .I0(n21368), .I1(encoder1_position[12]), 
            .CO(n53707));
    SB_LUT4 add_5393_11_lut (.I0(GND_net), .I1(n21369), .I2(encoder1_position[11]), 
            .I3(n53705), .O(n20163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_11 (.CI(n53705), .I0(n21369), .I1(encoder1_position[11]), 
            .CO(n53706));
    SB_LUT4 add_5393_10_lut (.I0(GND_net), .I1(n21370), .I2(encoder1_position[10]), 
            .I3(n53704), .O(n20164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_10 (.CI(n53704), .I0(n21370), .I1(encoder1_position[10]), 
            .CO(n53705));
    SB_LUT4 add_5393_9_lut (.I0(GND_net), .I1(n21371), .I2(encoder1_position[9]), 
            .I3(n53703), .O(n20165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_9 (.CI(n53703), .I0(n21371), .I1(encoder1_position[9]), 
            .CO(n53704));
    SB_LUT4 add_5393_8_lut (.I0(GND_net), .I1(n21372), .I2(encoder1_position[8]), 
            .I3(n53702), .O(n20166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_8 (.CI(n53702), .I0(n21372), .I1(encoder1_position[8]), 
            .CO(n53703));
    SB_LUT4 add_5393_7_lut (.I0(GND_net), .I1(n21373), .I2(encoder1_position[7]), 
            .I3(n53701), .O(n20167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_7 (.CI(n53701), .I0(n21373), .I1(encoder1_position[7]), 
            .CO(n53702));
    SB_LUT4 add_5393_6_lut (.I0(GND_net), .I1(n21374), .I2(encoder1_position[6]), 
            .I3(n53700), .O(n20168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_6 (.CI(n53700), .I0(n21374), .I1(encoder1_position[6]), 
            .CO(n53701));
    SB_LUT4 add_5393_5_lut (.I0(GND_net), .I1(n21375), .I2(encoder1_position[5]), 
            .I3(n53699), .O(n20169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_5 (.CI(n53699), .I0(n21375), .I1(encoder1_position[5]), 
            .CO(n53700));
    SB_LUT4 add_5393_4_lut (.I0(GND_net), .I1(n21376), .I2(encoder1_position[4]), 
            .I3(n53698), .O(n20170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_4 (.CI(n53698), .I0(n21376), .I1(encoder1_position[4]), 
            .CO(n53699));
    SB_LUT4 add_5393_3_lut (.I0(GND_net), .I1(n21377), .I2(encoder1_position[3]), 
            .I3(n53697), .O(n20171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_3 (.CI(n53697), .I0(n21377), .I1(encoder1_position[3]), 
            .CO(n53698));
    SB_LUT4 add_5393_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n20172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5393_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5393_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n53697));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5705), 
            .I3(n52785), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n52785), .I0(GND_net), .I1(n15_adj_5705), 
            .CO(n52786));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5706), 
            .I3(n52784), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n52784), .I0(GND_net), .I1(n16_adj_5706), 
            .CO(n52785));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5707), 
            .I3(n52783), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n52783), .I0(GND_net), .I1(n17_adj_5707), 
            .CO(n52784));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5708), 
            .I3(n52782), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n52782), .I0(GND_net), .I1(n18_adj_5708), 
            .CO(n52783));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5709), 
            .I3(n52781), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n52781), .I0(GND_net), .I1(n19_adj_5709), 
            .CO(n52782));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5710), 
            .I3(n52780), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n52780), .I0(GND_net), .I1(n20_adj_5710), 
            .CO(n52781));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5711), 
            .I3(n52779), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n52779), .I0(GND_net), .I1(n21_adj_5711), 
            .CO(n52780));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5712), 
            .I3(n52778), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n52778), .I0(GND_net), .I1(n22_adj_5712), 
            .CO(n52779));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5713), 
            .I3(n52777), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n52777), .I0(GND_net), .I1(n23_adj_5713), 
            .CO(n52778));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5714), 
            .I3(n52776), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n52776), .I0(GND_net), .I1(n24_adj_5714), 
            .CO(n52777));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n41880), .I1(GND_net), .I2(n25_adj_5715), 
            .I3(VCC_net), .O(n67594)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5715), 
            .CO(n52776));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n52534), .O(n1246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_19 (.CI(n52546), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n52547));
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n52545), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_18 (.CI(n52545), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n52546));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n52544), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n52544), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n52545));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5777), .I3(n52706), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3), .I3(n52705), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n52705), .I0(encoder0_position_scaled[22]), 
            .I1(n3), .CO(n52706));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5776), .I3(n52704), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n52704), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5776), .CO(n52705));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n52543), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5793), .I3(n52703), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n52703), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5793), .CO(n52704));
    SB_CARRY add_151_7 (.CI(n52534), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n52535));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5792), .I3(n52702), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n52702), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5792), .CO(n52703));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5791), .I3(n52701), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_16 (.CI(n52543), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n52544));
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n52530));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n52701), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5791), .CO(n52702));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5790), .I3(n52700), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n52533), .O(n1247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n52542), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_6 (.CI(n52533), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n52534));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n52700), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5790), .CO(n52701));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5789), .I3(n52699), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n52542), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n52543));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n52699), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5789), .CO(n52700));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n52541), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5775), .I3(n52698), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n52698), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5775), .CO(n52699));
    SB_LUT4 i12_2_lut (.I0(pwm_setpoint[6]), .I1(pwm_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5772));   // verilog/pwm.v(11[19:30])
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5774), .I3(n52697), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n52697), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5774), .CO(n52698));
    SB_LUT4 i13742_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3180), .I3(GND_net), 
            .O(n31687));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5773), .I3(n52696), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n52696), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5773), .CO(n52697));
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n23_adj_5843), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5232), .I3(o_Rx_DV_N_3488[8]), .O(n63043));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63043), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5771));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n59686), .O(n63193));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63193), .O(n63199));
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63453), .O(n63459));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63459), .O(n63465));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 i14000_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n63465), 
            .I3(n27), .O(n31945));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14000_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14724_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n32669));   // verilog/coms.v(130[12] 305[6])
    defparam i14724_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23520_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i23520_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23519_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i23519_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1801 (.I0(\data_out_frame[18] [6]), .I1(n28303), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5850));
    defparam i1_2_lut_adj_1801.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n55561), .I1(n28021), .I2(n60355), .I3(n6_adj_5850), 
            .O(n54982));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23649_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i23649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_1180_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5821));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1180_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45344_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64614));
    defparam i45344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i8_4_lut (.I0(displacement[7]), .I1(encoder0_position_scaled[7]), 
            .I2(n54181), .I3(n51206), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i45345_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64615));
    defparam i45345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45621_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64891));
    defparam i45621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45620_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64890));
    defparam i45620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13810_4_lut_4_lut (.I0(n29957), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n31755));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13810_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 mux_245_i9_4_lut (.I0(displacement[8]), .I1(encoder0_position_scaled[8]), 
            .I2(n54181), .I3(n51206), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(bit_ctr[3]), .I2(n41559), 
            .I3(bit_ctr[4]), .O(n4));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hd555;
    SB_LUT4 i14002_3_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(n62228), .I3(GND_net), .O(n31947));   // verilog/coms.v(130[12] 305[6])
    defparam i14002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48687_2_lut (.I0(n71521), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67759));
    defparam i48687_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5773));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5774));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5775));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5789));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5790));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5791));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5792));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5793));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i12_4_lut (.I0(displacement[11]), .I1(encoder0_position_scaled[11]), 
            .I2(n54181), .I3(n51206), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5776));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i13_4_lut (.I0(displacement[12]), .I1(encoder0_position_scaled[12]), 
            .I2(n54181), .I3(n51206), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i14_4_lut (.I0(displacement[13]), .I1(encoder0_position_scaled[13]), 
            .I2(n54181), .I3(n51206), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5777));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1802 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n63559));
    defparam i1_2_lut_adj_1802.LUT_INIT = 16'heeee;
    SB_LUT4 mux_245_i15_4_lut (.I0(displacement[14]), .I1(encoder0_position_scaled[14]), 
            .I2(n54181), .I3(n51206), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(r_SM_Main[1]), .I1(n6_adj_5846), .I2(r_Bit_Index[0]), 
            .I3(n63559), .O(n63545));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hffdf;
    SB_LUT4 mux_245_i16_4_lut (.I0(displacement[15]), .I1(encoder0_position_scaled[15]), 
            .I2(n54181), .I3(n51206), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 mux_245_i17_4_lut (.I0(displacement[16]), .I1(encoder0_position_scaled[16]), 
            .I2(n54181), .I3(n51206), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63545), .O(n63551));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i18_4_lut (.I0(displacement[17]), .I1(encoder0_position_scaled[17]), 
            .I2(n54181), .I3(n51206), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63551), .O(n63557));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i19_4_lut (.I0(displacement[18]), .I1(encoder0_position_scaled[18]), 
            .I2(n54181), .I3(n51206), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 mux_245_i20_4_lut (.I0(displacement[19]), .I1(encoder0_position_scaled[19]), 
            .I2(n54181), .I3(n51206), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(n3491), .I3(n10_adj_5717), .O(n60044));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 mux_245_i21_4_lut (.I0(displacement[20]), .I1(encoder0_position_scaled[20]), 
            .I2(n54181), .I3(n51206), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 mux_245_i22_4_lut (.I0(displacement[21]), .I1(encoder0_position_scaled[21]), 
            .I2(n54181), .I3(n51206), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i13757_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n63557), 
            .I3(n27), .O(n31702));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13757_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_245_i23_4_lut (.I0(displacement[22]), .I1(encoder0_position_scaled[22]), 
            .I2(n54181), .I3(n51206), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 mux_245_i24_4_lut (.I0(displacement[23]), .I1(encoder0_position_scaled[23]), 
            .I2(n54181), .I3(n51206), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'hf353;
    SB_LUT4 i1957_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1331), .I3(n41376), .O(n6917));   // verilog/TinyFPGA_B.v(363[5] 389[12])
    defparam i1957_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5711));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5710));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5709));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5708));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5707));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5706));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5705));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5704));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[1]), .I3(neopxl_color[3]), .O(n71422));
    defparam color_bit_N_502_1__bdd_4_lut_4_lut.LUT_INIT = 16'he6a2;
    SB_LUT4 i45609_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64879));
    defparam i45609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45610_4_lut (.I0(n64879), .I1(n30156), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1] [5]), .O(n64880));
    defparam i45610_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i45608_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64878));
    defparam i45608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1806 (.I0(\data_out_frame[18] [7]), .I1(n61989), 
            .I2(GND_net), .I3(GND_net), .O(n60355));
    defparam i1_2_lut_adj_1806.LUT_INIT = 16'h9999;
    SB_LUT4 i13647_3_lut_4_lut (.I0(n1755), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n31592));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13647_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i13645_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n31590));   // verilog/coms.v(130[12] 305[6])
    defparam i13645_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13634_3_lut_4_lut (.I0(n1805), .I1(b_prev_adj_5768), .I2(a_new_adj_5891[1]), 
            .I3(position_31__N_3836_adj_5770), .O(n31579));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13634_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i5558_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5558_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i5556_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5556_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i51672_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n41376), .I3(GND_net), .O(n29830));
    defparam i51672_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i5560_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i5560_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i49476_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n67643));
    defparam i49476_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i23634_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n41376), .I3(GND_net), .O(n41480));
    defparam i23634_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i5562_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i5562_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63435), .O(n63441));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63441), .O(n63447));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i14016_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n63447), 
            .I3(n27), .O(n31961));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14016_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13535_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5927[1]), 
            .I2(r_SM_Main_adj_5927[2]), .I3(n6_adj_5825), .O(n31480));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13535_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i13491_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n29776), .I3(GND_net), .O(n31436));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n59826));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n59825));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n59824));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63507), .O(n63513));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63513), .O(n63519));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i14075_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n63519), 
            .I3(n27), .O(n32020));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14075_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n59823));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n31262));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n59770));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63471), .O(n63477));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63477), .O(n63483));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i14076_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n63483), 
            .I3(n27), .O(n32021));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14076_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1818 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n59822));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1818.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1819 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n59821));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1819.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1820 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n59820));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1820.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n31257));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n59819));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n59818));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n59817));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h2300;
    SB_LUT4 i14554_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2889));   // verilog/coms.v(130[12] 305[6])
    defparam i14554_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n59816));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n59946));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n59945));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n59944));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n59815));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n59943));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n59942));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n59941));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n31251));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h2300;
    SB_LUT4 i49300_3_lut (.I0(enable_slow_N_4213), .I1(n41430), .I2(state_7__N_4110[0]), 
            .I3(GND_net), .O(n67768));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i49300_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_5937[0]), .I1(n67768), .I2(n6722), 
            .I3(n6_adj_5830), .O(n8_adj_5847));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n59947));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h2300;
    SB_LUT4 i14120_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[0]), 
            .I2(n10_adj_5824), .I3(n27672), .O(n32065));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n59814));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1836 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n59813));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1836.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n6_adj_5846), .I1(r_SM_Main[1]), .I2(n63559), 
            .I3(r_Bit_Index[0]), .O(n63565));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63565), .O(n63571));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1839 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63571), .O(n63577));
    defparam i1_4_lut_adj_1839.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n59812));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 i14142_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n63577), 
            .I3(n27), .O(n32087));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14142_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n59811));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1842 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n59810));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1842.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n59809));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n59808));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_adj_1845 (.I0(n15_adj_5760), .I1(n25001), .I2(dti), 
            .I3(GND_net), .O(n29728));
    defparam i1_2_lut_3_lut_adj_1845.LUT_INIT = 16'hbaba;
    SB_LUT4 i14156_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[0]), .I2(n11_adj_5779), 
            .I3(state_7__N_4319), .O(n32101));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14156_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n59807));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n59806));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n59805));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n59804));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1679_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n10012));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1850 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n59940));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1850.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1851 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n59939));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1851.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1852 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n59803));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1852.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1679_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n11494));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1853 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n31237));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1853.LUT_INIT = 16'h2300;
    SB_LUT4 i13558_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n30416), 
            .I3(GND_net), .O(n31503));   // verilog/coms.v(130[12] 305[6])
    defparam i13558_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13555_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n30416), 
            .I3(GND_net), .O(n31500));   // verilog/coms.v(130[12] 305[6])
    defparam i13555_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1679_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n11492));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1854 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n59802));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1854.LUT_INIT = 16'h2300;
    SB_LUT4 i13546_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n30416), 
            .I3(GND_net), .O(n31491));   // verilog/coms.v(130[12] 305[6])
    defparam i13546_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n59938));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n59937));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n59936));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n59935));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1859 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n59934));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1859.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1860 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n59933));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1860.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1861 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n59932));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1861.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1862 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n59931));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1862.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1863 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n59930));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1863.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1864 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n59929));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1864.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n59928));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n59927));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1867 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n59926));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1867.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n59925));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h2300;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n29817), .O(n55814));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n59924));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n59801));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n59800));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n59799));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n59798));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1874 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n59797));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1874.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n59796));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n59923));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n59795));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h2300;
    SB_LUT4 i19277_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n24903), .I3(GND_net), .O(n32185));
    defparam i19277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n59922));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h2300;
    SB_LUT4 i14241_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n24903), .I3(GND_net), .O(n32186));   // verilog/coms.v(130[12] 305[6])
    defparam i14241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14242_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n24903), .I3(GND_net), .O(n32187));   // verilog/coms.v(130[12] 305[6])
    defparam i14242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14243_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n24903), .I3(GND_net), .O(n32188));   // verilog/coms.v(130[12] 305[6])
    defparam i14243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14244_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n24903), .I3(GND_net), .O(n32189));   // verilog/coms.v(130[12] 305[6])
    defparam i14244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14245_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n24903), .I3(GND_net), .O(n32190));   // verilog/coms.v(130[12] 305[6])
    defparam i14245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14246_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n24903), .I3(GND_net), .O(n32191));   // verilog/coms.v(130[12] 305[6])
    defparam i14246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14247_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n24903), .I3(GND_net), .O(n32192));   // verilog/coms.v(130[12] 305[6])
    defparam i14247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5839));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i6917_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n24553));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i6917_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_adj_1879 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1331), .I3(n41376), .O(n24_adj_5835));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_adj_1879.LUT_INIT = 16'hffbf;
    SB_LUT4 i14248_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n24903), .I3(GND_net), .O(n32193));   // verilog/coms.v(130[12] 305[6])
    defparam i14248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14250_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n24903), .I3(GND_net), .O(n32195));   // verilog/coms.v(130[12] 305[6])
    defparam i14250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6174_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i6174_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14251_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n24903), .I3(GND_net), .O(n32196));   // verilog/coms.v(130[12] 305[6])
    defparam i14251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14252_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n24903), .I3(GND_net), .O(n32197));   // verilog/coms.v(130[12] 305[6])
    defparam i14252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14254_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n24903), .I3(GND_net), .O(n32199));   // verilog/coms.v(130[12] 305[6])
    defparam i14254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14255_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n24903), .I3(GND_net), .O(n32200));   // verilog/coms.v(130[12] 305[6])
    defparam i14255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13963_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n24553), .I3(n4_adj_5851), .O(n31908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i13963_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i14256_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n24903), .I3(GND_net), .O(n32201));   // verilog/coms.v(130[12] 305[6])
    defparam i14256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n59794));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i14257_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n24903), .I3(GND_net), .O(n32202));   // verilog/coms.v(130[12] 305[6])
    defparam i14257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14258_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n24903), .I3(GND_net), .O(n32203));   // verilog/coms.v(130[12] 305[6])
    defparam i14258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n59793));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n59921));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_LUT4 i18556_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n24877), .I3(GND_net), .O(n31462));
    defparam i18556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n59792));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 i13518_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n24903), .I3(GND_net), .O(n31463));   // verilog/coms.v(130[12] 305[6])
    defparam i13518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1679_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n11490));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n59791));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n59920));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n59790));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 i14261_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n24903), .I3(GND_net), .O(n32206));   // verilog/coms.v(130[12] 305[6])
    defparam i14261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18682_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n24877), .I3(GND_net), .O(n32207));
    defparam i18682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n59789));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 i14263_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n24877), .I3(GND_net), .O(n32208));   // verilog/coms.v(130[12] 305[6])
    defparam i14263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18704_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n24877), .I3(GND_net), .O(n32209));
    defparam i18704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18711_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n24877), .I3(GND_net), .O(n32210));
    defparam i18711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14266_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n24877), .I3(GND_net), .O(n32211));   // verilog/coms.v(130[12] 305[6])
    defparam i14266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14267_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n24877), .I3(GND_net), .O(n32212));   // verilog/coms.v(130[12] 305[6])
    defparam i14267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14268_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n24877), .I3(GND_net), .O(n32213));   // verilog/coms.v(130[12] 305[6])
    defparam i14268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14269_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n24877), .I3(GND_net), .O(n32214));   // verilog/coms.v(130[12] 305[6])
    defparam i14269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14270_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n24877), .I3(GND_net), .O(n32215));   // verilog/coms.v(130[12] 305[6])
    defparam i14270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13788_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n60042), 
            .I3(GND_net), .O(n31733));   // verilog/coms.v(130[12] 305[6])
    defparam i13788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14271_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n24877), .I3(GND_net), .O(n32216));   // verilog/coms.v(130[12] 305[6])
    defparam i14271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14272_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n24877), .I3(GND_net), .O(n32217));   // verilog/coms.v(130[12] 305[6])
    defparam i14272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14273_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n24877), .I3(GND_net), .O(n32218));   // verilog/coms.v(130[12] 305[6])
    defparam i14273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18636_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n24877), .I3(GND_net), .O(n32220));
    defparam i18636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18660_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n24877), .I3(GND_net), .O(n32221));
    defparam i18660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14277_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n24877), .I3(GND_net), .O(n32222));   // verilog/coms.v(130[12] 305[6])
    defparam i14277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n59788));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_LUT4 i13791_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n60042), 
            .I3(GND_net), .O(n31736));   // verilog/coms.v(130[12] 305[6])
    defparam i13791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14280_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n24877), .I3(GND_net), .O(n32225));   // verilog/coms.v(130[12] 305[6])
    defparam i14280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14281_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n24877), .I3(GND_net), .O(n32226));   // verilog/coms.v(130[12] 305[6])
    defparam i14281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n23_adj_5843), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5235), .I3(r_SM_Main_adj_5927[0]), .O(n63595));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfeff;
    SB_LUT4 i18510_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n24877), .I3(GND_net), .O(n32227));
    defparam i18510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18515_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n24877), .I3(GND_net), .O(n32228));
    defparam i18515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18516_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n24877), .I3(GND_net), .O(n32229));
    defparam i18516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13543_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n30416), 
            .I3(GND_net), .O(n31488));   // verilog/coms.v(130[12] 305[6])
    defparam i13543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n59787));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n59786));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63595), .O(n61652));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n59785));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63525), .O(n63531));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63531), .O(n63537));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 i14286_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n63537), 
            .I3(n27), .O(n32231));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14286_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n59784));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n59919));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n59783));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n59782));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n59781));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n59780));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n59779));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n59778));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n59777));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n59918));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n59776));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n59775));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n59774));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n41376), .O(n58154));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n59773));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n59772));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n59771));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n59832));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n59917));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n59916));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n59915));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n59914));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1917 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n59913));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1917.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n59912));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n59911));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n59910));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n59909));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n59908));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n59907));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n59906));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n59905));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n59904));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n59833));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n59903));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n59902));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n59901));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1931 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n59900));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1931.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n59899));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n59898));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n59897));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n59896));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n59895));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n59894));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n59893));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n59892));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n59891));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1941 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n59890));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1941.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1942 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n59889));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1942.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n59888));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n59887));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n59886));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n59885));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n59884));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n59883));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n59882));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n59881));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n59880));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n59879));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i14363_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n29776), .I3(GND_net), .O(n32308));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n59878));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 i13537_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n30416), 
            .I3(GND_net), .O(n31482));   // verilog/coms.v(130[12] 305[6])
    defparam i13537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n31321));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n59877));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 i14366_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n29776), .I3(GND_net), .O(n32311));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14367_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n338), 
            .I2(n29776), .I3(GND_net), .O(n32312));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14368_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n29776), .I3(GND_net), .O(n32313));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14369_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n29776), .I3(GND_net), .O(n32314));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n59876));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i14370_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n341), 
            .I2(n29776), .I3(GND_net), .O(n32315));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14371_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n29776), .I3(GND_net), .O(n32316));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14372_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n29776), .I3(GND_net), .O(n32317));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14373_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n29776), .I3(GND_net), .O(n32318));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n59875));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n59874));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n59873));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_LUT4 i14374_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n29776), .I3(GND_net), .O(n32319));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14375_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n29776), .I3(GND_net), .O(n32320));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n59872));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 i14376_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n29776), .I3(GND_net), .O(n32321));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14377_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n29776), .I3(GND_net), .O(n32322));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14378_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n29776), .I3(GND_net), .O(n32323));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14379_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n29776), .I3(GND_net), .O(n32324));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14380_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n29776), .I3(GND_net), .O(n32325));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14381_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n29776), .I3(GND_net), .O(n32326));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14382_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n29776), .I3(GND_net), .O(n32327));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14383_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n29776), .I3(GND_net), .O(n32328));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13982_3_lut (.I0(\data_in_frame[16] [0]), .I1(rx_data[0]), 
            .I2(n62228), .I3(GND_net), .O(n31927));   // verilog/coms.v(130[12] 305[6])
    defparam i13982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14384_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n29776), .I3(GND_net), .O(n32329));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14385_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n29776), .I3(GND_net), .O(n32330));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n59871));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i14386_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n29776), .I3(GND_net), .O(n32331));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n59870));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i14387_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n29776), .I3(GND_net), .O(n32332));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main_adj_5927[0]), .I1(o_Rx_DV_N_3488[24]), 
            .I2(n27), .I3(GND_net), .O(n14_adj_5832));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(o_Rx_DV_N_3488[12]), .I2(n23_adj_5843), 
            .I3(n5235), .O(n15_adj_5831));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5831), .I1(n1), .I2(n14_adj_5832), .I3(r_SM_Main_adj_5927[1]), 
            .O(n71705));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i14390_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[1]), 
            .I2(n10_adj_5824), .I3(n27624), .O(n32335));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14390_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14392_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[2]), 
            .I2(n4_adj_5761), .I3(n27672), .O(n32337));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14392_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14393_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[3]), 
            .I2(n4_adj_5761), .I3(n27624), .O(n32338));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14393_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14394_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[4]), 
            .I2(n4_adj_5762), .I3(n27672), .O(n32339));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14394_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n59869));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i49346_4_lut (.I0(data_ready), .I1(n6917), .I2(n24_adj_5835), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n67734));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i49346_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i49359_2_lut (.I0(n24_adj_5835), .I1(n6917), .I2(GND_net), 
            .I3(GND_net), .O(n67737));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i49359_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n67737), .I1(n67734), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5839), .O(n58068));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n59868));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n59867));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n59866));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n59865));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i13985_3_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n62228), .I3(GND_net), .O(n31930));   // verilog/coms.v(130[12] 305[6])
    defparam i13985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n59864));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n59863));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n59862));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n59861));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n59860));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n59859));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n59834));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n59858));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n31299));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i14411_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[5]), 
            .I2(n4_adj_5762), .I3(n27624), .O(n32356));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14411_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n59857));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n59856));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n59855));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n59854));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i14415_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[6]), 
            .I2(n41590), .I3(n27672), .O(n32360));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14415_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n31294));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n59853));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n59852));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 i14417_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5904[7]), 
            .I2(n41590), .I3(n27624), .O(n32362));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14417_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14147_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n30452), .I3(GND_net), .O(n32092));   // verilog/coms.v(130[12] 305[6])
    defparam i14147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13510_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n30414), 
            .I3(GND_net), .O(n31455));   // verilog/coms.v(130[12] 305[6])
    defparam i13510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14143_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n30452), .I3(GND_net), .O(n32088));   // verilog/coms.v(130[12] 305[6])
    defparam i14143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n59851));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i14138_4_lut (.I0(n63175), .I1(r_Bit_Index[0]), .I2(n60834), 
            .I3(n29821), .O(n32083));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14138_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i13507_3_lut (.I0(\data_in_frame[2] [4]), .I1(rx_data[4]), .I2(n30414), 
            .I3(GND_net), .O(n31452));   // verilog/coms.v(130[12] 305[6])
    defparam i13507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14133_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n30452), .I3(GND_net), .O(n32078));   // verilog/coms.v(130[12] 305[6])
    defparam i14133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14129_4_lut (.I0(n63177), .I1(r_Bit_Index_adj_5929[0]), .I2(n60832), 
            .I3(n29824), .O(n32074));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i14129_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i13504_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n30414), 
            .I3(GND_net), .O(n31449));   // verilog/coms.v(130[12] 305[6])
    defparam i13504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13501_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n30414), 
            .I3(GND_net), .O(n31446));   // verilog/coms.v(130[12] 305[6])
    defparam i13501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n59850));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 i14121_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n30452), .I3(GND_net), .O(n32066));   // verilog/coms.v(130[12] 305[6])
    defparam i14121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n59849));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n59848));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n59847));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n59846));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n59845));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5722));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14439_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[1]), .I2(n5_adj_5778), 
            .I3(n27680), .O(n32384));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14439_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14440_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[2]), .I2(n5_adj_5806), 
            .I3(n27680), .O(n32385));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14440_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6_4_lut_adj_1991 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5721));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_1991.LUT_INIT = 16'hfffe;
    SB_LUT4 i14441_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[3]), .I2(n41527), 
            .I3(n27680), .O(n32386));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14441_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14442_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[4]), .I2(n9_adj_5780), 
            .I3(n27667), .O(n32387));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14442_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14443_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[5]), .I2(n5_adj_5778), 
            .I3(n27667), .O(n32388));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14443_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14444_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[6]), .I2(n5_adj_5806), 
            .I3(n27667), .O(n32389));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14444_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n31284));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n59844));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i14445_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[7]), .I2(n41527), 
            .I3(n27667), .O(n32390));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14445_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14446_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[8]), .I2(n9_adj_5780), 
            .I3(n27643), .O(n32391));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14446_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14447_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[9]), .I2(n5_adj_5778), 
            .I3(n27643), .O(n32392));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14447_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14448_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[10]), .I2(n5_adj_5806), 
            .I3(n27643), .O(n32393));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14448_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n59843));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i7_4_lut_adj_1995 (.I0(dti_counter[0]), .I1(n14_adj_5721), .I2(n10_adj_5722), 
            .I3(dti_counter[3]), .O(n25001));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_1995.LUT_INIT = 16'hfffe;
    SB_LUT4 i14449_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[11]), .I2(n41527), 
            .I3(n27643), .O(n32394));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14449_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14450_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[12]), .I2(n9_adj_5780), 
            .I3(n27661), .O(n32395));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14450_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n59842));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n59841));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1998 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5718));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1998.LUT_INIT = 16'h7bde;
    SB_LUT4 i14451_4_lut (.I0(CS_MISO_c), .I1(data_adj_5911[15]), .I2(n41527), 
            .I3(n27661), .O(n32396));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14451_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n59840));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n59839));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n31277));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n59838));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i13988_3_lut (.I0(\data_in_frame[16] [2]), .I1(rx_data[2]), 
            .I2(n62228), .I3(GND_net), .O(n31933));   // verilog/coms.v(130[12] 305[6])
    defparam i13988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_2003 (.I0(commutation_state[0]), .I1(n4_adj_5718), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5760));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut_adj_2003.LUT_INIT = 16'hdede;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n59837));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n59836));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n59835));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n59831));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n59830));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 i51861_2_lut (.I0(n25001), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i51861_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n59829));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i13498_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n30414), 
            .I3(GND_net), .O(n31443));   // verilog/coms.v(130[12] 305[6])
    defparam i13498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n31269));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n59828));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n59827));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2013 (.I0(\data_in_frame[19] [7]), .I1(n30366), 
            .I2(n30449), .I3(rx_data[7]), .O(n59136));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2013.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13495_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n30414), 
            .I3(GND_net), .O(n31440));   // verilog/coms.v(130[12] 305[6])
    defparam i13495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_2014 (.I0(\data_in_frame[19] [2]), .I1(n30366), 
            .I2(n30449), .I3(rx_data[2]), .O(n59138));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2014.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2015 (.I0(\data_in_frame[19] [0]), .I1(n30366), 
            .I2(n30449), .I3(rx_data[0]), .O(n59140));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2015.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[18] [6]), .I1(n30368), .I2(n30447), 
            .I3(rx_data[6]), .O(n59142));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14051_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n30447), .I3(GND_net), .O(n31996));   // verilog/coms.v(130[12] 305[6])
    defparam i14051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_2016 (.I0(\data_in_frame[18] [4]), .I1(n30368), 
            .I2(n30447), .I3(rx_data[4]), .O(n59144));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2016.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14045_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n30447), .I3(GND_net), .O(n31990));   // verilog/coms.v(130[12] 305[6])
    defparam i14045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2017 (.I0(\data_in_frame[18] [2]), .I1(n30368), 
            .I2(n30447), .I3(rx_data[2]), .O(n59146));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2017.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2018 (.I0(\data_in_frame[18] [1]), .I1(n30368), 
            .I2(n30447), .I3(rx_data[1]), .O(n59148));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2018.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2019 (.I0(\data_in_frame[18] [0]), .I1(n30368), 
            .I2(n30447), .I3(rx_data[0]), .O(n59150));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2019.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14032_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n62670), .I3(GND_net), .O(n31977));   // verilog/coms.v(130[12] 305[6])
    defparam i14032_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14029_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n62670), .I3(GND_net), .O(n31974));   // verilog/coms.v(130[12] 305[6])
    defparam i14029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14026_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n62670), .I3(GND_net), .O(n31971));   // verilog/coms.v(130[12] 305[6])
    defparam i14026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14023_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n62670), .I3(GND_net), .O(n31968));   // verilog/coms.v(130[12] 305[6])
    defparam i14023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14020_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n62670), .I3(GND_net), .O(n31965));   // verilog/coms.v(130[12] 305[6])
    defparam i14020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1679_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n11488));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13526_3_lut (.I0(current[0]), .I1(data_adj_5911[0]), .I2(n29799), 
            .I3(GND_net), .O(n31471));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14009_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n62670), .I3(GND_net), .O(n31954));   // verilog/coms.v(130[12] 305[6])
    defparam i14009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1679_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n11486));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13536_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3180), .I3(GND_net), 
            .O(n31481));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1679_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n11484));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n11482));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n11480));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n11478));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n11476));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_2_lut_adj_2020 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_2020.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut_adj_2021 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_2021.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_4_lut_adj_2022 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2836), .O(n25_adj_5834));   // verilog/TinyFPGA_B.v(378[7:11])
    defparam i1_4_lut_4_lut_adj_2022.LUT_INIT = 16'h5450;
    SB_LUT4 i12914_2_lut (.I0(n29752), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n30865));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i12914_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51631_4_lut (.I0(commutation_state[1]), .I1(n25001), .I2(dti), 
            .I3(commutation_state[2]), .O(n29752));
    defparam i51631_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 mux_1679_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n11474));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n11472));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i5566_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5566_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i5564_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5564_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i13794_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n60042), 
            .I3(GND_net), .O(n31739));   // verilog/coms.v(130[12] 305[6])
    defparam i13794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1679_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n11470));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13193_4_lut (.I0(n29830), .I1(n1331), .I2(n67643), .I3(n41480), 
            .O(n31109));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i13193_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1679_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n11468));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n11466));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n11464));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n11462));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i51898_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5852));
    defparam i51898_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 mux_1679_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n11460));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n11458));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n11456));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1679_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n11454));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1679_i22_3_lut.LUT_INIT = 16'h3535;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1800(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .\a_new[1] (a_new_adj_5891[1]), 
            .\b_new[1] (b_new_adj_5892[1]), .n31593(n31593), .a_prev(a_prev_adj_5767), 
            .n31582(n31582), .b_prev(b_prev_adj_5768), .n31579(n31579), 
            .n1805(n1805), .position_31__N_3836(position_31__N_3836_adj_5770), 
            .encoder1_position({encoder1_position}), .GND_net(GND_net), 
            .VCC_net(VCC_net), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5769)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i41631_3_lut (.I0(n4_adj_5851), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n60846));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i41631_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n62898));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i13637_3_lut (.I0(b_prev_adj_5768), .I1(b_new_adj_5892[1]), 
            .I2(debounce_cnt_N_3833_adj_5769), .I3(GND_net), .O(n31582));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13644_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n31589));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13646_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n31591));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13646_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1800(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .\a_new[1] (a_new[1]), 
            .\b_new[1] (b_new[1]), .n1757(n1757), .GND_net(GND_net), .n1759(n1759), 
            .n1761(n1761), .n1763(n1763), .n1765(n1765), .n1767(n1767), 
            .n1769(n1769), .n1771(n1771), .n1773(n1773), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .n31592(n31592), 
            .n1755(n1755), .n31591(n31591), .a_prev(a_prev), .n31589(n31589), 
            .b_prev(b_prev), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net), .position_31__N_3836(position_31__N_3836), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 i13648_3_lut (.I0(a_prev_adj_5767), .I1(a_new_adj_5891[1]), 
            .I2(debounce_cnt_N_3833_adj_5769), .I3(GND_net), .O(n31593));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19096_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(\data_in_frame[22] [6]), 
            .I3(rx_data[6]), .O(n32350));
    defparam i19096_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i14173_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n32118));
    defparam i14173_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14170_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n32115));
    defparam i14170_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14167_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n32112));
    defparam i14167_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14163_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n32108));
    defparam i14163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23529_2_lut (.I0(control_mode[7]), .I1(control_mode[6]), .I2(GND_net), 
            .I3(GND_net), .O(n41374));
    defparam i23529_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_2023 (.I0(control_mode[4]), .I1(control_mode[2]), 
            .I2(control_mode[3]), .I3(control_mode[5]), .O(n59660));
    defparam i2_4_lut_adj_2023.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut_4_lut (.I0(reset), .I1(n30362), .I2(\data_in_frame[22] [0]), 
            .I3(rx_data[0]), .O(n59062));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_4_lut_adj_2024 (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), 
            .I2(n6_adj_5846), .I3(n4_adj_5764), .O(n63507));
    defparam i1_2_lut_4_lut_adj_2024.LUT_INIT = 16'hfff7;
    SB_LUT4 i14005_3_lut (.I0(\data_in_frame[16] [7]), .I1(rx_data[7]), 
            .I2(n62228), .I3(GND_net), .O(n31950));   // verilog/coms.v(130[12] 305[6])
    defparam i14005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_2025 (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), 
            .I2(n6_adj_5846), .I3(n41584), .O(n63525));
    defparam i1_2_lut_4_lut_adj_2025.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_4_lut_adj_2026 (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), 
            .I2(n6_adj_5846), .I3(n4_adj_5763), .O(n63489));
    defparam i1_2_lut_4_lut_adj_2026.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_2027 (.I0(hall1), .I1(hall2), .I2(n24553), 
            .I3(GND_net), .O(n4_adj_5851));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_2027.LUT_INIT = 16'hf2f2;
    SB_LUT4 i13797_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n60042), 
            .I3(GND_net), .O(n31742));   // verilog/coms.v(130[12] 305[6])
    defparam i13797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13800_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n60042), 
            .I3(GND_net), .O(n31745));   // verilog/coms.v(130[12] 305[6])
    defparam i13800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71422_bdd_4_lut (.I0(n71422), .I1(neopxl_color[2]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[0]), .O(n71425));
    defparam n71422_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_2028 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5828));
    defparam i5_4_lut_adj_2028.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_2029 (.I0(delay_counter[28]), .I1(n12_adj_5828), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n27501));
    defparam i6_4_lut_adj_2029.LUT_INIT = 16'hfffe;
    SB_LUT4 i4293_4_lut (.I0(n27497), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5716));
    defparam i4293_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_2030 (.I0(n24_adj_5716), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n62593));
    defparam i2_4_lut_adj_2030.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_2031 (.I0(n62593), .I1(delay_counter[18]), .I2(n27494), 
            .I3(GND_net), .O(n62537));
    defparam i2_3_lut_adj_2031.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_2032 (.I0(n62537), .I1(delay_counter[23]), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5844));
    defparam i2_4_lut_adj_2032.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_2033 (.I0(n7_adj_5844), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n27501), .O(n62));
    defparam i4_4_lut_adj_2033.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2034 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n27494));
    defparam i2_3_lut_adj_2034.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut_adj_2035 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_5838));
    defparam i5_3_lut_adj_2035.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_2036 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5837));
    defparam i6_4_lut_adj_2036.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_2037 (.I0(n15_adj_5837), .I1(delay_counter[2]), 
            .I2(n14_adj_5838), .I3(delay_counter[6]), .O(n27497));
    defparam i8_4_lut_adj_2037.LUT_INIT = 16'hfffe;
    SB_LUT4 i13930_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n31875));
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13933_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n31878));
    defparam i13933_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_2038 (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5719));   // verilog/TinyFPGA_B.v(379[12:17])
    defparam i6_4_lut_adj_2038.LUT_INIT = 16'hfffe;
    SB_LUT4 i13936_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n31881));
    defparam i13936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13942_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n31887));
    defparam i13942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13945_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n31890));
    defparam i13945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13948_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n31893));
    defparam i13948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_2039 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5720));   // verilog/TinyFPGA_B.v(379[12:17])
    defparam i5_4_lut_adj_2039.LUT_INIT = 16'hfffe;
    SB_LUT4 i23531_4_lut (.I0(n13_adj_5720), .I1(baudrate[0]), .I2(n14_adj_5719), 
            .I3(n27632), .O(n41376));
    defparam i23531_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i13952_3_lut_4_lut (.I0(reset), .I1(n163), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n31897));
    defparam i13952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_2040 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5829));
    defparam i1_2_lut_adj_2040.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_2041 (.I0(delay_counter[9]), .I1(n4_adj_5829), 
            .I2(delay_counter[10]), .I3(n27497), .O(n62592));
    defparam i2_4_lut_adj_2041.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_3_lut_4_lut_adj_2042 (.I0(n161), .I1(n3491), .I2(n10), 
            .I3(n167), .O(n30370));
    defparam i2_3_lut_4_lut_adj_2042.LUT_INIT = 16'hf7ff;
    SB_LUT4 i2_4_lut_adj_2043 (.I0(n62592), .I1(n27494), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n62445));
    defparam i2_4_lut_adj_2043.LUT_INIT = 16'hffec;
    SB_LUT4 i2_3_lut_4_lut_adj_2044 (.I0(n161), .I1(n3491), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n1_adj_5809), .O(n152));
    defparam i2_3_lut_4_lut_adj_2044.LUT_INIT = 16'hf7ff;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5826));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_2045 (.I0(delay_counter[22]), .I1(n62445), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5827));
    defparam i2_4_lut_adj_2045.LUT_INIT = 16'ha8a0;
    SB_LUT4 i23534_4_lut (.I0(n7_adj_5827), .I1(delay_counter[31]), .I2(n27501), 
            .I3(n8_adj_5826), .O(n1331));   // verilog/TinyFPGA_B.v(381[14:38])
    defparam i23534_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i23606_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(367[12:35])
    defparam i23606_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i591_2_lut (.I0(n1331), .I1(n41376), .I2(GND_net), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(385[18] 387[12])
    defparam i591_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5758));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45208_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64469));
    defparam i45208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5754));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51872_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6917), .I2(n64469), 
            .I3(n25_adj_5834), .O(n17_adj_5833));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i51872_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5756));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_4_lut_adj_2046 (.I0(n260), .I1(n64457), .I2(duty[23]), 
            .I3(n22_adj_5845), .O(n9947));
    defparam i1_4_lut_4_lut_adj_2046.LUT_INIT = 16'h1505;
    SB_LUT4 i49312_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n68582));
    defparam i49312_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45076_2_lut (.I0(color_bit_N_502[2]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n64335));
    defparam i45076_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48890_4_lut (.I0(n64335), .I1(n54699), .I2(n54679), .I3(color_bit_N_502[1]), 
            .O(n67748));   // verilog/neopixel.v(34[12] 113[6])
    defparam i48890_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5742));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i26_4_lut (.I0(n27099), .I1(n67748), .I2(state[1]), .I3(n4), 
            .O(n58944));   // verilog/neopixel.v(34[12] 113[6])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i49125_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n68395));
    defparam i49125_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5740));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49143_2_lut_4_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(current[5]), .I3(current_limit[5]), .O(n68413));
    defparam i49143_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i10_3_lut_3_lut (.I0(current_limit[5]), .I1(current_limit[6]), 
            .I2(current[6]), .I3(GND_net), .O(n10_adj_5738));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48715_4_lut (.I0(n10_adj_5717), .I1(\FRAME_MATCHER.i [0]), 
            .I2(rx_data[6]), .I3(n1_adj_5809), .O(n67750));   // verilog/coms.v(130[12] 305[6])
    defparam i48715_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i16_3_lut (.I0(\data_in_frame[6] [6]), .I1(n67750), .I2(n30423), 
            .I3(GND_net), .O(n58986));   // verilog/coms.v(130[12] 305[6])
    defparam i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2047 (.I0(\data_in_frame[6] [5]), .I1(n30382), 
            .I2(n30423), .I3(rx_data[5]), .O(n59110));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2047.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13621_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n30423), 
            .I3(GND_net), .O(n31566));   // verilog/coms.v(130[12] 305[6])
    defparam i13621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2048 (.I0(\data_in_frame[6] [3]), .I1(n30382), 
            .I2(n30423), .I3(rx_data[3]), .O(n59114));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2048.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2049 (.I0(\data_in_frame[6] [2]), .I1(n30382), 
            .I2(n30423), .I3(rx_data[2]), .O(n59126));
    defparam i12_4_lut_adj_2049.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13612_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n30423), 
            .I3(GND_net), .O(n31557));   // verilog/coms.v(130[12] 305[6])
    defparam i13612_3_lut.LUT_INIT = 16'hcaca;
    coms neopxl_color_23__I_0 (.n2889(n2889), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .clk16MHz(clk16MHz), .n59826(n59826), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n60431(n60431), .GND_net(GND_net), .n31950(n31950), .VCC_net(VCC_net), 
         .\data_in_frame[16] ({\data_in_frame[16] }), .n59825(n59825), .n59824(n59824), 
         .n31947(n31947), .n59823(n59823), .n31262(n31262), .n59770(n59770), 
         .n59822(n59822), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n59821(n59821), .n59820(n59820), .n31257(n31257), .n59819(n59819), 
         .n59818(n59818), .rx_data({rx_data}), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .byte_transmit_counter({Open_3, 
         Open_4, Open_5, Open_6, Open_7, byte_transmit_counter[2:0]}), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n59817(n59817), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n31942(n31942), 
         .n59816(n59816), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n59946(n59946), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n59945(n59945), .control_mode({control_mode}), .n27629(n27629), 
         .n51206(n51206), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n59944(n59944), .n31939(n31939), .n59815(n59815), .displacement({displacement}), 
         .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), .n54181(n54181), 
         .n8(n8_adj_5808), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n59943(n59943), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n59942(n59942), .n31936(n31936), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n59941(n59941), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), .pwm_setpoint({pwm_setpoint}), 
         .n31251(n31251), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n60434(n60434), .n54659(n54659), .LED_c(LED_c), .n59947(n59947), 
         .n59814(n59814), .n59813(n59813), .n59812(n59812), .n59811(n59811), 
         .n59810(n59810), .n59809(n59809), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n59808(n59808), .n59807(n59807), .n60592(n60592), .n59806(n59806), 
         .n59805(n59805), .n59804(n59804), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n59940(n59940), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .n59939(n59939), .n59803(n59803), .n31237(n31237), .n10(n10_adj_5717), 
         .n152(n152), .n30382(n30382), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .n28303(n28303), .n59802(n59802), .n31933(n31933), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n59938(n59938), .n28963(n28963), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .setpoint({setpoint}), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n59937(n59937), .n27161(n27161), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n31930(n31930), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .n59936(n59936), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .n59935(n59935), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .n59934(n59934), .n31927(n31927), .\data_out_frame[3][7] (\data_out_frame[3] [7]), 
         .n59933(n59933), .\data_out_frame[4] ({\data_out_frame[4] }), .n59932(n59932), 
         .n59931(n59931), .n59930(n59930), .n55737(n55737), .n59929(n59929), 
         .n59928(n59928), .n59927(n59927), .n59926(n59926), .n59925(n59925), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .n59924(n59924), .n59801(n59801), 
         .n59800(n59800), .n59799(n59799), .n59798(n59798), .n59797(n59797), 
         .n59796(n59796), .n59923(n59923), .n59795(n59795), .n59922(n59922), 
         .n59794(n59794), .n59793(n59793), .\data_in_frame[3] ({\data_in_frame[3] [7:6], 
         Open_8, Open_9, Open_10, Open_11, Open_12, Open_13}), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n59921(n59921), .n59792(n59792), .n59791(n59791), .n59920(n59920), 
         .n59790(n59790), .n59789(n59789), .n59788(n59788), .n59787(n59787), 
         .n59786(n59786), .n59785(n59785), .n59784(n59784), .n59919(n59919), 
         .n59783(n59783), .\data_in_frame[1] ({\data_in_frame[1] [7:4], 
         Open_14, Open_15, Open_16, Open_17}), .n59782(n59782), .n59781(n59781), 
         .n59780(n59780), .n61872(n61872), .n59779(n59779), .\current[15] (current[15]), 
         .n59778(n59778), .n59777(n59777), .n59918(n59918), .n55561(n55561), 
         .\current[11] (current[11]), .n31897(n31897), .\data_in_frame[14] ({\data_in_frame[14] [7:4], 
         Open_18, Open_19, Open_20, Open_21}), .\current[10] (current[10]), 
         .n59776(n59776), .n59775(n59775), .n24(n24_adj_5841), .\current[9] (current[9]), 
         .n55706(n55706), .n23(n23_adj_5842), .n25(n25_adj_5840), .n59774(n59774), 
         .n59773(n59773), .\current[8] (current[8]), .n59772(n59772), 
         .n59771(n59771), .n59832(n59832), .\data_in_frame[5][4] (\data_in_frame[5] [4]), 
         .\data_in_frame[2][1] (\data_in_frame[2] [1]), .n60470(n60470), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), 
         .n31893(n31893), .n59917(n59917), .\data_out_frame[26][1] (\data_out_frame[26] [1]), 
         .\data_out_frame[26][2] (\data_out_frame[26] [2]), .reset(reset), 
         .n31890(n31890), .\data_in_frame[21] ({\data_in_frame[21] [7], 
         Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, Open_28}), 
         .n59916(n59916), .\data_out_frame[27][1] (\data_out_frame[27] [1]), 
         .\data_out_frame[27][2] (\data_out_frame[27] [2]), .n31887(n31887), 
         .\data_out_frame[11][7] (\data_out_frame[11] [7]), .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), 
         .\data_out_frame[11][6] (\data_out_frame[11] [6]), .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), 
         .\data_out_frame[11][5] (\data_out_frame[11] [5]), .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), 
         .\data_out_frame[11][4] (\data_out_frame[11] [4]), .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), 
         .\data_out_frame[11][3] (\data_out_frame[11] [3]), .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), 
         .\data_out_frame[11][2] (\data_out_frame[11] [2]), .\encoder0_position_scaled[2] (encoder0_position_scaled[2]), 
         .\data_out_frame[11][1] (\data_out_frame[11] [1]), .\encoder0_position_scaled[1] (encoder0_position_scaled[1]), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n59915(n59915), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), 
         .n59914(n59914), .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), 
         .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), 
         .n31881(n31881), .\data_in_frame[14][2] (\data_in_frame[14] [2]), 
         .n31878(n31878), .\data_in_frame[14][1] (\data_in_frame[14] [1]), 
         .n59913(n59913), .n31875(n31875), .\data_in_frame[14][0] (\data_in_frame[14] [0]), 
         .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), 
         .n59912(n59912), .n59911(n59911), .\data_in_frame[5][5] (\data_in_frame[5] [5]), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\encoder0_position_scaled[23] (encoder0_position_scaled[23]), 
         .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), .\encoder0_position_scaled[21] (encoder0_position_scaled[21]), 
         .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), 
         .n60254(n60254), .\data_in_frame[20] ({\data_in_frame[20] }), .\data_in_frame[21][0] (\data_in_frame[21] [0]), 
         .\data_in_frame[18] ({Open_29, \data_in_frame[18] [6:5], Open_30, 
         Open_31, Open_32, Open_33, Open_34}), .\data_in_frame[21][1] (\data_in_frame[21] [1]), 
         .\data_in_frame[21][4] (\data_in_frame[21] [4]), .\data_in_frame[19] ({Open_35, 
         Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, \data_in_frame[19] [0]}), 
         .\data_in_frame[21][5] (\data_in_frame[21] [5]), .\data_in_frame[18][1] (\data_in_frame[18] [1]), 
         .\data_in_frame[18][3] (\data_in_frame[18] [3]), .\data_in_frame[18][0] (\data_in_frame[18] [0]), 
         .\data_in_frame[17][5] (\data_in_frame[17] [5]), .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), 
         .\data_in_frame[18][4] (\data_in_frame[18] [4]), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[19][7] (\data_in_frame[19] [7]), .\data_in_frame[17][7] (\data_in_frame[17] [7]), 
         .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), .\data_in_frame[18][2] (\data_in_frame[18] [2]), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[6][3] (\data_in_frame[6] [3]), 
         .n31847(n31847), .\data_in_frame[6][5] (\data_in_frame[6] [5]), 
         .\data_in_frame[5][0] (\data_in_frame[5] [0]), .n31844(n31844), 
         .n31841(n31841), .\data_out_frame[8][7] (\data_out_frame[8] [7]), 
         .\data_in_frame[5][6] (\data_in_frame[5] [6]), .\data_in_frame[5][7] (\data_in_frame[5] [7]), 
         .n31836(n31836), .n59910(n59910), .\data_out_frame[8][6] (\data_out_frame[8] [6]), 
         .n31833(n31833), .n59909(n59909), .n31830(n31830), .n31827(n31827), 
         .n31824(n31824), .\data_out_frame[8][5] (\data_out_frame[8] [5]), 
         .\data_in_frame[19][2] (\data_in_frame[19] [2]), .\data_in_frame[21][3] (\data_in_frame[21] [3]), 
         .\data_in_frame[17][0] (\data_in_frame[17] [0]), .\data_out_frame[8][4] (\data_out_frame[8] [4]), 
         .\data_in_frame[17][6] (\data_in_frame[17] [6]), .\data_out_frame[8][3] (\data_out_frame[8] [3]), 
         .n31797(n31797), .n31794(n31794), .n31791(n31791), .n31788(n31788), 
         .n31785(n31785), .\data_out_frame[8][2] (\data_out_frame[8] [2]), 
         .n31782(n31782), .\data_out_frame[8][1] (\data_out_frame[8] [1]), 
         .n31779(n31779), .n31776(n31776), .n31773(n31773), .n31770(n31770), 
         .n31767(n31767), .\data_out_frame[7] ({\data_out_frame[7] }), .n59122(n59122), 
         .\data_in_frame[6][0] (\data_in_frame[6] [0]), .n31557(n31557), 
         .\data_in_frame[6][1] (\data_in_frame[6] [1]), .n59126(n59126), 
         .\data_in_frame[6][2] (\data_in_frame[6] [2]), .n59114(n59114), 
         .n31566(n31566), .\data_in_frame[6][4] (\data_in_frame[6] [4]), 
         .n59110(n59110), .n58986(n58986), .\data_in_frame[6][6] (\data_in_frame[6] [6]), 
         .n59908(n59908), .n31745(n31745), .n31742(n31742), .n31739(n31739), 
         .n31736(n31736), .n31733(n31733), .n59907(n59907), .\data_in_frame[17][3] (\data_in_frame[17] [3]), 
         .DE_c(DE_c), .\data_in_frame[2][0] (\data_in_frame[2] [0]), .\data_in_frame[17][4] (\data_in_frame[17] [4]), 
         .n59906(n59906), .n59905(n59905), .n59904(n59904), .n59833(n59833), 
         .n59903(n59903), .n59902(n59902), .n59901(n59901), .n59900(n59900), 
         .n59899(n59899), .n59898(n59898), .n59897(n59897), .n59896(n59896), 
         .n59895(n59895), .n59894(n59894), .n59893(n59893), .n59892(n59892), 
         .n59891(n59891), .n59890(n59890), .n59889(n59889), .n59888(n59888), 
         .n59887(n59887), .n59886(n59886), .n59885(n59885), .n59884(n59884), 
         .n59883(n59883), .n59882(n59882), .n59881(n59881), .n59880(n59880), 
         .n59879(n59879), .n59878(n59878), .n32669(n32669), .n31321(n31321), 
         .n59877(n59877), .n59876(n59876), .n59875(n59875), .n59874(n59874), 
         .n59873(n59873), .n59872(n59872), .n59871(n59871), .n59870(n59870), 
         .n59869(n59869), .n59868(n59868), .n59867(n59867), .n59866(n59866), 
         .n59865(n59865), .n59864(n59864), .n59863(n59863), .n59862(n59862), 
         .n59861(n59861), .n59860(n59860), .n59859(n59859), .n59834(n59834), 
         .n59858(n59858), .n32691(n32691), .n31299(n31299), .n59857(n59857), 
         .n59856(n59856), .n59855(n59855), .n59854(n59854), .n31294(n31294), 
         .n59853(n59853), .n59852(n59852), .n59851(n59851), .n59850(n59850), 
         .n59849(n59849), .n59848(n59848), .n59847(n59847), .n59846(n59846), 
         .n59845(n59845), .n32706(n32706), .n31284(n31284), .n59844(n59844), 
         .n59843(n59843), .n59842(n59842), .n31590(n31590), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n59841(n59841), .n59840(n59840), .n59839(n59839), .n31277(n31277), 
         .n59838(n59838), .n59837(n59837), .n59836(n59836), .n59835(n59835), 
         .n59831(n59831), .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .n59830(n59830), 
         .\data_in_frame[2][4] (\data_in_frame[2] [4]), .\data_in_frame[5][1] (\data_in_frame[5] [1]), 
         .\data_in_frame[2][5] (\data_in_frame[2] [5]), .n59829(n59829), 
         .\data_in_frame[5][2] (\data_in_frame[5] [2]), .ID({ID}), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .\data_in_frame[1][1] (\data_in_frame[1] [1]), .\data_in_frame[3][0] (\data_in_frame[3] [0]), 
         .\data_in_frame[3][2] (\data_in_frame[3] [2]), .\data_in_frame[1][0] (\data_in_frame[1] [0]), 
         .\data_in_frame[2][2] (\data_in_frame[2] [2]), .deadband({deadband}), 
         .n71521(n71521), .\data_in_frame[22][4] (\data_in_frame[22] [4]), 
         .\data_in_frame[22][6] (\data_in_frame[22] [6]), .\data_in_frame[22][1] (\data_in_frame[22] [1]), 
         .\data_in_frame[22][0] (\data_in_frame[22] [0]), .\data_in_frame[22][3] (\data_in_frame[22] [3]), 
         .\data_in_frame[22][2] (\data_in_frame[22] [2]), .IntegralLimit({IntegralLimit}), 
         .\Kp[0] (Kp[0]), .\Ki[0] (Ki[0]), .PWMLimit({PWMLimit}), .n31269(n31269), 
         .n161(n161), .n59828(n59828), .n31954(n31954), .n60741(n60741), 
         .n62047(n62047), .n31965(n31965), .n31968(n31968), .n31971(n31971), 
         .n31974(n31974), .n31977(n31977), .n59150(n59150), .n59148(n59148), 
         .n59146(n59146), .n31990(n31990), .n59144(n59144), .n31996(n31996), 
         .n59142(n59142), .n59140(n59140), .n59138(n59138), .n31440(n31440), 
         .n59136(n59136), .n31443(n31443), .n32066(n32066), .n31446(n31446), 
         .n31449(n31449), .\data_in_frame[2][3] (\data_in_frame[2] [3]), 
         .n32078(n32078), .n31452(n31452), .n32088(n32088), .n31455(n31455), 
         .n32092(n32092), .n59062(n59062), .n32108(n32108), .n32112(n32112), 
         .n32115(n32115), .n32118(n32118), .n32350(n32350), .n31482(n31482), 
         .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
         .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), 
         .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), 
         .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), 
         .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
         .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), 
         .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
         .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .n31488(n31488), .n32229(n32229), 
         .neopxl_color({neopxl_color}), .n32228(n32228), .n32227(n32227), 
         .n32226(n32226), .n32225(n32225), .n32222(n32222), .n32221(n32221), 
         .n32220(n32220), .n32218(n32218), .n32217(n32217), .n32216(n32216), 
         .n32215(n32215), .n32214(n32214), .n32213(n32213), .n32212(n32212), 
         .n32211(n32211), .n32210(n32210), .n32209(n32209), .n32208(n32208), 
         .n32207(n32207), .n32206(n32206), .current_limit({current_limit}), 
         .n31463(n31463), .n31462(n31462), .n59827(n59827), .n32203(n32203), 
         .n32202(n32202), .n32201(n32201), .n32200(n32200), .n32199(n32199), 
         .n32197(n32197), .n32196(n32196), .n32195(n32195), .n32193(n32193), 
         .n32192(n32192), .n32191(n32191), .n32190(n32190), .n32189(n32189), 
         .n32188(n32188), .n32187(n32187), .n32186(n32186), .n32185(n32185), 
         .n31491(n31491), .n31500(n31500), .n31503(n31503), .n60669(n60669), 
         .n167(n167), .n28330(n28330), .n54982(n54982), .n60241(n60241), 
         .n54578(n54578), .n3491(n3491), .rx_data_ready(rx_data_ready), 
         .n61989(n61989), .n71389(n71389), .n71401(n71401), .n30156(n30156), 
         .n60391(n60391), .n1(n1_adj_5809), .n144(n144), .n163(n163), 
         .n60044(n60044), .n60042(n60042), .n60039(n60039), .n67759(n67759), 
         .n28021(n28021), .n30370(n30370), .n10_adj_6(n10), .n30449(n30449), 
         .n70677(n70677), .n30366(n30366), .n30416(n30416), .\current[7] (current[7]), 
         .n24903(n24903), .\current[6] (current[6]), .\current[5] (current[5]), 
         .n24877(n24877), .\current[4] (current[4]), .\current[3] (current[3]), 
         .\current[2] (current[2]), .\current[1] (current[1]), .\current[0] (current[0]), 
         .n30414(n30414), .n30362(n30362), .n30452(n30452), .n30447(n30447), 
         .n62670(n62670), .n62228(n62228), .n30368(n30368), .control_update(control_update), 
         .n41374(n41374), .n27538(n27538), .tx_active(tx_active), .n45(n45), 
         .n31(n31), .n28(n28), .n30(n30_adj_5807), .n30423(n30423), 
         .n60355(n60355), .n60038(n60038), .n64880(n64880), .n64878(n64878), 
         .n64890(n64890), .n64891(n64891), .n64615(n64615), .n64614(n64614), 
         .n1_adj_7(n1), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_5927}), 
         .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), .r_Clock_Count({r_Clock_Count_adj_5928}), 
         .n29824(n29824), .\r_Bit_Index[0] (r_Bit_Index_adj_5929[0]), .n59688(n59688), 
         .n31480(n31480), .n63187(n63187), .n27(n27), .n32074(n32074), 
         .n71705(n71705), .n63177(n63177), .n5235(n5235), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
         .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n29(n29), .n23_adj_8(n23_adj_5843), 
         .n61652(n61652), .n6(n6_adj_5825), .n60832(n60832), .tx_enable(tx_enable), 
         .n31953(n31953), .baudrate({baudrate}), .n31945(n31945), .n27632(n27632), 
         .\r_SM_Main[2]_adj_9 (r_SM_Main[2]), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
         .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), 
         .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), 
         .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .r_Clock_Count_adj_22({r_Clock_Count}), 
         .n31702(n31702), .\r_SM_Main[1]_adj_18 (r_SM_Main[1]), .n29821(n29821), 
         .r_Bit_Index({r_Bit_Index}), .n32083(n32083), .n55814(n55814), 
         .n32231(n32231), .n32087(n32087), .n32021(n32021), .n32020(n32020), 
         .n31961(n31961), .n6_adj_20(n6_adj_5846), .n5232(n5232), .n4(n4_adj_5763), 
         .n59686(n59686), .n63199(n63199), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .n4_adj_21(n4_adj_5764), .n63175(n63175), .n41584(n41584), .n29817(n29817), 
         .n60834(n60834)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 LessThan_1180_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5819));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1180_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48548_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n67818));   // verilog/uart_rx.v(119[17:57])
    defparam i48548_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i13214_2_lut_3_lut (.I0(n25001), .I1(dti), .I2(n15_adj_5760), 
            .I3(GND_net), .O(n31159));
    defparam i13214_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_3_lut_adj_2050 (.I0(n25001), .I1(dti), .I2(n15_adj_5760), 
            .I3(GND_net), .O(n29976));
    defparam i1_2_lut_3_lut_adj_2050.LUT_INIT = 16'hf8f8;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_2051 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(n28963), .I3(n54578), .O(n4_adj_5836));
    defparam i1_2_lut_3_lut_4_lut_adj_2051.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_1180_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5818));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1180_i4_4_lut.LUT_INIT = 16'h4d0c;
    TLI4970 tli (.clk16MHz(clk16MHz), .n29799(n29799), .\current[15] (current[15]), 
            .n31638(n31638), .\current[1] (current[1]), .n31637(n31637), 
            .\current[2] (current[2]), .n31636(n31636), .\current[3] (current[3]), 
            .n31635(n31635), .\current[4] (current[4]), .n31634(n31634), 
            .\current[5] (current[5]), .n31633(n31633), .\current[6] (current[6]), 
            .n31632(n31632), .\current[7] (current[7]), .n31631(n31631), 
            .\current[8] (current[8]), .n31630(n31630), .\current[9] (current[9]), 
            .n31629(n31629), .\current[10] (current[10]), .n31628(n31628), 
            .\current[11] (current[11]), .state_7__N_4319(state_7__N_4319), 
            .GND_net(GND_net), .VCC_net(VCC_net), .CS_c(CS_c), .n31471(n31471), 
            .\current[0] (current[0]), .n32396(n32396), .\data[15] (data_adj_5911[15]), 
            .n32395(n32395), .\data[12] (data_adj_5911[12]), .n32394(n32394), 
            .\data[11] (data_adj_5911[11]), .n32393(n32393), .\data[10] (data_adj_5911[10]), 
            .n32392(n32392), .\data[9] (data_adj_5911[9]), .n32391(n32391), 
            .\data[8] (data_adj_5911[8]), .n32390(n32390), .\data[7] (data_adj_5911[7]), 
            .n32389(n32389), .\data[6] (data_adj_5911[6]), .n32388(n32388), 
            .\data[5] (data_adj_5911[5]), .n32387(n32387), .\data[4] (data_adj_5911[4]), 
            .n32386(n32386), .\data[3] (data_adj_5911[3]), .n32385(n32385), 
            .\data[2] (data_adj_5911[2]), .n32384(n32384), .\data[1] (data_adj_5911[1]), 
            .n32101(n32101), .\data[0] (data_adj_5911[0]), .CS_CLK_c(CS_CLK_c), 
            .n27661(n27661), .n27667(n27667), .n11(n11_adj_5779), .n27680(n27680), 
            .n27643(n27643), .n5(n5_adj_5778), .n5_adj_4(n5_adj_5806), 
            .n41527(n41527), .n9(n9_adj_5780)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(406[11] 412[4])
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n71392));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 LessThan_1180_i8_3_lut (.I0(n6_adj_5819), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5821), .I3(GND_net), .O(n8_adj_5820));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1180_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51454_4_lut (.I0(n8_adj_5820), .I1(n4_adj_5818), .I2(n9_adj_5821), 
            .I3(n67818), .O(n70724));   // verilog/uart_rx.v(119[17:57])
    defparam i51454_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51455_3_lut (.I0(n70724), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n70725));   // verilog/uart_rx.v(119[17:57])
    defparam i51455_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_2052 (.I0(n6_adj_5846), .I1(r_SM_Main[1]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5764), .O(n63435));
    defparam i1_2_lut_4_lut_adj_2052.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_2053 (.I0(n6_adj_5846), .I1(r_SM_Main[1]), 
            .I2(r_Bit_Index[0]), .I3(n41584), .O(n63471));
    defparam i1_2_lut_4_lut_adj_2053.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_2054 (.I0(n6_adj_5846), .I1(r_SM_Main[1]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5763), .O(n63453));
    defparam i1_2_lut_4_lut_adj_2054.LUT_INIT = 16'hfffb;
    SB_LUT4 i51352_3_lut (.I0(n70725), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n70622));   // verilog/uart_rx.v(119[17:57])
    defparam i51352_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51218_3_lut (.I0(n70622), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5232));   // verilog/uart_rx.v(119[17:57])
    defparam i51218_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut (.I0(control_mode[7]), .I1(control_mode[6]), 
            .I2(n59660), .I3(control_mode[1]), .O(n54181));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2055 (.I0(o_Rx_DV_N_3488[12]), .I1(n5232), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63489), .O(n63495));
    defparam i1_4_lut_adj_2055.LUT_INIT = 16'hfffe;
    SB_LUT4 i14761_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n32706));   // verilog/coms.v(130[12] 305[6])
    defparam i14761_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2056 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5843), 
            .I3(n63495), .O(n63501));
    defparam i1_4_lut_adj_2056.LUT_INIT = 16'hfffe;
    SB_LUT4 i14008_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n63501), 
            .I3(n27), .O(n31953));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14008_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_4_lut_adj_2057 (.I0(control_mode[1]), .I1(n59660), 
            .I2(control_mode[7]), .I3(control_mode[6]), .O(n27629));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_3_lut_4_lut_adj_2057.LUT_INIT = 16'hfffd;
    pwm PWM (.n2889(n2889), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .reset(reset), 
        .GND_net(GND_net), .\pwm_counter[6] (pwm_counter[6]), .\pwm_counter[8] (pwm_counter[8]), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint}), .n17(n17_adj_5771), 
        .n13(n13_adj_5772)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    motorControl control (.\Ki[8] (Ki[8]), .n335({n336, n337, n338, 
            n339, n340, n341, n342, n343, n344, n345, n346, 
            n347, n348, n349, n350, n351, n352, n353, n354, 
            n355, n356, n357, n358, n359}), .GND_net(GND_net), .\Ki[9] (Ki[9]), 
            .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .setpoint({setpoint}), 
            .IntegralLimit({IntegralLimit}), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Kp[6] (Kp[6]), .\Ki[2] (Ki[2]), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .\Ki[3] (Ki[3]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Ki[4] (Ki[4]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .n8(n8_adj_5808), .\motor_state[9] (motor_state[9]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Ki[5] (Ki[5]), .\Kp[15] (Kp[15]), 
            .\motor_state[8] (motor_state[8]), .\Ki[6] (Ki[6]), .\motor_state[7] (motor_state[7]), 
            .\Ki[7] (Ki[7]), .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .\motor_state[1] (motor_state[1]), 
            .VCC_net(VCC_net), .PWMLimit({PWMLimit}), .n32332(n32332), 
            .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), .n32331(n32331), 
            .n32330(n32330), .n32329(n32329), .n32328(n32328), .n32327(n32327), 
            .n32326(n32326), .n32325(n32325), .n32324(n32324), .n32323(n32323), 
            .n32322(n32322), .n32321(n32321), .n32320(n32320), .n32319(n32319), 
            .n32318(n32318), .n32317(n32317), .n32316(n32316), .n32315(n32315), 
            .n32314(n32314), .n32313(n32313), .n32312(n32312), .n32311(n32311), 
            .n32308(n32308), .n31436(n31436), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .\motor_state[11] (motor_state[11]), 
            .deadband({deadband}), .n41880(n41880), .\control_mode[7] (control_mode[7]), 
            .\control_mode[6] (control_mode[6]), .\control_mode[1] (control_mode[1]), 
            .\control_mode[0] (control_mode[0]), .n27629(n27629), .n29776(n29776), 
            .n54181(n54181), .\displacement[0] (displacement[0]), .n59660(n59660), 
            .n27538(n27538), .n28(n28), .n31(n31), .n45(n45), .n30(n30_adj_5807), 
            .n70677(n70677)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    EEPROM eeprom (.enable_slow_N_4213(enable_slow_N_4213), .clk16MHz(clk16MHz), 
           .n29874(n29874), .data({data_adj_5904}), .ID({ID}), .GND_net(GND_net), 
           .baudrate({baudrate}), .n31646(n31646), .n31645(n31645), .n31644(n31644), 
           .n31643(n31643), .n31642(n31642), .n31641(n31641), .n31640(n31640), 
           .n31639(n31639), .\state_7__N_3918[0] (state_7__N_3918[0]), .data_ready(data_ready), 
           .\state_7__N_4110[0] (state_7__N_4110[0]), .\state[0] (state_adj_5937[0]), 
           .scl_enable(scl_enable), .VCC_net(VCC_net), .sda_enable(sda_enable), 
           .n32362(n32362), .n32360(n32360), .n32356(n32356), .n32339(n32339), 
           .n32338(n32338), .n32337(n32337), .n32335(n32335), .n32065(n32065), 
           .n8(n8_adj_5847), .n6722(n6722), .scl(scl), .sda_out(sda_out), 
           .\state_7__N_4126[3] (state_7__N_4126[3]), .n41430(n41430), .n6(n6_adj_5830), 
           .n4(n4_adj_5761), .n4_adj_3(n4_adj_5762), .n41590(n41590), 
           .n10(n10_adj_5824), .n27672(n27672), .n27624(n27624)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(392[10] 404[6])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (n29957, bit_ctr, clk16MHz, 
            GND_net, state, \neopxl_color[5] , \neopxl_color[4] , \color_bit_N_502[1] , 
            n31755, VCC_net, n58944, n31687, t0, n31686, n31685, 
            timer, n31684, n31683, n31682, \bit_ctr[3] , n31681, 
            n31680, n31679, n31678, \bit_ctr[0] , NEOPXL_c, n31481, 
            n27099, LED_c, n41559, n54699, \color_bit_N_502[2] , n3180, 
            \neopxl_color[14] , \neopxl_color[15] , \neopxl_color[12] , 
            \neopxl_color[13] , n71341, n54679, n71425, n71395, \neopxl_color[6] , 
            \neopxl_color[7] ) /* synthesis syn_module_defined=1 */ ;
    output n29957;
    output [4:0]bit_ctr;
    input clk16MHz;
    input GND_net;
    output [1:0]state;
    input \neopxl_color[5] ;
    input \neopxl_color[4] ;
    output \color_bit_N_502[1] ;
    input n31755;
    input VCC_net;
    input n58944;
    input n31687;
    output [10:0]t0;
    input n31686;
    input n31685;
    output [10:0]timer;
    input n31684;
    input n31683;
    input n31682;
    output \bit_ctr[3] ;
    input n31681;
    input n31680;
    input n31679;
    input n31678;
    output \bit_ctr[0] ;
    output NEOPXL_c;
    input n31481;
    output n27099;
    input LED_c;
    output n41559;
    output n54699;
    output \color_bit_N_502[2] ;
    output n3180;
    input \neopxl_color[14] ;
    input \neopxl_color[15] ;
    input \neopxl_color[12] ;
    input \neopxl_color[13] ;
    input n71341;
    output n54679;
    input n71425;
    input n71395;
    input \neopxl_color[6] ;
    input \neopxl_color[7] ;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n149;
    
    wire n31392;
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n62542, \neo_pixel_transmitter.done , 
        start_N_507, n59204, start, n27640, n6, n27655, n27657, 
        n59976, n61029, n15, n53, n32, n62951, n71356, n71359;
    wire [10:0]n49;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    
    wire n23169, n29951, n30869;
    wire [1:0]state_1__N_451;
    
    wire n29766, n30868, one_wire_N_499, n44, n62668, n61035, n15_adj_5699, 
        n62044, n41482, n81, n60950, n6_adj_5700, n41947;
    wire [10:0]n1;
    
    wire n52820, n52819, n52818, n53342, n53341, n52817, n52816, 
        n53340, n53339, n52815, n52814, n53338, n53337, n53336, 
        n52813, n53335, n53334, n52812, n52811, n53333, n41715, 
        n7217, n27611, n27532, n25, n60014, n22, n67783, n67781, 
        n8_adj_5703, n24776, n67422, n60952, n62577, n67790, n68, 
        n64708, n64707, n64709, n64642, n64641, n64643;
    
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr[4]), .C(clk16MHz), .E(n29957), .D(n149[4]), 
            .R(n31392));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n62542), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n59204), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i1_2_lut (.I0(n27640), .I1(t1[8]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/neopixel.v(100[14:42])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(t1[10]), .I1(n27655), .I2(t1[2]), .I3(n6), 
            .O(n27657));   // verilog/neopixel.v(100[14:42])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i22_4_lut (.I0(n59976), .I1(n61029), .I2(state[1]), .I3(start), 
            .O(n59204));
    defparam i22_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i51801_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i51801_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n15), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n53));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i3_4_lut (.I0(n27640), .I1(n32), .I2(t1[10]), .I3(t1[8]), 
            .O(n62951));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut (.I0(state[1]), .I1(n62951), .I2(start), .I3(GND_net), 
            .O(n62542));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_1__I_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 n71356_bdd_4_lut (.I0(n71356), .I1(\neopxl_color[5] ), .I2(\neopxl_color[4] ), 
            .I3(\color_bit_N_502[1] ), .O(n71359));
    defparam n71356_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(VCC_net), .D(n31755));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n58944));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n31687));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n31686));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n31685));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2040__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n31684));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n31683));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n31682));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n29957), 
            .D(n149[2]), .R(n31392));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(\bit_ctr[3] ), .C(clk16MHz), .E(n29957), 
            .D(n149[3]), .R(n31392));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n31681));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n31680));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n31679));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n31678));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i0 (.Q(\bit_ctr[0] ), .C(clk16MHz), .E(n29951), 
            .D(n23169), .R(n30869));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n29766), .D(state_1__N_451[0]), 
            .S(n30868));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n44), .D(one_wire_N_499), 
            .R(n62668));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n27657), .I3(state[1]), .O(n62668));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1774 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n61035), .I3(n15_adj_5699), .O(n62044));
    defparam i2_3_lut_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i41806_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n27657), .I3(GND_net), .O(n61029));
    defparam i41806_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n31481));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_LUT4 i1_4_lut_4_lut (.I0(n27099), .I1(state[1]), .I2(n41482), .I3(state[0]), 
            .O(n29766));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hee2e;
    SB_LUT4 i1_2_lut_3_lut (.I0(n27099), .I1(state[1]), .I2(n29951), .I3(GND_net), 
            .O(n29957));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n29951));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i12924_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n30869));   // verilog/neopixel.v(35[4] 112[11])
    defparam i12924_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_adj_1775 (.I0(\bit_ctr[3] ), .I1(n41559), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n54699));
    defparam i1_2_lut_3_lut_adj_1775.LUT_INIT = 16'h7878;
    SB_LUT4 i41729_2_lut (.I0(t1[10]), .I1(t1[9]), .I2(GND_net), .I3(GND_net), 
            .O(n60950));
    defparam i41729_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41812_4_lut (.I0(t1[8]), .I1(n60950), .I2(n6_adj_5700), .I3(t1[5]), 
            .O(n61035));
    defparam i41812_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF timer_2040__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 i24096_2_lut_3_lut (.I0(\bit_ctr[3] ), .I1(n41559), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n41947));
    defparam i24096_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF timer_2040__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2040__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n52820), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1776 (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr_c[2]), .I3(GND_net), .O(\color_bit_N_502[2] ));
    defparam i1_2_lut_3_lut_adj_1776.LUT_INIT = 16'h1e1e;
    SB_LUT4 i23713_2_lut_3_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n41559));
    defparam i23713_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n52819), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n52819), .I0(timer[9]), .I1(n1[9]), 
            .CO(n52820));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n52818), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n52818), .I0(timer[8]), .I1(n1[8]), 
            .CO(n52819));
    SB_LUT4 timer_2040_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n53342), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2040_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n53341), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n52817), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n52817), .I0(timer[7]), .I1(n1[7]), 
            .CO(n52818));
    SB_CARRY timer_2040_add_4_11 (.CI(n53341), .I0(GND_net), .I1(timer[9]), 
            .CO(n53342));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n52816), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2040_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n53340), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_10 (.CI(n53340), .I0(GND_net), .I1(timer[8]), 
            .CO(n53341));
    SB_LUT4 timer_2040_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n53339), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n52816), .I0(timer[6]), .I1(n1[6]), 
            .CO(n52817));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n52815), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n52815), .I0(timer[5]), .I1(n1[5]), 
            .CO(n52816));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n52814), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n52814), .I0(timer[4]), .I1(n1[4]), 
            .CO(n52815));
    SB_CARRY timer_2040_add_4_9 (.CI(n53339), .I0(GND_net), .I1(timer[7]), 
            .CO(n53340));
    SB_LUT4 timer_2040_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n53338), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_8 (.CI(n53338), .I0(GND_net), .I1(timer[6]), 
            .CO(n53339));
    SB_LUT4 timer_2040_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n53337), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_7 (.CI(n53337), .I0(GND_net), .I1(timer[5]), 
            .CO(n53338));
    SB_LUT4 timer_2040_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n53336), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n52813), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_6 (.CI(n53336), .I0(GND_net), .I1(timer[4]), 
            .CO(n53337));
    SB_LUT4 timer_2040_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n53335), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_5 (.CI(n53335), .I0(GND_net), .I1(timer[3]), 
            .CO(n53336));
    SB_LUT4 timer_2040_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n53334), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n52813), .I0(timer[3]), .I1(n1[3]), 
            .CO(n52814));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n52812), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n52812), .I0(timer[2]), .I1(n1[2]), 
            .CO(n52813));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n52811), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_4 (.CI(n53334), .I0(GND_net), .I1(timer[2]), 
            .CO(n53335));
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n52811), .I0(timer[1]), .I1(n1[1]), 
            .CO(n52812));
    SB_LUT4 timer_2040_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n53333), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_3 (.CI(n53333), .I0(GND_net), .I1(timer[1]), 
            .CO(n53334));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n52811));
    SB_LUT4 timer_2040_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2040_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n53333));
    SB_LUT4 i23869_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n41715));
    defparam i23869_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2212_2_lut_3_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2212_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2214_2_lut_3_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n7217));   // verilog/neopixel.v(65[23:32])
    defparam i2214_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1777 (.I0(n15), .I1(n15_adj_5699), .I2(state[0]), 
            .I3(n27611), .O(n59976));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut_adj_1777.LUT_INIT = 16'h3500;
    SB_LUT4 i1_2_lut_4_lut_adj_1778 (.I0(n15), .I1(n15_adj_5699), .I2(state[0]), 
            .I3(n27532), .O(n27099));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut_adj_1778.LUT_INIT = 16'h3500;
    SB_LUT4 i46_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25));
    defparam i46_3_lut_4_lut_3_lut.LUT_INIT = 16'h1818;
    SB_LUT4 i3_3_lut_4_lut (.I0(t1[1]), .I1(t1[3]), .I2(t1[2]), .I3(n60014), 
            .O(n15));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i47_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n22));
    defparam i47_3_lut_4_lut_3_lut.LUT_INIT = 16'h8181;
    SB_LUT4 i49189_4_lut (.I0(n22), .I1(n25), .I2(n41715), .I3(state[0]), 
            .O(n67783));
    defparam i49189_4_lut.LUT_INIT = 16'h0c0a;
    SB_LUT4 i50381_4_lut (.I0(n67783), .I1(t1[4]), .I2(t1[2]), .I3(n61035), 
            .O(n67781));
    defparam i50381_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i45_3_lut (.I0(n67781), .I1(state[1]), .I2(start), .I3(GND_net), 
            .O(n3180));
    defparam i45_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i3_3_lut_4_lut_adj_1779 (.I0(\bit_ctr[3] ), .I1(n41559), .I2(n54699), 
            .I3(\bit_ctr[0] ), .O(n8_adj_5703));
    defparam i3_3_lut_4_lut_adj_1779.LUT_INIT = 16'hff9f;
    SB_LUT4 i2_3_lut_4_lut_adj_1780 (.I0(t1[1]), .I1(t1[0]), .I2(t1[4]), 
            .I3(t1[3]), .O(n27655));   // verilog/neopixel.v(60[15:45])
    defparam i2_3_lut_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_4_lut_adj_1781 (.I0(t1[9]), .I1(t1[6]), .I2(t1[7]), 
            .I3(t1[5]), .O(n27640));   // verilog/neopixel.v(100[14:42])
    defparam i3_3_lut_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i5579_3_lut_4_lut (.I0(\bit_ctr[0] ), .I1(start), .I2(n27611), 
            .I3(n24776), .O(n23169));   // verilog/neopixel.v(35[4] 112[11])
    defparam i5579_3_lut_4_lut.LUT_INIT = 16'haa9a;
    SB_LUT4 state_1__I_0_103_Mux_0_i1_3_lut_4_lut (.I0(n15), .I1(t1[2]), 
            .I2(n27655), .I3(state[0]), .O(n24776));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_103_Mux_0_i1_3_lut_4_lut.LUT_INIT = 16'hf3aa;
    SB_LUT4 i48152_2_lut_3_lut (.I0(n54699), .I1(\bit_ctr[3] ), .I2(n41559), 
            .I3(GND_net), .O(n67422));   // verilog/neopixel.v(24[26:38])
    defparam i48152_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i41731_2_lut_3_lut (.I0(n27657), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n60952));
    defparam i41731_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1782 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(t1[2]), .I3(n27655), .O(n62577));
    defparam i2_3_lut_4_lut_adj_1782.LUT_INIT = 16'h0080;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49482_3_lut (.I0(n27657), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n67790));
    defparam i49482_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i72_4_lut (.I0(n62044), .I1(n67790), .I2(state[1]), .I3(start), 
            .O(n68));
    defparam i72_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i51890_4_lut (.I0(n61035), .I1(n68), .I2(n62577), .I3(n53), 
            .O(n44));
    defparam i51890_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23636_2_lut (.I0(n27657), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n41482));
    defparam i23636_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(start), .I1(n60952), .I2(state[1]), .I3(n59976), 
            .O(n30868));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i45438_3_lut (.I0(\neopxl_color[14] ), .I1(\neopxl_color[15] ), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n64708));
    defparam i45438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45437_3_lut (.I0(\neopxl_color[12] ), .I1(\neopxl_color[13] ), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n64707));
    defparam i45437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45439_4_lut (.I0(n64708), .I1(n71341), .I2(n54699), .I3(n54679), 
            .O(n64709));
    defparam i45439_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45372_4_lut (.I0(n64709), .I1(n64707), .I2(n54699), .I3(\color_bit_N_502[1] ), 
            .O(n64642));
    defparam i45372_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i45371_3_lut (.I0(n71425), .I1(n71359), .I2(\color_bit_N_502[2] ), 
            .I3(GND_net), .O(n64641));
    defparam i45371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45373_4_lut (.I0(n64642), .I1(n71395), .I2(n54699), .I3(\color_bit_N_502[2] ), 
            .O(n64643));
    defparam i45373_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i23535_4_lut (.I0(n64643), .I1(n81), .I2(n64641), .I3(n67422), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i23535_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2219_2_lut_4_lut (.I0(\bit_ctr[3] ), .I1(bit_ctr[1]), .I2(\bit_ctr[0] ), 
            .I3(bit_ctr_c[2]), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2219_2_lut_4_lut.LUT_INIT = 16'h6aaa;
    SB_LUT4 bit_ctr_0__bdd_4_lut_52082_4_lut (.I0(\bit_ctr[0] ), .I1(\neopxl_color[6] ), 
            .I2(\neopxl_color[7] ), .I3(bit_ctr[1]), .O(n71356));
    defparam bit_ctr_0__bdd_4_lut_52082_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_4_lut_4_lut_adj_1783 (.I0(n15), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(n15_adj_5699), .O(n32));
    defparam i1_4_lut_4_lut_adj_1783.LUT_INIT = 16'h14d7;
    SB_LUT4 i2_2_lut (.I0(t1[6]), .I1(t1[7]), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5700));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1784 (.I0(\neo_pixel_transmitter.done ), .I1(n27640), 
            .I2(t1[10]), .I3(t1[8]), .O(n27611));
    defparam i3_4_lut_adj_1784.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_1785 (.I0(t1[0]), .I1(t1[4]), .I2(GND_net), .I3(GND_net), 
            .O(n60014));
    defparam i1_2_lut_adj_1785.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1786 (.I0(t1[2]), .I1(n27655), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5699));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1786.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1787 (.I0(start), .I1(n27611), .I2(GND_net), 
            .I3(GND_net), .O(n27532));
    defparam i1_2_lut_adj_1787.LUT_INIT = 16'h4444;
    SB_LUT4 i2205_2_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));   // verilog/neopixel.v(65[23:32])
    defparam i2205_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1788 (.I0(\bit_ctr[3] ), .I1(n41559), .I2(GND_net), 
            .I3(GND_net), .O(n54679));
    defparam i1_2_lut_adj_1788.LUT_INIT = 16'h6666;
    SB_LUT4 i1176_4_lut (.I0(\color_bit_N_502[1] ), .I1(n41947), .I2(n8_adj_5703), 
            .I3(\color_bit_N_502[2] ), .O(n81));   // verilog/neopixel.v(24[26:38])
    defparam i1176_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i13447_2_lut (.I0(n29957), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n31392));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2226_3_lut (.I0(bit_ctr[4]), .I1(\bit_ctr[3] ), .I2(n7217), 
            .I3(GND_net), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2226_3_lut.LUT_INIT = 16'h6a6a;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1800, ENCODER1_A_N_keep, 
            \a_new[1] , \b_new[1] , n31593, a_prev, n31582, b_prev, 
            n31579, n1805, position_31__N_3836, encoder1_position, GND_net, 
            VCC_net, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1800;
    input ENCODER1_A_N_keep;
    output \a_new[1] ;
    output \b_new[1] ;
    input n31593;
    output a_prev;
    input n31582;
    output b_prev;
    input n31579;
    output n1805;
    output position_31__N_3836;
    output [31:0]encoder1_position;
    input GND_net;
    input VCC_net;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n53396, n53395, n53394, n53393, n53392, 
        n53391, n53390, n53389, n53388, n53387, n53386, n53385, 
        n53384, n53383, n53382, n53381, n53380, n53379, n53378, 
        n53377, n53376, n53375, n53374, n53373, n53372, n53371, 
        n53370, n53369, n53368, n53367, n53366;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1800), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1800), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1800), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1800), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1800), .D(n31593));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1800), .D(n31582));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1805), .C(n1800), .D(n31579));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2042__i0 (.Q(encoder1_position[0]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_2042_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[31]), .I3(n53396), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2042_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[30]), .I3(n53395), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_32 (.CI(n53395), .I0(direction_N_3840), 
            .I1(encoder1_position[30]), .CO(n53396));
    SB_LUT4 position_2042_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[29]), .I3(n53394), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_31 (.CI(n53394), .I0(direction_N_3840), 
            .I1(encoder1_position[29]), .CO(n53395));
    SB_LUT4 position_2042_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[28]), .I3(n53393), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_30 (.CI(n53393), .I0(direction_N_3840), 
            .I1(encoder1_position[28]), .CO(n53394));
    SB_LUT4 position_2042_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[27]), .I3(n53392), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_29 (.CI(n53392), .I0(direction_N_3840), 
            .I1(encoder1_position[27]), .CO(n53393));
    SB_LUT4 position_2042_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[26]), .I3(n53391), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_28 (.CI(n53391), .I0(direction_N_3840), 
            .I1(encoder1_position[26]), .CO(n53392));
    SB_LUT4 position_2042_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[25]), .I3(n53390), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_27 (.CI(n53390), .I0(direction_N_3840), 
            .I1(encoder1_position[25]), .CO(n53391));
    SB_LUT4 position_2042_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[24]), .I3(n53389), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_26 (.CI(n53389), .I0(direction_N_3840), 
            .I1(encoder1_position[24]), .CO(n53390));
    SB_LUT4 position_2042_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[23]), .I3(n53388), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_25 (.CI(n53388), .I0(direction_N_3840), 
            .I1(encoder1_position[23]), .CO(n53389));
    SB_LUT4 position_2042_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[22]), .I3(n53387), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_24 (.CI(n53387), .I0(direction_N_3840), 
            .I1(encoder1_position[22]), .CO(n53388));
    SB_LUT4 position_2042_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[21]), .I3(n53386), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_23 (.CI(n53386), .I0(direction_N_3840), 
            .I1(encoder1_position[21]), .CO(n53387));
    SB_LUT4 position_2042_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[20]), .I3(n53385), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_22 (.CI(n53385), .I0(direction_N_3840), 
            .I1(encoder1_position[20]), .CO(n53386));
    SB_LUT4 position_2042_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[19]), .I3(n53384), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_21 (.CI(n53384), .I0(direction_N_3840), 
            .I1(encoder1_position[19]), .CO(n53385));
    SB_LUT4 position_2042_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[18]), .I3(n53383), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_20 (.CI(n53383), .I0(direction_N_3840), 
            .I1(encoder1_position[18]), .CO(n53384));
    SB_LUT4 position_2042_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[17]), .I3(n53382), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_19 (.CI(n53382), .I0(direction_N_3840), 
            .I1(encoder1_position[17]), .CO(n53383));
    SB_LUT4 position_2042_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[16]), .I3(n53381), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_18 (.CI(n53381), .I0(direction_N_3840), 
            .I1(encoder1_position[16]), .CO(n53382));
    SB_LUT4 position_2042_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[15]), .I3(n53380), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_17 (.CI(n53380), .I0(direction_N_3840), 
            .I1(encoder1_position[15]), .CO(n53381));
    SB_LUT4 position_2042_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[14]), .I3(n53379), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_16 (.CI(n53379), .I0(direction_N_3840), 
            .I1(encoder1_position[14]), .CO(n53380));
    SB_LUT4 position_2042_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[13]), .I3(n53378), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_15 (.CI(n53378), .I0(direction_N_3840), 
            .I1(encoder1_position[13]), .CO(n53379));
    SB_LUT4 position_2042_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[12]), .I3(n53377), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_14 (.CI(n53377), .I0(direction_N_3840), 
            .I1(encoder1_position[12]), .CO(n53378));
    SB_LUT4 position_2042_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[11]), .I3(n53376), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_13 (.CI(n53376), .I0(direction_N_3840), 
            .I1(encoder1_position[11]), .CO(n53377));
    SB_LUT4 position_2042_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[10]), .I3(n53375), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_12 (.CI(n53375), .I0(direction_N_3840), 
            .I1(encoder1_position[10]), .CO(n53376));
    SB_LUT4 position_2042_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[9]), .I3(n53374), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_11 (.CI(n53374), .I0(direction_N_3840), 
            .I1(encoder1_position[9]), .CO(n53375));
    SB_LUT4 position_2042_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[8]), .I3(n53373), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_10 (.CI(n53373), .I0(direction_N_3840), 
            .I1(encoder1_position[8]), .CO(n53374));
    SB_LUT4 position_2042_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[7]), .I3(n53372), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_9 (.CI(n53372), .I0(direction_N_3840), 
            .I1(encoder1_position[7]), .CO(n53373));
    SB_LUT4 position_2042_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[6]), .I3(n53371), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_8 (.CI(n53371), .I0(direction_N_3840), 
            .I1(encoder1_position[6]), .CO(n53372));
    SB_LUT4 position_2042_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[5]), .I3(n53370), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_7 (.CI(n53370), .I0(direction_N_3840), 
            .I1(encoder1_position[5]), .CO(n53371));
    SB_LUT4 position_2042_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[4]), .I3(n53369), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_6 (.CI(n53369), .I0(direction_N_3840), 
            .I1(encoder1_position[4]), .CO(n53370));
    SB_LUT4 position_2042_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[3]), .I3(n53368), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_5 (.CI(n53368), .I0(direction_N_3840), 
            .I1(encoder1_position[3]), .CO(n53369));
    SB_LUT4 position_2042_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[2]), .I3(n53367), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_4 (.CI(n53367), .I0(direction_N_3840), 
            .I1(encoder1_position[2]), .CO(n53368));
    SB_LUT4 position_2042_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[1]), .I3(n53366), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_3 (.CI(n53366), .I0(direction_N_3840), 
            .I1(encoder1_position[1]), .CO(n53367));
    SB_LUT4 position_2042_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2042_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2042_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n53366));
    SB_DFFE position_2042__i1 (.Q(encoder1_position[1]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i2 (.Q(encoder1_position[2]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i3 (.Q(encoder1_position[3]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i4 (.Q(encoder1_position[4]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i5 (.Q(encoder1_position[5]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i6 (.Q(encoder1_position[6]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i7 (.Q(encoder1_position[7]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i8 (.Q(encoder1_position[8]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i9 (.Q(encoder1_position[9]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i10 (.Q(encoder1_position[10]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i11 (.Q(encoder1_position[11]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i12 (.Q(encoder1_position[12]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i13 (.Q(encoder1_position[13]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i14 (.Q(encoder1_position[14]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i15 (.Q(encoder1_position[15]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i16 (.Q(encoder1_position[16]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i17 (.Q(encoder1_position[17]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i18 (.Q(encoder1_position[18]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i19 (.Q(encoder1_position[19]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i20 (.Q(encoder1_position[20]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i21 (.Q(encoder1_position[21]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i22 (.Q(encoder1_position[22]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i23 (.Q(encoder1_position[23]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i24 (.Q(encoder1_position[24]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i25 (.Q(encoder1_position[25]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i26 (.Q(encoder1_position[26]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i27 (.Q(encoder1_position[27]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i28 (.Q(encoder1_position[28]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i29 (.Q(encoder1_position[29]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i30 (.Q(encoder1_position[30]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2042__i31 (.Q(encoder1_position[31]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1800, ENCODER0_A_N_keep, 
            \a_new[1] , \b_new[1] , n1757, GND_net, n1759, n1761, 
            n1763, n1765, n1767, n1769, n1771, n1773, \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , n31592, n1755, 
            n31591, a_prev, n31589, b_prev, \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , VCC_net, position_31__N_3836, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1800;
    input ENCODER0_A_N_keep;
    output \a_new[1] ;
    output \b_new[1] ;
    output n1757;
    input GND_net;
    output n1759;
    output n1761;
    output n1763;
    output n1765;
    output n1767;
    output n1769;
    output n1771;
    output n1773;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    input n31592;
    output n1755;
    input n31591;
    output a_prev;
    input n31589;
    output b_prev;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    output position_31__N_3836;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n53498, n53497, n53496, n53495, n53494, 
        n53493, n53492, n53491, n53490, n53489, n53488, n53487, 
        n53486, n53485, n53484, n53483, n53482, n53481, n53480, 
        n53479, n53478, n53477, n53476, n53475, n53474, n53473, 
        n53472, n53471, n53470, n53469, n53468;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1800), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1800), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1800), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1800), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2055_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1757), .I3(n53498), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2055_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1759), .I3(n53497), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_32 (.CI(n53497), .I0(direction_N_3840), 
            .I1(n1759), .CO(n53498));
    SB_LUT4 position_2055_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1761), .I3(n53496), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_31 (.CI(n53496), .I0(direction_N_3840), 
            .I1(n1761), .CO(n53497));
    SB_LUT4 position_2055_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1763), .I3(n53495), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_30 (.CI(n53495), .I0(direction_N_3840), 
            .I1(n1763), .CO(n53496));
    SB_LUT4 position_2055_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1765), .I3(n53494), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_29 (.CI(n53494), .I0(direction_N_3840), 
            .I1(n1765), .CO(n53495));
    SB_LUT4 position_2055_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1767), .I3(n53493), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_28 (.CI(n53493), .I0(direction_N_3840), 
            .I1(n1767), .CO(n53494));
    SB_LUT4 position_2055_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1769), .I3(n53492), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_27 (.CI(n53492), .I0(direction_N_3840), 
            .I1(n1769), .CO(n53493));
    SB_LUT4 position_2055_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1771), .I3(n53491), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_26 (.CI(n53491), .I0(direction_N_3840), 
            .I1(n1771), .CO(n53492));
    SB_LUT4 position_2055_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1773), .I3(n53490), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_25 (.CI(n53490), .I0(direction_N_3840), 
            .I1(n1773), .CO(n53491));
    SB_LUT4 position_2055_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n53489), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_24 (.CI(n53489), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n53490));
    SB_LUT4 position_2055_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n53488), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_23 (.CI(n53488), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n53489));
    SB_LUT4 position_2055_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n53487), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_22 (.CI(n53487), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n53488));
    SB_LUT4 position_2055_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n53486), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_21 (.CI(n53486), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n53487));
    SB_LUT4 position_2055_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n53485), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_20 (.CI(n53485), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n53486));
    SB_LUT4 position_2055_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n53484), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_19 (.CI(n53484), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n53485));
    SB_LUT4 position_2055_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n53483), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_18 (.CI(n53483), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n53484));
    SB_LUT4 position_2055_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n53482), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_17 (.CI(n53482), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n53483));
    SB_LUT4 position_2055_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n53481), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_16 (.CI(n53481), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n53482));
    SB_LUT4 position_2055_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n53480), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_15 (.CI(n53480), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n53481));
    SB_LUT4 position_2055_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n53479), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_14 (.CI(n53479), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n53480));
    SB_LUT4 position_2055_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n53478), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_13 (.CI(n53478), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n53479));
    SB_LUT4 position_2055_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n53477), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_12 (.CI(n53477), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n53478));
    SB_LUT4 position_2055_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n53476), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_11 (.CI(n53476), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n53477));
    SB_LUT4 position_2055_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n53475), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_10 (.CI(n53475), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n53476));
    SB_LUT4 position_2055_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n53474), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_9 (.CI(n53474), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n53475));
    SB_LUT4 position_2055_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n53473), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_8 (.CI(n53473), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n53474));
    SB_LUT4 position_2055_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n53472), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_7 (.CI(n53472), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n53473));
    SB_DFF direction_42 (.Q(n1755), .C(n1800), .D(n31592));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1800), .D(n31591));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1800), .D(n31589));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2055_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n53471), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_6 (.CI(n53471), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n53472));
    SB_LUT4 position_2055_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n53470), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_5 (.CI(n53470), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n53471));
    SB_LUT4 position_2055_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n53469), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_4 (.CI(n53469), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n53470));
    SB_LUT4 position_2055_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n53468), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_3 (.CI(n53468), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n53469));
    SB_LUT4 position_2055_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2055_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2055_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n53468));
    SB_DFFE position_2055__i0 (.Q(\encoder0_position[0] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i1 (.Q(\encoder0_position[1] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i2 (.Q(\encoder0_position[2] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i3 (.Q(\encoder0_position[3] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i4 (.Q(\encoder0_position[4] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i5 (.Q(\encoder0_position[5] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i6 (.Q(\encoder0_position[6] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i7 (.Q(\encoder0_position[7] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i8 (.Q(\encoder0_position[8] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i9 (.Q(\encoder0_position[9] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i10 (.Q(\encoder0_position[10] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i11 (.Q(\encoder0_position[11] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i12 (.Q(\encoder0_position[12] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i13 (.Q(\encoder0_position[13] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i14 (.Q(\encoder0_position[14] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i15 (.Q(\encoder0_position[15] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i16 (.Q(\encoder0_position[16] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i17 (.Q(\encoder0_position[17] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i18 (.Q(\encoder0_position[18] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i19 (.Q(\encoder0_position[19] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i20 (.Q(\encoder0_position[20] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i21 (.Q(\encoder0_position[21] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i22 (.Q(\encoder0_position[22] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i23 (.Q(n1773), .C(n1800), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i24 (.Q(n1771), .C(n1800), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i25 (.Q(n1769), .C(n1800), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i26 (.Q(n1767), .C(n1800), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i27 (.Q(n1765), .C(n1800), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i28 (.Q(n1763), .C(n1800), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i29 (.Q(n1761), .C(n1800), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i30 (.Q(n1759), .C(n1800), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2055__i31 (.Q(n1757), .C(n1800), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n2889, \data_out_frame[18] , clk16MHz, n59826, \FRAME_MATCHER.state[3] , 
            n60431, GND_net, n31950, VCC_net, \data_in_frame[16] , 
            n59825, n59824, n31947, n59823, n31262, n59770, n59822, 
            \data_out_frame[19] , n59821, n59820, n31257, n59819, 
            n59818, rx_data, \data_out_frame[14] , \data_out_frame[15] , 
            byte_transmit_counter, \data_out_frame[12] , \data_out_frame[13] , 
            n59817, \data_out_frame[20] , \data_out_frame[22] , n31942, 
            n59816, \data_out_frame[0][2] , n59946, \data_out_frame[0][3] , 
            n59945, control_mode, n27629, n51206, \data_out_frame[0][4] , 
            n59944, n31939, n59815, displacement, \encoder0_position_scaled[10] , 
            n54181, n8, \data_out_frame[1][0] , n59943, \data_out_frame[1][1] , 
            n59942, n31936, \data_out_frame[1][3] , n59941, \data_out_frame[17] , 
            \FRAME_MATCHER.i_31__N_2509 , pwm_setpoint, n31251, \data_out_frame[25] , 
            n60434, n54659, LED_c, n59947, n59814, n59813, n59812, 
            n59811, n59810, n59809, \data_out_frame[21] , n59808, 
            n59807, n60592, n59806, n59805, n59804, \data_out_frame[1][5] , 
            n59940, \data_out_frame[1][6] , n59939, n59803, n31237, 
            n10, n152, n30382, \data_out_frame[23] , n28303, n59802, 
            n31933, \data_out_frame[1][7] , n59938, n28963, \data_out_frame[16] , 
            setpoint, \data_out_frame[3][1] , n59937, n27161, \data_out_frame[24] , 
            n31930, \data_out_frame[3][3] , n59936, \data_out_frame[3][4] , 
            n59935, \data_out_frame[3][6] , n59934, n31927, \data_out_frame[3][7] , 
            n59933, \data_out_frame[4] , n59932, n59931, n59930, n55737, 
            n59929, n59928, n59927, n59926, n59925, \data_out_frame[5] , 
            n59924, n59801, n59800, n59799, n59798, n59797, n59796, 
            n59923, n59795, n59922, n59794, n59793, \data_in_frame[3] , 
            \data_in_frame[4] , n59921, n59792, n59791, n59920, n59790, 
            n59789, n59788, n59787, n59786, n59785, n59784, n59919, 
            n59783, \data_in_frame[1] , n59782, n59781, n59780, n61872, 
            n59779, \current[15] , n59778, n59777, n59918, n55561, 
            \current[11] , n31897, \data_in_frame[14] , \current[10] , 
            n59776, n59775, n24, \current[9] , n55706, n23, n25, 
            n59774, n59773, \current[8] , n59772, n59771, n59832, 
            \data_in_frame[5][4] , \data_in_frame[2][1] , n60470, \data_out_frame[6] , 
            \encoder0_position_scaled[16] , n31893, n59917, \data_out_frame[26][1] , 
            \data_out_frame[26][2] , reset, n31890, \data_in_frame[21] , 
            n59916, \data_out_frame[27][1] , \data_out_frame[27][2] , 
            n31887, \data_out_frame[11][7] , \encoder0_position_scaled[7] , 
            \data_out_frame[11][6] , \encoder0_position_scaled[6] , \data_out_frame[11][5] , 
            \encoder0_position_scaled[5] , \data_out_frame[11][4] , \encoder0_position_scaled[4] , 
            \data_out_frame[11][3] , \encoder0_position_scaled[3] , \data_out_frame[11][2] , 
            \encoder0_position_scaled[2] , \data_out_frame[11][1] , \encoder0_position_scaled[1] , 
            \data_in_frame[10] , n59915, \data_out_frame[10] , \encoder0_position_scaled[15] , 
            \encoder0_position_scaled[14] , n59914, \encoder0_position_scaled[13] , 
            \encoder0_position_scaled[12] , \encoder0_position_scaled[11] , 
            n31881, \data_in_frame[14][2] , n31878, \data_in_frame[14][1] , 
            n59913, n31875, \data_in_frame[14][0] , \encoder0_position_scaled[9] , 
            \encoder0_position_scaled[8] , n59912, n59911, \data_in_frame[5][5] , 
            \data_out_frame[9] , \encoder0_position_scaled[23] , \encoder0_position_scaled[22] , 
            \encoder0_position_scaled[21] , \encoder0_position_scaled[20] , 
            \encoder0_position_scaled[19] , n60254, \data_in_frame[20] , 
            \data_in_frame[21][0] , \data_in_frame[18] , \data_in_frame[21][1] , 
            \data_in_frame[21][4] , \data_in_frame[19] , \data_in_frame[21][5] , 
            \data_in_frame[18][1] , \data_in_frame[18][3] , \data_in_frame[18][0] , 
            \data_in_frame[17][5] , \encoder0_position_scaled[18] , \data_in_frame[18][4] , 
            \data_in_frame[12] , \data_in_frame[19][7] , \data_in_frame[17][7] , 
            \encoder0_position_scaled[17] , \data_in_frame[18][2] , \data_in_frame[9] , 
            \data_in_frame[6][3] , n31847, \data_in_frame[6][5] , \data_in_frame[5][0] , 
            n31844, n31841, \data_out_frame[8][7] , \data_in_frame[5][6] , 
            \data_in_frame[5][7] , n31836, n59910, \data_out_frame[8][6] , 
            n31833, n59909, n31830, n31827, n31824, \data_out_frame[8][5] , 
            \data_in_frame[19][2] , \data_in_frame[21][3] , \data_in_frame[17][0] , 
            \data_out_frame[8][4] , \data_in_frame[17][6] , \data_out_frame[8][3] , 
            n31797, n31794, n31791, n31788, n31785, \data_out_frame[8][2] , 
            n31782, \data_out_frame[8][1] , n31779, n31776, n31773, 
            n31770, n31767, \data_out_frame[7] , n59122, \data_in_frame[6][0] , 
            n31557, \data_in_frame[6][1] , n59126, \data_in_frame[6][2] , 
            n59114, n31566, \data_in_frame[6][4] , n59110, n58986, 
            \data_in_frame[6][6] , n59908, n31745, n31742, n31739, 
            n31736, n31733, n59907, \data_in_frame[17][3] , DE_c, 
            \data_in_frame[2][0] , \data_in_frame[17][4] , n59906, n59905, 
            n59904, n59833, n59903, n59902, n59901, n59900, n59899, 
            n59898, n59897, n59896, n59895, n59894, n59893, n59892, 
            n59891, n59890, n59889, n59888, n59887, n59886, n59885, 
            n59884, n59883, n59882, n59881, n59880, n59879, n59878, 
            n32669, n31321, n59877, n59876, n59875, n59874, n59873, 
            n59872, n59871, n59870, n59869, n59868, n59867, n59866, 
            n59865, n59864, n59863, n59862, n59861, n59860, n59859, 
            n59834, n59858, n32691, n31299, n59857, n59856, n59855, 
            n59854, n31294, n59853, n59852, n59851, n59850, n59849, 
            n59848, n59847, n59846, n59845, n32706, n31284, n59844, 
            n59843, n59842, n31590, \FRAME_MATCHER.rx_data_ready_prev , 
            n59841, n59840, n59839, n31277, n59838, n59837, n59836, 
            n59835, n59831, \FRAME_MATCHER.i[0] , n59830, \data_in_frame[2][4] , 
            \data_in_frame[5][1] , \data_in_frame[2][5] , n59829, \data_in_frame[5][2] , 
            ID, \data_in_frame[3][3] , \data_in_frame[1][1] , \data_in_frame[3][0] , 
            \data_in_frame[3][2] , \data_in_frame[1][0] , \data_in_frame[2][2] , 
            deadband, n71521, \data_in_frame[22][4] , \data_in_frame[22][6] , 
            \data_in_frame[22][1] , \data_in_frame[22][0] , \data_in_frame[22][3] , 
            \data_in_frame[22][2] , IntegralLimit, \Kp[0] , \Ki[0] , 
            PWMLimit, n31269, n161, n59828, n31954, n60741, n62047, 
            n31965, n31968, n31971, n31974, n31977, n59150, n59148, 
            n59146, n31990, n59144, n31996, n59142, n59140, n59138, 
            n31440, n59136, n31443, n32066, n31446, n31449, \data_in_frame[2][3] , 
            n32078, n31452, n32088, n31455, n32092, n59062, n32108, 
            n32112, n32115, n32118, n32350, n31482, \Kp[1] , \Kp[2] , 
            \Kp[3] , \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , 
            \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , 
            \Kp[15] , \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , 
            \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , n31488, n32229, 
            neopxl_color, n32228, n32227, n32226, n32225, n32222, 
            n32221, n32220, n32218, n32217, n32216, n32215, n32214, 
            n32213, n32212, n32211, n32210, n32209, n32208, n32207, 
            n32206, current_limit, n31463, n31462, n59827, n32203, 
            n32202, n32201, n32200, n32199, n32197, n32196, n32195, 
            n32193, n32192, n32191, n32190, n32189, n32188, n32187, 
            n32186, n32185, n31491, n31500, n31503, n60669, n167, 
            n28330, n54982, n60241, n54578, n3491, rx_data_ready, 
            n61989, n71389, n71401, n30156, n60391, n1, n144, 
            n163, n60044, n60042, n60039, n67759, n28021, n30370, 
            n10_adj_6, n30449, n70677, n30366, n30416, \current[7] , 
            n24903, \current[6] , \current[5] , n24877, \current[4] , 
            \current[3] , \current[2] , \current[1] , \current[0] , 
            n30414, n30362, n30452, n30447, n62670, n62228, n30368, 
            control_update, n41374, n27538, tx_active, n45, n31, 
            n28, n30, n30423, n60355, n60038, n64880, n64878, 
            n64890, n64891, n64615, n64614, n1_adj_7, tx_o, r_SM_Main, 
            \r_SM_Main_2__N_3536[1] , r_Clock_Count, n29824, \r_Bit_Index[0] , 
            n59688, n31480, n63187, n27, n32074, n71705, n63177, 
            n5235, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , n29, 
            n23_adj_8, n61652, n6, n60832, tx_enable, n31953, baudrate, 
            n31945, n27632, \r_SM_Main[2]_adj_9 , r_Rx_Data, RX_N_2, 
            \o_Rx_DV_N_3488[8] , \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            r_Clock_Count_adj_22, n31702, \r_SM_Main[1]_adj_18 , n29821, 
            r_Bit_Index, n32083, n55814, n32231, n32087, n32021, 
            n32020, n31961, n6_adj_20, n5232, n4, n59686, n63199, 
            \r_SM_Main_2__N_3446[1] , n4_adj_21, n63175, n41584, n29817, 
            n60834) /* synthesis syn_module_defined=1 */ ;
    input n2889;
    output [7:0]\data_out_frame[18] ;
    input clk16MHz;
    input n59826;
    output \FRAME_MATCHER.state[3] ;
    output n60431;
    input GND_net;
    input n31950;
    input VCC_net;
    output [7:0]\data_in_frame[16] ;
    input n59825;
    input n59824;
    input n31947;
    input n59823;
    input n31262;
    input n59770;
    input n59822;
    output [7:0]\data_out_frame[19] ;
    input n59821;
    input n59820;
    input n31257;
    input n59819;
    input n59818;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    input n59817;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[22] ;
    input n31942;
    input n59816;
    output \data_out_frame[0][2] ;
    input n59946;
    output \data_out_frame[0][3] ;
    input n59945;
    output [7:0]control_mode;
    input n27629;
    output n51206;
    output \data_out_frame[0][4] ;
    input n59944;
    input n31939;
    input n59815;
    input [23:0]displacement;
    input \encoder0_position_scaled[10] ;
    input n54181;
    output n8;
    output \data_out_frame[1][0] ;
    input n59943;
    output \data_out_frame[1][1] ;
    input n59942;
    input n31936;
    output \data_out_frame[1][3] ;
    input n59941;
    output [7:0]\data_out_frame[17] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]pwm_setpoint;
    input n31251;
    output [7:0]\data_out_frame[25] ;
    output n60434;
    output n54659;
    output LED_c;
    input n59947;
    input n59814;
    input n59813;
    input n59812;
    input n59811;
    input n59810;
    input n59809;
    output [7:0]\data_out_frame[21] ;
    input n59808;
    input n59807;
    output n60592;
    input n59806;
    input n59805;
    input n59804;
    output \data_out_frame[1][5] ;
    input n59940;
    output \data_out_frame[1][6] ;
    input n59939;
    input n59803;
    input n31237;
    output n10;
    input n152;
    output n30382;
    output [7:0]\data_out_frame[23] ;
    output n28303;
    input n59802;
    input n31933;
    output \data_out_frame[1][7] ;
    input n59938;
    output n28963;
    output [7:0]\data_out_frame[16] ;
    output [23:0]setpoint;
    output \data_out_frame[3][1] ;
    input n59937;
    input n27161;
    output [7:0]\data_out_frame[24] ;
    input n31930;
    output \data_out_frame[3][3] ;
    input n59936;
    output \data_out_frame[3][4] ;
    input n59935;
    output \data_out_frame[3][6] ;
    input n59934;
    input n31927;
    output \data_out_frame[3][7] ;
    input n59933;
    output [7:0]\data_out_frame[4] ;
    input n59932;
    input n59931;
    input n59930;
    input n55737;
    input n59929;
    input n59928;
    input n59927;
    input n59926;
    input n59925;
    output [7:0]\data_out_frame[5] ;
    input n59924;
    input n59801;
    input n59800;
    input n59799;
    input n59798;
    input n59797;
    input n59796;
    input n59923;
    input n59795;
    input n59922;
    input n59794;
    input n59793;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[4] ;
    input n59921;
    input n59792;
    input n59791;
    input n59920;
    input n59790;
    input n59789;
    input n59788;
    input n59787;
    input n59786;
    input n59785;
    input n59784;
    input n59919;
    input n59783;
    output [7:0]\data_in_frame[1] ;
    input n59782;
    input n59781;
    input n59780;
    output n61872;
    input n59779;
    input \current[15] ;
    input n59778;
    input n59777;
    input n59918;
    output n55561;
    input \current[11] ;
    input n31897;
    output [7:0]\data_in_frame[14] ;
    input \current[10] ;
    input n59776;
    input n59775;
    output n24;
    input \current[9] ;
    output n55706;
    output n23;
    output n25;
    input n59774;
    input n59773;
    input \current[8] ;
    input n59772;
    input n59771;
    input n59832;
    output \data_in_frame[5][4] ;
    output \data_in_frame[2][1] ;
    output n60470;
    output [7:0]\data_out_frame[6] ;
    input \encoder0_position_scaled[16] ;
    input n31893;
    input n59917;
    output \data_out_frame[26][1] ;
    output \data_out_frame[26][2] ;
    input reset;
    input n31890;
    output [7:0]\data_in_frame[21] ;
    input n59916;
    output \data_out_frame[27][1] ;
    output \data_out_frame[27][2] ;
    input n31887;
    output \data_out_frame[11][7] ;
    input \encoder0_position_scaled[7] ;
    output \data_out_frame[11][6] ;
    input \encoder0_position_scaled[6] ;
    output \data_out_frame[11][5] ;
    input \encoder0_position_scaled[5] ;
    output \data_out_frame[11][4] ;
    input \encoder0_position_scaled[4] ;
    output \data_out_frame[11][3] ;
    input \encoder0_position_scaled[3] ;
    output \data_out_frame[11][2] ;
    input \encoder0_position_scaled[2] ;
    output \data_out_frame[11][1] ;
    input \encoder0_position_scaled[1] ;
    output [7:0]\data_in_frame[10] ;
    input n59915;
    output [7:0]\data_out_frame[10] ;
    input \encoder0_position_scaled[15] ;
    input \encoder0_position_scaled[14] ;
    input n59914;
    input \encoder0_position_scaled[13] ;
    input \encoder0_position_scaled[12] ;
    input \encoder0_position_scaled[11] ;
    input n31881;
    output \data_in_frame[14][2] ;
    input n31878;
    output \data_in_frame[14][1] ;
    input n59913;
    input n31875;
    output \data_in_frame[14][0] ;
    input \encoder0_position_scaled[9] ;
    input \encoder0_position_scaled[8] ;
    input n59912;
    input n59911;
    output \data_in_frame[5][5] ;
    output [7:0]\data_out_frame[9] ;
    input \encoder0_position_scaled[23] ;
    input \encoder0_position_scaled[22] ;
    input \encoder0_position_scaled[21] ;
    input \encoder0_position_scaled[20] ;
    input \encoder0_position_scaled[19] ;
    input n60254;
    output [7:0]\data_in_frame[20] ;
    output \data_in_frame[21][0] ;
    output [7:0]\data_in_frame[18] ;
    output \data_in_frame[21][1] ;
    output \data_in_frame[21][4] ;
    output [7:0]\data_in_frame[19] ;
    output \data_in_frame[21][5] ;
    output \data_in_frame[18][1] ;
    output \data_in_frame[18][3] ;
    output \data_in_frame[18][0] ;
    output \data_in_frame[17][5] ;
    input \encoder0_position_scaled[18] ;
    output \data_in_frame[18][4] ;
    output [7:0]\data_in_frame[12] ;
    output \data_in_frame[19][7] ;
    output \data_in_frame[17][7] ;
    input \encoder0_position_scaled[17] ;
    output \data_in_frame[18][2] ;
    output [7:0]\data_in_frame[9] ;
    output \data_in_frame[6][3] ;
    input n31847;
    output \data_in_frame[6][5] ;
    output \data_in_frame[5][0] ;
    input n31844;
    input n31841;
    output \data_out_frame[8][7] ;
    output \data_in_frame[5][6] ;
    output \data_in_frame[5][7] ;
    input n31836;
    input n59910;
    output \data_out_frame[8][6] ;
    input n31833;
    input n59909;
    input n31830;
    input n31827;
    input n31824;
    output \data_out_frame[8][5] ;
    output \data_in_frame[19][2] ;
    output \data_in_frame[21][3] ;
    output \data_in_frame[17][0] ;
    output \data_out_frame[8][4] ;
    output \data_in_frame[17][6] ;
    output \data_out_frame[8][3] ;
    input n31797;
    input n31794;
    input n31791;
    input n31788;
    input n31785;
    output \data_out_frame[8][2] ;
    input n31782;
    output \data_out_frame[8][1] ;
    input n31779;
    input n31776;
    input n31773;
    input n31770;
    input n31767;
    output [7:0]\data_out_frame[7] ;
    input n59122;
    output \data_in_frame[6][0] ;
    input n31557;
    output \data_in_frame[6][1] ;
    input n59126;
    output \data_in_frame[6][2] ;
    input n59114;
    input n31566;
    output \data_in_frame[6][4] ;
    input n59110;
    input n58986;
    output \data_in_frame[6][6] ;
    input n59908;
    input n31745;
    input n31742;
    input n31739;
    input n31736;
    input n31733;
    input n59907;
    output \data_in_frame[17][3] ;
    output DE_c;
    output \data_in_frame[2][0] ;
    output \data_in_frame[17][4] ;
    input n59906;
    input n59905;
    input n59904;
    input n59833;
    input n59903;
    input n59902;
    input n59901;
    input n59900;
    input n59899;
    input n59898;
    input n59897;
    input n59896;
    input n59895;
    input n59894;
    input n59893;
    input n59892;
    input n59891;
    input n59890;
    input n59889;
    input n59888;
    input n59887;
    input n59886;
    input n59885;
    input n59884;
    input n59883;
    input n59882;
    input n59881;
    input n59880;
    input n59879;
    input n59878;
    input n32669;
    input n31321;
    input n59877;
    input n59876;
    input n59875;
    input n59874;
    input n59873;
    input n59872;
    input n59871;
    input n59870;
    input n59869;
    input n59868;
    input n59867;
    input n59866;
    input n59865;
    input n59864;
    input n59863;
    input n59862;
    input n59861;
    input n59860;
    input n59859;
    input n59834;
    input n59858;
    input n32691;
    input n31299;
    input n59857;
    input n59856;
    input n59855;
    input n59854;
    input n31294;
    input n59853;
    input n59852;
    input n59851;
    input n59850;
    input n59849;
    input n59848;
    input n59847;
    input n59846;
    input n59845;
    input n32706;
    input n31284;
    input n59844;
    input n59843;
    input n59842;
    input n31590;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n59841;
    input n59840;
    input n59839;
    input n31277;
    input n59838;
    input n59837;
    input n59836;
    input n59835;
    input n59831;
    output \FRAME_MATCHER.i[0] ;
    input n59830;
    output \data_in_frame[2][4] ;
    output \data_in_frame[5][1] ;
    output \data_in_frame[2][5] ;
    input n59829;
    output \data_in_frame[5][2] ;
    input [7:0]ID;
    output \data_in_frame[3][3] ;
    output \data_in_frame[1][1] ;
    output \data_in_frame[3][0] ;
    output \data_in_frame[3][2] ;
    output \data_in_frame[1][0] ;
    output \data_in_frame[2][2] ;
    output [23:0]deadband;
    output n71521;
    output \data_in_frame[22][4] ;
    output \data_in_frame[22][6] ;
    output \data_in_frame[22][1] ;
    output \data_in_frame[22][0] ;
    output \data_in_frame[22][3] ;
    output \data_in_frame[22][2] ;
    output [23:0]IntegralLimit;
    output \Kp[0] ;
    output \Ki[0] ;
    output [23:0]PWMLimit;
    input n31269;
    output n161;
    input n59828;
    input n31954;
    input n60741;
    output n62047;
    input n31965;
    input n31968;
    input n31971;
    input n31974;
    input n31977;
    input n59150;
    input n59148;
    input n59146;
    input n31990;
    input n59144;
    input n31996;
    input n59142;
    input n59140;
    input n59138;
    input n31440;
    input n59136;
    input n31443;
    input n32066;
    input n31446;
    input n31449;
    output \data_in_frame[2][3] ;
    input n32078;
    input n31452;
    input n32088;
    input n31455;
    input n32092;
    input n59062;
    input n32108;
    input n32112;
    input n32115;
    input n32118;
    input n32350;
    input n31482;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    output \Kp[13] ;
    output \Kp[14] ;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    input n31488;
    input n32229;
    output [23:0]neopxl_color;
    input n32228;
    input n32227;
    input n32226;
    input n32225;
    input n32222;
    input n32221;
    input n32220;
    input n32218;
    input n32217;
    input n32216;
    input n32215;
    input n32214;
    input n32213;
    input n32212;
    input n32211;
    input n32210;
    input n32209;
    input n32208;
    input n32207;
    input n32206;
    output [15:0]current_limit;
    input n31463;
    input n31462;
    input n59827;
    input n32203;
    input n32202;
    input n32201;
    input n32200;
    input n32199;
    input n32197;
    input n32196;
    input n32195;
    input n32193;
    input n32192;
    input n32191;
    input n32190;
    input n32189;
    input n32188;
    input n32187;
    input n32186;
    input n32185;
    input n31491;
    input n31500;
    input n31503;
    output n60669;
    output n167;
    input n28330;
    input n54982;
    input n60241;
    output n54578;
    output n3491;
    output rx_data_ready;
    output n61989;
    input n71389;
    input n71401;
    output n30156;
    output n60391;
    output n1;
    output n144;
    output n163;
    input n60044;
    output n60042;
    output n60039;
    input n67759;
    output n28021;
    input n30370;
    output n10_adj_6;
    output n30449;
    input n70677;
    output n30366;
    output n30416;
    input \current[7] ;
    output n24903;
    input \current[6] ;
    input \current[5] ;
    output n24877;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    output n30414;
    output n30362;
    output n30452;
    output n30447;
    output n62670;
    output n62228;
    output n30368;
    input control_update;
    input n41374;
    output n27538;
    output tx_active;
    output n45;
    output n31;
    input n28;
    output n30;
    input n30423;
    input n60355;
    output n60038;
    input n64880;
    input n64878;
    input n64890;
    input n64891;
    input n64615;
    input n64614;
    output n1_adj_7;
    output tx_o;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    output [8:0]r_Clock_Count;
    output n29824;
    output \r_Bit_Index[0] ;
    output n59688;
    input n31480;
    input n63187;
    output n27;
    input n32074;
    input n71705;
    output n63177;
    input n5235;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23_adj_8;
    input n61652;
    output n6;
    output n60832;
    output tx_enable;
    input n31953;
    input [31:0]baudrate;
    input n31945;
    output n27632;
    output \r_SM_Main[2]_adj_9 ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output [7:0]r_Clock_Count_adj_22;
    input n31702;
    output \r_SM_Main[1]_adj_18 ;
    output n29821;
    output [2:0]r_Bit_Index;
    input n32083;
    input n55814;
    input n32231;
    input n32087;
    input n32021;
    input n32020;
    input n31961;
    output n6_adj_20;
    input n5232;
    output n4;
    output n59686;
    input n63199;
    input \r_SM_Main_2__N_3446[1] ;
    output n4_adj_21;
    output n63175;
    output n41584;
    output n29817;
    output n60834;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2, n55784, n3, n2_adj_5291, n2_adj_5292, n2_adj_5293, 
        n2_adj_5294, n2_adj_5295, n31539;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5296, n2_adj_5297, n2_adj_5298, n2_adj_5299, n2_adj_5300, 
        n2_adj_5301, n8_c, n60036;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n31866, n31869, n64588, n64587, n2_adj_5302, n31872, n54636, 
        n55690, n62640, n5, n60437, n61755, n3_adj_5303, n2_adj_5304, 
        n2_adj_5305, n55641, n55627, n2_adj_5306, n60634, n60635, 
        n2_adj_5307, n2_adj_5308, n2_adj_5310, n2_adj_5311, n2_adj_5312, 
        n28889, n60775;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5313, n60381, n6_c, n2_adj_5314, n62178, n3_adj_5315, 
        n2_adj_5316, n55008, n3_adj_5317, n60322, n60695, LED_N_3408, 
        LED_N_3407, n27913, n55659, n55663, n2_adj_5318, n29481, 
        \FRAME_MATCHER.i_31__N_2513 , n31050, n3_adj_5319, Kp_23__N_1748, 
        Kp_23__N_612, n5_adj_5320, n2_adj_5321, n2_adj_5322, n2_adj_5323, 
        n2_adj_5324, n2_adj_5325, n2_adj_5326, n2_adj_5327, n2_adj_5328, 
        n2_adj_5329, n60227, n54689, n2_adj_5330, n2_adj_5331, n2_adj_5332, 
        n55665, n60359, n8_adj_5333, n2_adj_5334, n2_adj_5335, n8_adj_5336, 
        n3_adj_5337, n2_adj_5338, n2_adj_5339, n2_adj_5340, n2_adj_5341, 
        n2_adj_5342, n2_adj_5343, n60440, n55546, n3_adj_5344, n60689, 
        n55645, n18, n60449, n20, n60692, n16, n60672, n55719, 
        n62514, n16_adj_5345, n2_adj_5346, n2_adj_5347, n2_adj_5348, 
        n28864, n60452, n60756, n16_adj_5349, n15, n60362, n60797, 
        n28869, n17, n54936, n18_adj_5350, n2_adj_5351, n60076, 
        n20_adj_5352, n55770, n2_adj_5353, n6_adj_5354, n2_adj_5355, 
        n2_adj_5356, n2_adj_5357, n2_adj_5358, n2_adj_5359, n2_adj_5360, 
        n2_adj_5361, n2_adj_5362, n31924;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5363, n12, n31921, n2_adj_5364, n2_adj_5365, n31918, 
        n2_adj_5366, n31915, n2_adj_5367, n31912, n2_adj_5368, n31909, 
        n2_adj_5369, n2_adj_5370, n2_adj_5371, n2_adj_5372, n2_adj_5373, 
        n2_adj_5374, n2_adj_5375, n2_adj_5376, n2_adj_5377, n2_adj_5378, 
        n2_adj_5379, n2_adj_5380, n60142, n60331, Kp_23__N_872, n2_adj_5381, 
        n2_adj_5382, n2_adj_5383, n31903, n2_adj_5384, n2_adj_5385, 
        n2_adj_5386, n2_adj_5387, n2_adj_5388, n2_adj_5389, n2_adj_5390, 
        n2_adj_5391, n2_adj_5392, n2_adj_5393, n31900, n2_adj_5394, 
        n2_adj_5395, n3_adj_5396, n2_adj_5397, n60545, n60073, n2_adj_5398, 
        n2_adj_5399, n2_adj_5400, n3_adj_5401, n2_adj_5402, n2_adj_5403, 
        n2_adj_5404, n2_adj_5405, n2_adj_5406, n55776, n60794, n60478, 
        n14, n2_adj_5407, n9, n28608, n13, n2_adj_5408, n2_adj_5409, 
        n2_adj_5410, n2_adj_5411, n60643, n54606, n22, n2_adj_5412, 
        n60424, n55550, n54695, n2_adj_5413, n2_adj_5414, n2_adj_5415, 
        n2_adj_5416, n2_adj_5417, n2_adj_5418, n2_adj_5419, n2_adj_5420, 
        n2_adj_5421, n31542, n2_adj_5422, n6_adj_5423, n3_adj_5424, 
        n3_adj_5425;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n59968;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    
    wire n60272, Kp_23__N_748, n16_adj_5426, n60337, n55542, n60416, 
        n62335, n60548, n60115, n28027, n3_adj_5427, n2_adj_5428, 
        n2_adj_5429, n60487, n3_adj_5430, n2_adj_5431, n2_adj_5432, 
        n3_adj_5433, n59967, n10_adj_5434, Kp_23__N_869, n3_adj_5435, 
        n59966, n2081;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n71380, n28432, n60296, n36324;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    
    wire n7;
    wire [23:0]n4947;
    
    wire n29831, n2_adj_5436, n55186, n55565, n3_adj_5437, n59965;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    
    wire n27900, n60584, n60723, n60562, n28386, n3_adj_5438, n59964, 
        n2_adj_5439, n59962, n55653, n60150, n6_adj_5440, n59963, 
        n2_adj_5441, n59970, n59956, n71383, n59961, n62393;
    wire [7:0]\data_in_frame[21]_c ;   // verilog/coms.v(99[12:25])
    
    wire n8_adj_5442, n59957, n59958, n2_adj_5443, n2_adj_5444, n2_adj_5445, 
        n59955, n59959, n2_adj_5446, n2_adj_5447, n2_adj_5448, n2_adj_5449, 
        n59960, n71374, n2_adj_5450, n2_adj_5451, n28529, n4_c, 
        n28134, n59969, n1_c, n59759, n2_adj_5452, n1_adj_5453, 
        n59760, n1_adj_5454;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n59762, n60607, n60309, n64019, n2_adj_5455, n31886;
    wire [7:0]\data_in_frame[14]_c ;   // verilog/coms.v(99[12:25])
    
    wire n64915, n64914, n71377, n2_adj_5456, n2_adj_5457, n2_adj_5458, 
        n71368, n2_adj_5459, n1_adj_5460, n59763, n2_adj_5461, n1_adj_5462, 
        n59764, n28055, n28074;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    
    wire n64173, n71371, n1_adj_5463, n59761, n2_adj_5464, n2_adj_5465, 
        n2_adj_5466;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n7_adj_5467, n2_adj_5468, n2_adj_5469, n2_adj_5470, n31545, 
        n1_adj_5471, n59765, n31862, n2_adj_5472, n31859, n2_adj_5473, 
        Kp_23__N_1389, n4_adj_5474, n2_adj_5475, n2_adj_5476, n2_adj_5477, 
        n2_adj_5478, n60659, n64167, n55739, n64584, n64585, n71362, 
        n25812, n60763, n28877, n64037, n27332, n60601, n60248, 
        n55671, n6_adj_5479, n55778, n54264, n60306, n60260, n55708, 
        n64213, n60604, n64219, n60540, n60495, n60656, n64225, 
        n60800;
    wire [7:0]\data_in_frame[18]_c ;   // verilog/coms.v(99[12:25])
    
    wire n60579, n64229, n54773, n60765, n60275, n64235, n55766, 
        n60458, n64241, n61855, n62783, n60388, n62602, n60443, 
        n54740;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n28247, n26003, n28753, n28002, n28507, n60278, n64882, 
        n64881, n71365, n54742, n54649, n60785, n64011, n60759, 
        n60701, n8_adj_5480, n60190, n6_adj_5481, n60368, n64003, 
        n60698, n60662, n55643, n62107, n54647, n64057, n64005, 
        n64061, n60817, n28908, n60461, n64081, n55556, n64089, 
        n10_adj_5482, n60473, n61729, n14_adj_5483, n9_adj_5484, n61984, 
        n60682, n2_adj_5485, n60512, n54563, n60374, n55712, n62306, 
        n62554, n27873, n2_adj_5486, n31856, n31853, n54662, n60622, 
        n60396;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    
    wire n12_adj_5487, n60319, n27223, n27843, n60791, n10_adj_5488, 
        n27865, n60508, n10_adj_5489, n2_adj_5490, n60619, n27294, 
        n60132, n28126, n54620, n27810, n60312, n28559, n20_adj_5491, 
        n60094, n19, n60105, n21, n31850, n62103, Kp_23__N_1271, 
        n6_adj_5492, n2_adj_5493, n60484, n26, n54872, n55163, n60428, 
        n16_adj_5494, n28572, n60176, n24_adj_5495, n20_adj_5496, 
        n28_c, Kp_23__N_1080, Kp_23__N_875, n28_adj_5497, n60726, 
        n60287, n54597, n26_adj_5498, n60467, n60217, n27_c, n54746, 
        n60208, n25_adj_5499, n27251, n2_adj_5500, n31548, n31551, 
        n2_adj_5501, \FRAME_MATCHER.i_31__N_2511 , n1_adj_5502, n31821, 
        n2_adj_5503, n6_adj_5504, n60235, n31818, n27264, n12_adj_5505, 
        n54624, n60518, n31815, n54626, n60649, n28583, n31812, 
        n31809, n2_adj_5506, n6_adj_5507, n60224, n60481, n2_adj_5508, 
        n31806, n31803, n31800, n2_adj_5509, n64187, n2_adj_5510, 
        n55482, n60646, n26045, n26041, n2_adj_5511, n60806, n60167, 
        n64067, Kp_23__N_1067, n55710, n60051, n70909, n64195, n64197, 
        n60559, n64203, n64073, n64647, n64648, n71350, n64717, 
        n64716, n71353, n2_adj_5512, n60720, n64209, n31576, n60102, 
        n60769, n31583;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n31586, n31625, n2_adj_5513, n60135, n12_adj_5514, n24_adj_5515, 
        n58710, n60613, n10_adj_5516, n54602, n28834, n71700, \FRAME_MATCHER.i_31__N_2507 , 
        n29158, \FRAME_MATCHER.i_31__N_2508 , n2061, n2062, n23276, 
        n58832, \FRAME_MATCHER.i_31__N_2512 , n2073, n29161, \FRAME_MATCHER.i_31__N_2514 , 
        n54857, n2_adj_5517, n31730, n31727, n2_adj_5518, n62185, 
        n31724, n60220, n28041, n31721, n31718, n31715, n31712, 
        n52659, n59757, n52658, n55574, n60772, n31709, n2_adj_5519, 
        n31688, n60738, n64179, n31705, n31691, n2_adj_5520, n31694, 
        n60524, n27956, n12_adj_5521, n31697, n28366, n52657, Kp_23__N_1085, 
        n60587, n52656, Kp_23__N_974, n28398, n60284, n60293, n27971, 
        n60631, n28490, n27992, n2_adj_5522, n64638, n64639, n71332, 
        n60251, n64624, n64623, n71335, n52655, n29032, n31014, 
        n7_adj_5523, n64025, n27211, n52654, n28463, n52653, n59758, 
        tx_transmit_N_3416, n8_adj_5524, n61746, n55599, n31624;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n31623, n31622, n31621, n31620, n31619, n31618, n31617;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n31616, n31615, n31614, n31613, n31612, n31611, n31610, 
        n31609;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n31608, n31607, n31606, n31605, n31604, n31603, n2_adj_5525, 
        n31602, n31601;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n31600, n31599, n31598, n31597, n2_adj_5526, n31596, n31595, 
        n31594, n2_adj_5527, n2_adj_5528, n2_adj_5529, n2_adj_5530, 
        n2_adj_5531, n2_adj_5532, n2_adj_5533, n2_adj_5534, n2_adj_5535, 
        n2_adj_5536, n64896, n64897, n71326, n1_adj_5537;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n31004, n28435, n60576, n30058, n28296, n60173, n6_adj_5538, 
        n60111, n2_adj_5539;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n60122, n28018, n64603, n64602, n71329, n28006, n14_adj_5540, 
        n60079, n15_adj_5541, n2_adj_5542, n28694, n60365, n10_adj_5543, 
        n11, n12_adj_5544, n71320, n27849, n28009, n12_adj_5545, 
        n10_adj_5546, n11_adj_5547, n9_adj_5548, n62747;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3]_c ;   // verilog/coms.v(99[12:25])
    
    wire n60202, n71518, n28930, n6_adj_5549, n27996, Kp_23__N_799, 
        n64047, Kp_23__N_767, n14_adj_5550, n10_adj_5551, n60199, 
        n67645, n67644, n71323, n28429, Kp_23__N_753, n30148, n30361, 
        n53427, n67576, n64125, n30146, n53426, n67577, n30144, 
        n53425, n67579, n64129, n64133, n30142, n53424, n67580, 
        n30140, n53423, n67581, n64147, n64139, n64151, n64157, 
        n60750, n30138, n53422, n67588, n60747, n15_adj_5552, n14_adj_5553, 
        n62486, n21_adj_5554, n27_adj_5555, n26_adj_5556, n64318, 
        n64467, n30136, n53421, n67591, n30134, n53420, n67592, 
        n31458, n31_c, n7_adj_5557, n8_adj_5558;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n62764;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n64331, n30132, n53419, n67595, n30130, n53418, n67596, 
        n30128, n53417, n67601, n64093, n62652, n62789, n64099, 
        n60257, n10_adj_5559, n30126, n53416, n67602, n30124, n53415, 
        n67646, n64101, n30122, n53414, n67647, n64103, n8_adj_5560, 
        n64105, n12_adj_5561, n64249, n10_adj_5562, n30120, n53413, 
        n67648, n30118, n53412, n67649, n12_adj_5563, n64107, n60735, 
        n62338, n62155, n62150, n64113, n62272, n30116, n53411, 
        n67650, n30114, n53410, n67651, n64115, n71512, n64185, 
        n64119, n31459, n31460, n31461, n30112, n53409, n67659, 
        n30110, n53408, n67671, n71515, n32162, n32163, n32164, 
        n2_adj_5564, n30108, n53407, n67672, n44, n32165, n42, 
        n30106, n53406, n67673, n30104, n53405, n67676, n43, n41, 
        n40, n30102, n53404, n67677, n39, n69670, n67758, n71506, 
        n71437;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n69637, n67745, n71500, n71431, n71494, n71497, n30100, 
        n53403, n67678, n71482, n71485, n71476, n30098, n53402, 
        n67679, n30096, n53401, n67682, n30094, n53400, n67683, 
        n50, n30092, n53399, n67689, n30090, n53398, n67690, n30088, 
        n53397, n67691;
    wire [31:0]n133;
    
    wire n45_c, n6_adj_5565, n60011, n32166, n27621, n4452, n71479, 
        n32167, n71314, n71317, n31478, n32168, n2_adj_5566, n32169, 
        n60782, n8_adj_5567, n54653, n32170, n32171, n32172, n55280, 
        n32173, n54618, n7_adj_5568, n55614, n55544, n55570, n14_adj_5569, 
        n62106, n15_adj_5570, n31957, n31962, n31426, n31429, n59064, 
        n31433, n31437, n59106, n32437, n32435, n59052, n59118, 
        n32038, n32427, n59316, n59308, n32418, n32415, n32412, 
        n32409, n54771, n32406, n32403, n32400, n32397, n32041, 
        n59322, n32048, n32051, n59214, n32059, n32062, n59050, 
        n59046, n59058, n32098, n59060, n32351, n32349, n32130, 
        n32133, n59220, n32140, n32143, n32146, n32149, n59230, 
        n31467, n32334, n31485, n32307, n32306, n32305, n32304, 
        n32303, n32302, n32301, n32300, n32299, n32298, n32297, 
        n32296, n32295, n32294, n32293, n32292, n32291, n32290, 
        n32289, n32288, n32287, n32286, n32285, n32284, n32283, 
        n32282, n32281, n32280, n32279, n32278, n32277, n32276, 
        n32275, n32274, n32273, n32272, n32271, n32270, n32269, 
        n32268, n32267, n32266, n32265, n32264, n32263, n32262, 
        n32261, n32260, n32259, n32258, n32257, n32256, n32255, 
        n32254, n32253, n32252, n32251, n32250, n32249, n32248, 
        n32247, n32246, n32245, n32244, n32243, n32242, n32241, 
        n32240, n32239, n32238, n32237, n32236, n32235, n32234, 
        n32233, n32232, n32224, n32223, n32219, n32205, n32204, 
        n31465, n71173, n67746, n71470, n31464, n2_adj_5571, n32198, 
        n32194, n32184, n32183, n32182, n32181, n32180, n32179, 
        n32178, n32177, n32176, n32175, n32174, n59294, n59298, 
        n55554, n31506, n28707, n60032, n59304, n62354, n60185, 
        n27799, n31512, n62117, n31515, n31518, n31521, n31524, 
        n31527, n31530, n31533, n31536, n60625, n60182, n60717, 
        n10_adj_5572, n60230, n5_adj_5573, n60345, n54752, n40_adj_5574, 
        n60281, n38, n39_adj_5575, n60637, n60054, n37, n60342, 
        n42_adj_5576, n46, n55303, n60145, n41_adj_5577, n60679, 
        n60446, n13_adj_5578, n11_adj_5579, n6_adj_5580, n60325, n60729, 
        n7_adj_5581, n60595, n6_adj_5582, n60568, n64308, n54638, 
        n60410, n55105, n60352, n10_adj_5583, n60349, n37_adj_5584, 
        n28169, n60290, n54789, n60640, n60161, n28198, n18_adj_5585, 
        n27770, n16_adj_5586, n20_adj_5587, n60753, n45_adj_5588, 
        n20_adj_5589, n55703, n1130, n6_adj_5590, n28188, n60565, 
        n60328, n12_adj_5591, n60244, n1835, n7_adj_5592, n8_adj_5593, 
        n55625, n6_adj_5594, n60464, n12_adj_5595, n8_adj_5596, n60002, 
        n39975, n60616, n60268, n12_adj_5597, n60515, n60211, n64887, 
        n54585, n60153, n60490, n64888, n64909, n64908, n60521, 
        n60809, n10_adj_5598, n60066, n6_adj_5599, n27774, n60530, 
        n64722, n64723, n60711, n28524, n28620, n12_adj_5600, n64621, 
        n64620, n64698, n64699, n64711, n64710, n62456, n62385, 
        n64605, n61660, n28347, n12_adj_5601, n64606, n64618, n55167, 
        n64617, n64911, n64912, n64903, n27767, n60170, n60705, 
        n1191, n60708, n10_adj_5602, n64902, n27907, n1516, n60533, 
        n28205, n67616, n67617, n5_adj_5603, n4_adj_5604, n64590, 
        n64591, n60385, n64900, n64899, n1_adj_5605, n67615, n5_adj_5606, 
        n4_adj_5607, n30071, n64870, n64871, n64869, n67755, n67741, 
        n64663, n64664, n64662, n6_adj_5608, n67743, n64705, n64706, 
        n64704, n67730, n30026, n64681, n64682, n64680, n67742, 
        n30024, n64678, n64679, n64677, n14_adj_5609, n28714, n8_adj_5610, 
        n60139, n1655, n60573, n38_adj_5611, n60196, n28918, n45_adj_5612, 
        n60598, n60744, n42_adj_5613, n60062, n60108, n44_adj_5615, 
        n50_adj_5616, n10_adj_5617, n67722, n40004, n48, n32, n1182, 
        n49, n47, n60788, n60156, n15_adj_5618, n14_adj_5619, n60553, 
        n6_adj_5620, n28769, n60214, n28445, n27763, n6_adj_5621, 
        n60316, n60082, n60125, n60556, n12_adj_5622, n12_adj_5623, 
        n60714, n62204, n60778, n6_adj_5624, n60610, n10_adj_5625, 
        n60812, n28_adj_5626, n29000, n38_adj_5627, n36, n42_adj_5628, 
        n40_adj_5629, n60675, n60048, n41_adj_5630, n39_adj_5631, 
        n62609, n10_adj_5632, n30400, n60527, n6_adj_5633, n60455, 
        n10_adj_5634, n60164, n6_adj_5635, n71179, n71464, n10_adj_5636, 
        n8_adj_5637, n771, n27595, n4_adj_5638, n40142, n6_adj_5640, 
        n8_adj_5641, n8_adj_5642, n86, n64302, n4_adj_5643, n80, 
        n60026, n60017, n30380, n7_adj_5644, n71407, n71185, n71458, 
        n7_adj_5645, n30390, n1964, n61882, n23271, n24814, n3303, 
        n1967, n1970, n64276, n62294, n1968, n6_adj_5646, n27491, 
        n71191, n71452, n7_adj_5647, n71197, n71446, n96, n39989, 
        n40019, n29711, n61670, n27610, n10_adj_5648, n4_adj_5649, 
        n14_adj_5650, n27634, n27521, n20_adj_5651, n19_adj_5652, 
        n7_adj_5653, n64483, n27684, n18_adj_5654, n27658, n20_adj_5655, 
        n71203, n71440, n71305, n7_adj_5656, n15_adj_5657, n71434, 
        n4_adj_5658, n53, n40172, n40157, n10_adj_5659, n14_adj_5660, 
        n15_adj_5661, n71302, n16_adj_5662, n17_adj_5663, n16_adj_5664, 
        n71413, n71299, n71419, n17_adj_5665, n15_adj_5666, n16_adj_5667, 
        n71428, n71296, n4_adj_5668, n4_adj_5669, n41899, n5_adj_5670, 
        n62599, n7_adj_5674, n71416, n71410, n71404, n10_adj_5675, 
        n26037, n22_adj_5676, n20_adj_5677, n24_adj_5678, n6_adj_5679, 
        n71200, n71194, n71188, n71182, n71176, n71170;
    
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2), .S(n59826));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_223_i3_3_lut (.I0(n55784), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60431), .I3(GND_net), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_223_i3_3_lut.LUT_INIT = 16'h8484;
    SB_DFFE data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31950));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5291), .S(n59825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5292), .S(n59824));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31947));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5293), .S(n59823));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5294), .S(n31262));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5295), .S(n59770));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n31539));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5296), .S(n59822));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5297), .S(n59821));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5298), .S(n59820));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5299), .S(n31257));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5300), .S(n59819));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5301), .S(n59818));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13921_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n31866));
    defparam i13921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13924_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n31869));
    defparam i13924_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i45318_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64588));
    defparam i45318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45317_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64587));
    defparam i45317_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5302), .S(n59817));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13927_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n31872));
    defparam i13927_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[20] [2]), .I1(n54636), .I2(n55690), 
            .I3(\data_out_frame[22] [3]), .O(n62640));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_222_i3_4_lut (.I0(n5), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60437), .I3(n61755), .O(n3_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFE data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5304), .S(n59816));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5305), .S(n59946));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[20] [2]), .I1(n54636), 
            .I2(n55641), .I3(\data_out_frame[20] [3]), .O(n55627));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5306), .S(n59945));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut (.I0(control_mode[0]), .I1(n27629), .I2(GND_net), 
            .I3(GND_net), .O(n51206));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[20] [3]), .I1(n55641), .I2(n60634), 
            .I3(GND_net), .O(n60635));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5307), .S(n59944));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5308), .S(n59815));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i34347_4_lut (.I0(displacement[10]), .I1(\encoder0_position_scaled[10] ), 
            .I2(n54181), .I3(n51206), .O(n8));
    defparam i34347_4_lut.LUT_INIT = 16'hf353;
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5310), .S(n59943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5311), .S(n59942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5312), .S(n59941));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1084 (.I0(\data_out_frame[17] [7]), .I1(n28889), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n60775));
    defparam i1_2_lut_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1085 (.I0(\data_out_frame[17] [7]), .I1(n28889), 
            .I2(n60381), .I3(GND_net), .O(n6_c));
    defparam i1_2_lut_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5314), .S(n31251));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_221_i3_4_lut (.I0(n62178), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60437), .I3(\data_out_frame[25] [3]), .O(n3_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_789_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_220_i3_4_lut (.I0(n62178), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60434), .I3(n55008), .O(n3_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1086 (.I0(n60322), .I1(n60695), .I2(\data_out_frame[18] [4]), 
            .I3(GND_net), .O(n54659));
    defparam i1_2_lut_3_lut_adj_1086.LUT_INIT = 16'h9696;
    SB_LUT4 i23560_2_lut (.I0(LED_c), .I1(LED_N_3408), .I2(GND_net), .I3(GND_net), 
            .O(LED_N_3407));   // verilog/coms.v(253[15] 255[9])
    defparam i23560_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1087 (.I0(n60322), .I1(n60695), .I2(n27913), 
            .I3(n55659), .O(n55663));
    defparam i2_3_lut_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13105_4_lut (.I0(n2889), .I1(LED_N_3407), .I2(n29481), .I3(\FRAME_MATCHER.i_31__N_2513 ), 
            .O(n31050));   // verilog/coms.v(130[12] 305[6])
    defparam i13105_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 select_1745_Select_0_i3_3_lut (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n3_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i3_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut (.I0(LED_c), .I1(n3_adj_5319), .I2(Kp_23__N_1748), 
            .I3(Kp_23__N_612), .O(n5_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5321), .S(n59947));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5322), .S(n59814));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5323), .S(n59813));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5324), .S(n59812));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5325), .S(n59811));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5326), .S(n59810));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5327), .S(n59809));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5328), .S(n59808));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5329), .S(n59807));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n60227), .I1(n60592), .I2(n54689), .I3(\data_out_frame[25] [4]), 
            .O(n60437));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5330), .S(n59806));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5331), .S(n59805));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut (.I0(n55665), .I1(n55663), .I2(n60359), .I3(GND_net), 
            .O(n8_adj_5333));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5334), .S(n59804));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5335), .S(n59940));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1088 (.I0(n60227), .I1(n60592), .I2(n54689), 
            .I3(n60359), .O(n8_adj_5336));
    defparam i1_2_lut_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_219_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5333), .I3(\data_out_frame[25] [2]), 
            .O(n3_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_219_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5338), .S(n59939));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5340), .S(n59803));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5341), .S(n31237));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1089 (.I0(n10), .I1(n152), .I2(GND_net), .I3(GND_net), 
            .O(n30382));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'heeee;
    SB_LUT4 select_789_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n60440), .I3(n55546), .O(n3_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[23] [2]), .I1(n28303), .I2(n60689), 
            .I3(n55645), .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut (.I0(n27913), .I1(n18), .I2(n60449), .I3(n60695), 
            .O(n20));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n60692), .I1(n20), .I2(n16), .I3(n60672), 
            .O(n62178));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[18] [5]), .I1(n55719), .I2(n62514), 
            .I3(GND_net), .O(n16_adj_5345));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5346), .S(n59802));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5347), .S(n59938));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut (.I0(n28864), .I1(n60452), .I2(n60756), .I3(n60672), 
            .O(n16_adj_5349));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[19] [2]), .I1(n28963), .I2(GND_net), 
            .I3(GND_net), .O(n15));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1090 (.I0(n60362), .I1(n60797), .I2(\data_out_frame[16] [7]), 
            .I3(n28869), .O(n17));
    defparam i7_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(\data_out_frame[23] [0]), .I1(n17), .I2(n15), 
            .I3(n16_adj_5349), .O(n55546));
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i7_4_lut_adj_1092 (.I0(n55546), .I1(n60692), .I2(n54936), 
            .I3(n60227), .O(n18_adj_5350));
    defparam i7_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1093 (.I0(\data_out_frame[16] [3]), .I1(n18_adj_5350), 
            .I2(\data_out_frame[22] [7]), .I3(n60076), .O(n20_adj_5352));
    defparam i9_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1094 (.I0(n55770), .I1(n20_adj_5352), .I2(n16_adj_5345), 
            .I3(\data_out_frame[16] [4]), .O(n55008));
    defparam i10_4_lut_adj_1094.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5353), .S(n59937));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_out_frame[21] [0]), .I1(n27161), 
            .I2(GND_net), .I3(GND_net), .O(n60227));
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[22] [6]), .I1(n55008), .I2(\data_out_frame[24] [7]), 
            .I3(n6_adj_5354), .O(n60359));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5357), .S(n59936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5358), .S(n59935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5359), .S(n59934));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5360), .S(n59933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5361), .S(n59932));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5362), .S(n59931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5363), .S(n59930));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut (.I0(n55665), .I1(n55663), .I2(n55737), .I3(n62178), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5364), .S(n59929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5365), .S(n59928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5366), .S(n59927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5367), .S(n59926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5368), .S(n59925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5369), .S(n59924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5370), .S(n59801));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5371), .S(n59800));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5372), .S(n59799));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5373), .S(n59798));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5374), .S(n59797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5375), .S(n59796));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5376), .S(n59923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5377), .S(n59795));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5378), .S(n59922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5379), .S(n59794));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5380), .S(n59793));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1096 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(n60142), .I3(n60331), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5381), .S(n59921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5382), .S(n59792));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5383), .S(n59791));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5384), .S(n59920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5385), .S(n59790));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5386), .S(n59789));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5387), .S(n59788));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5388), .S(n59787));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5389), .S(n59786));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5390), .S(n59785));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5391), .S(n59784));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5393), .S(n59919));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5394), .S(n59783));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_217_i3_4_lut (.I0(n55784), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12), .I3(n8_adj_5336), .O(n3_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_217_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_3_lut_adj_1097 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n60331));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1097.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1098 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n60545));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[25] [0]), .I1(n55665), .I2(\data_out_frame[24] [6]), 
            .I3(n60073), .O(n60440));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5398), .S(n59782));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5399), .S(n59781));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5400), .S(n59780));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_216_i3_4_lut (.I0(n61872), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60440), .I3(n55737), .O(n3_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_216_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5402), .S(n59779));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5404), .S(n59778));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5405), .S(n59777));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60434));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1100 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60592));
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5406), .S(n59918));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_out_frame[22] [5]), .I1(n55776), 
            .I2(GND_net), .I3(GND_net), .O(n60794));
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1102 (.I0(n60478), .I1(n55561), .I2(\data_out_frame[19] [0]), 
            .I3(\data_out_frame[21] [1]), .O(n14));
    defparam i6_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1103 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1103.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1104 (.I0(n9), .I1(n14), .I2(n62514), .I3(n55719), 
            .O(n28608));
    defparam i7_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1105 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [7]), 
            .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n13));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1105.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31897));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60431));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1107 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [6]), 
            .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1107.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5409), .S(n59776));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1108 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(n27161), .I3(\data_out_frame[20] [6]), .O(n60756));
    defparam i3_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n60643), .I1(n55663), .I2(\data_out_frame[23] [0]), 
            .I3(n54606), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_2_lut_3_lut_adj_1109 (.I0(\data_out_frame[18] [5]), .I1(n55719), 
            .I2(\data_out_frame[21] [1]), .I3(GND_net), .O(n16));
    defparam i5_2_lut_3_lut_adj_1109.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5412), .S(n59775));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut_adj_1110 (.I0(n60424), .I1(\data_out_frame[22] [7]), 
            .I2(n55550), .I3(n60756), .O(n24));
    defparam i10_4_lut_adj_1110.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1111 (.I0(\data_out_frame[21] [0]), .I1(n55706), 
            .I2(n28608), .I3(n60794), .O(n23));
    defparam i9_4_lut_adj_1111.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut (.I0(n60634), .I1(n22), .I2(n54695), .I3(GND_net), 
            .O(n25));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1112 (.I0(n28608), .I1(\data_out_frame[23] [3]), 
            .I2(\data_out_frame[25] [5]), .I3(GND_net), .O(n5));
    defparam i1_2_lut_3_lut_adj_1112.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5414), .S(n59774));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5415), .S(n59773));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5417), .S(n59772));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5418), .S(n59771));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5420), .S(n59832));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5][4] ), .C(clk16MHz), 
           .D(n31542));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_215_i3_4_lut (.I0(n55737), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5423), .I3(\data_out_frame[24] [5]), .O(n3_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_789_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5425), .S(n59968));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in_frame[2] [6]), .I1(n60272), .I2(\data_in_frame[2][1] ), 
            .I3(Kp_23__N_748), .O(n16_adj_5426));   // verilog/coms.v(99[12:25])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0990;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[1] [4]), .I1(n60337), .I2(n55542), 
            .I3(n60416), .O(n62335));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1113 (.I0(\data_in_frame[1] [4]), .I1(n60337), 
            .I2(n60548), .I3(n60115), .O(n28027));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60470));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1115 (.I0(\FRAME_MATCHER.state[3] ), .I1(n62640), 
            .I2(n60470), .I3(n60635), .O(n3_adj_5427));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1115.LUT_INIT = 16'h2882;
    SB_LUT4 select_789_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5428));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5429));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_213_i3_4_lut (.I0(n62640), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60487), .I3(\data_out_frame[24] [4]), .O(n3_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5431), .S(n59917));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26][1] ), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5433), .S(n59967));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(n10_adj_5434), .I3(\data_in_frame[3] [6]), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26][2] ), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5435), .S(n59966));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2081), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52077 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n71380));
    defparam byte_transmit_counter_0__bdd_4_lut_52077.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_4_lut (.I0(n28432), .I1(n60296), .I2(n36324), .I3(\data_in_frame[8] [7]), 
            .O(n7));   // verilog/coms.v(18[27:29])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1116 (.I0(n28608), .I1(\data_out_frame[23] [3]), 
            .I2(n61872), .I3(GND_net), .O(n55784));
    defparam i1_2_lut_3_lut_adj_1116.LUT_INIT = 16'h6969;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n29831), 
            .D(n4947[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1117 (.I0(n28432), .I1(n60296), .I2(n36324), 
            .I3(n55186), .O(n55565));   // verilog/coms.v(18[27:29])
    defparam i1_2_lut_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5437), .S(n59965));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1118 (.I0(\data_in_frame[6] [7]), .I1(n27900), 
            .I2(n28432), .I3(GND_net), .O(n60584));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1118.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1119 (.I0(\data_in_frame[6] [7]), .I1(n27900), 
            .I2(n60723), .I3(n60562), .O(n28386));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5438), .S(n59964));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31890));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5430), .S(n59962));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1120 (.I0(\data_in_frame[21] [7]), .I1(n55653), 
            .I2(n60150), .I3(GND_net), .O(n6_adj_5440));
    defparam i1_2_lut_3_lut_adj_1120.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5428), .S(n59916));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5427), .S(n59963));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5424), .S(n59970));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5401), .S(n59956));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71380_bdd_4_lut (.I0(n71380), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n71383));
    defparam n71380_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27][1] ), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5396), .S(n59961));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_3_lut_4_lut_adj_1121 (.I0(\data_in_frame[21] [7]), .I1(n55653), 
            .I2(n62393), .I3(\data_in_frame[21]_c [6]), .O(n8_adj_5442));
    defparam i3_3_lut_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27][2] ), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5344), .S(n59957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5337), .S(n59958));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2889), .D(n5_adj_5320), 
            .S(n31050));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1122 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [1]), 
            .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1122.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_95_i2_4_lut (.I0(\data_out_frame[11][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5317), .S(n59955));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5315), .S(n59959));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_94_i2_4_lut (.I0(\data_out_frame[11][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_93_i2_4_lut (.I0(\data_out_frame[11][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_92_i2_4_lut (.I0(\data_out_frame[11][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_91_i2_4_lut (.I0(\data_out_frame[11][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2889), .D(n3_adj_5303), .S(n59960));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52087 (.I0(byte_transmit_counter[1]), 
            .I1(n64587), .I2(n64588), .I3(byte_transmit_counter[2]), .O(n71374));
    defparam byte_transmit_counter_1__bdd_4_lut_52087.LUT_INIT = 16'he4aa;
    SB_LUT4 select_789_Select_90_i2_4_lut (.I0(\data_out_frame[11][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_89_i2_4_lut (.I0(\data_out_frame[11][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(n28529), .I1(n4_c), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n28134));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2889), .D(n3), .S(n59969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2889), .D(n1_c), .S(n59759));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5452), .S(n59915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2889), .D(n1_adj_5453), .S(n59760));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(clk16MHz), .E(n2889), .D(n1_adj_5454), .S(n59762));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1124 (.I0(n28529), .I1(n4_c), .I2(n60607), 
            .I3(n60309), .O(n64019));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31886));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71374_bdd_4_lut (.I0(n71374), .I1(n64915), .I2(n64914), .I3(byte_transmit_counter[2]), 
            .O(n71377));
    defparam n71374_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5457), .S(n59914));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_789_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_789_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52072 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n71368));
    defparam byte_transmit_counter_0__bdd_4_lut_52072.LUT_INIT = 16'he4aa;
    SB_LUT4 select_789_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(clk16MHz), .E(n2889), .D(n1_adj_5460), .S(n59763));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2889), .D(n1_adj_5462), .S(n59764));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1125 (.I0(n28055), .I1(n28074), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[14] [7]), .O(n64173));   // verilog/coms.v(78[16:43])
    defparam i1_3_lut_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 n71368_bdd_4_lut (.I0(n71368), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71371));
    defparam n71368_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2889), .D(n1_adj_5463), .S(n59761));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14][2] ), .C(clk16MHz), 
            .E(VCC_net), .D(n31881));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n31878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5465), .S(n59913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n31875));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31872));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5467));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'hbbbb;
    SB_DFFE data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31869));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5469), .S(n59912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31866));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5470), .S(n59911));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5][5] ), .C(clk16MHz), 
           .D(n31545));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2889), .D(n1_adj_5471), .S(n59765));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31862));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31859));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1127 (.I0(n28055), .I1(n28074), .I2(Kp_23__N_1389), 
            .I3(\data_in_frame[13] [5]), .O(n4_adj_5474));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5478));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1128 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[14] [6]), .I3(n60659), .O(n64167));
    defparam i1_3_lut_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_out_frame[24] [3]), .I1(n55739), 
            .I2(GND_net), .I3(GND_net), .O(n60487));
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52067 (.I0(byte_transmit_counter[1]), 
            .I1(n64584), .I2(n64585), .I3(byte_transmit_counter[2]), .O(n71362));
    defparam byte_transmit_counter_1__bdd_4_lut_52067.LUT_INIT = 16'he4aa;
    SB_LUT4 select_789_Select_211_i3_4_lut (.I0(n25812), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60254), .I3(\data_out_frame[24] [1]), .O(n3_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1130 (.I0(n60763), .I1(n28877), .I2(\data_in_frame[20] [6]), 
            .I3(\data_in_frame[21][0] ), .O(n64037));
    defparam i1_4_lut_adj_1130.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1131 (.I0(n27332), .I1(n60601), .I2(n60248), 
            .I3(n64037), .O(n55671));
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5479));
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(n55778), .I1(n54264), .I2(\data_in_frame[20] [5]), 
            .I3(n6_adj_5479), .O(n60306));
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1134 (.I0(\data_in_frame[21][1] ), .I1(\data_in_frame[21][4] ), 
            .I2(n60260), .I3(n6_adj_5440), .O(n55708));
    defparam i4_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n64213));
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5306));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1136 (.I0(n60604), .I1(\data_in_frame[19] [0]), 
            .I2(n64213), .I3(\data_in_frame[20] [7]), .O(n64219));
    defparam i1_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1137 (.I0(n60540), .I1(n60495), .I2(n64219), 
            .I3(n60656), .O(n64225));
    defparam i1_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1138 (.I0(n60800), .I1(\data_in_frame[18]_c [7]), 
            .I2(n64225), .I3(n60579), .O(n64229));
    defparam i1_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1139 (.I0(n54773), .I1(n60765), .I2(n64229), 
            .I3(n60275), .O(n64235));
    defparam i1_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1140 (.I0(n55766), .I1(n60458), .I2(n60306), 
            .I3(n64235), .O(n64241));
    defparam i1_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1141 (.I0(n61855), .I1(n62783), .I2(n64241), 
            .I3(n60388), .O(n62602));
    defparam i1_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(n62602), .I1(n55708), .I2(GND_net), 
            .I3(GND_net), .O(n60443));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h9999;
    SB_LUT4 select_789_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5304));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut (.I0(n54740), .I1(\data_in_frame[19]_c [5]), .I2(n28247), 
            .I3(n55653), .O(n55766));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[21][5] ), .I1(n55766), .I2(\data_in_frame[21]_c [6]), 
            .I3(GND_net), .O(n60260));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(n55653), .I1(n61855), .I2(GND_net), 
            .I3(GND_net), .O(n26003));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[19]_c [6]), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n60495));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[18][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28753));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1146 (.I0(n28753), .I1(n28002), .I2(n28507), 
            .I3(\data_in_frame[18] [5]), .O(n60278));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 n71362_bdd_4_lut (.I0(n71362), .I1(n64882), .I2(n64881), .I3(byte_transmit_counter[2]), 
            .O(n71365));
    defparam n71362_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(n54742), .I1(n54649), .I2(n60785), 
            .I3(\data_in_frame[14] [7]), .O(n64011));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1148 (.I0(n60759), .I1(n60701), .I2(n60765), 
            .I3(GND_net), .O(n8_adj_5480));
    defparam i3_3_lut_adj_1148.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n60190), .I1(\data_in_frame[16] [0]), 
            .I2(n6_adj_5481), .I3(n60368), .O(n64003));
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1150 (.I0(n60698), .I1(n60662), .I2(n55643), 
            .I3(n64011), .O(n62107));
    defparam i1_4_lut_adj_1150.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1151 (.I0(n54647), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [3]), .I3(\data_in_frame[15] [6]), .O(n64057));
    defparam i1_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1152 (.I0(\data_in_frame[16] [7]), .I1(n64003), 
            .I2(n8_adj_5480), .I3(Kp_23__N_1389), .O(n64005));
    defparam i1_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1153 (.I0(n64005), .I1(n64057), .I2(n64061), 
            .I3(n62107), .O(n60817));
    defparam i1_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1154 (.I0(n28908), .I1(n60461), .I2(\data_in_frame[18][0] ), 
            .I3(\data_in_frame[17][5] ), .O(n64081));
    defparam i1_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1155 (.I0(n55556), .I1(n64089), .I2(n64081), 
            .I3(n60817), .O(n10_adj_5482));
    defparam i2_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1156 (.I0(n54264), .I1(\data_in_frame[16] [5]), 
            .I2(n60473), .I3(n61729), .O(n14_adj_5483));
    defparam i6_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(n62783), .I1(n60278), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5484));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1158 (.I0(n61984), .I1(n9_adj_5484), .I2(n14_adj_5483), 
            .I3(n10_adj_5482), .O(n60682));
    defparam i1_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\data_in_frame[13] [7]), .I1(n60698), 
            .I2(GND_net), .I3(GND_net), .O(n27332));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[18][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n60512));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[17] [1]), .I1(n54563), 
            .I2(GND_net), .I3(GND_net), .O(n54647));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1162 (.I0(\data_in_frame[16] [7]), .I1(n60374), 
            .I2(n55712), .I3(\data_in_frame[12] [3]), .O(n62306));
    defparam i3_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(n62554), .I1(n60461), .I2(GND_net), 
            .I3(GND_net), .O(n27873));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(n62393), .I1(n28247), .I2(GND_net), 
            .I3(GND_net), .O(n28908));
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_in_frame[19][7] ), .I1(\data_in_frame[19]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60604));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5486));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31853));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n60368));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n60656));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1168 (.I0(n54662), .I1(n60622), .I2(n60396), 
            .I3(\data_in_frame[11] [5]), .O(n12_adj_5487));
    defparam i5_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1169 (.I0(n60319), .I1(n12_adj_5487), .I2(\data_in_frame[13] [7]), 
            .I3(n60656), .O(n27223));
    defparam i6_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1170 (.I0(n55565), .I1(n27843), .I2(\data_in_frame[14][1] ), 
            .I3(n60791), .O(n10_adj_5488));
    defparam i4_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n27865), .I1(n10_adj_5488), .I2(n55542), .I3(GND_net), 
            .O(n60508));
    defparam i5_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1171 (.I0(n60508), .I1(\data_in_frame[13] [5]), 
            .I2(n28055), .I3(n60622), .O(n10_adj_5489));
    defparam i4_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1172 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[20] [4]), 
            .I2(n27223), .I3(\data_in_frame[20] [3]), .O(n54773));
    defparam i3_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1173 (.I0(n60619), .I1(\data_in_frame[14][0] ), 
            .I2(n28074), .I3(GND_net), .O(n60785));
    defparam i2_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1174 (.I0(n27294), .I1(n60132), .I2(n28126), 
            .I3(\data_in_frame[15] [7]), .O(n54620));
    defparam i3_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(n54620), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[16] [0]), .I3(GND_net), .O(n60396));
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1176 (.I0(n27810), .I1(n60312), .I2(n28559), 
            .I3(GND_net), .O(n60619));
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1177 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [6]), 
            .I2(n60396), .I3(\data_in_frame[13] [3]), .O(n20_adj_5491));   // verilog/coms.v(88[17:63])
    defparam i8_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1178 (.I0(\data_in_frame[14][0] ), .I1(n60619), 
            .I2(n60094), .I3(\data_in_frame[13] [5]), .O(n19));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1179 (.I0(\data_in_frame[13] [7]), .I1(n60105), 
            .I2(n54620), .I3(n28055), .O(n21));   // verilog/coms.v(88[17:63])
    defparam i9_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31850));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_3_lut_adj_1180 (.I0(n21), .I1(n19), .I2(n20_adj_5491), 
            .I3(GND_net), .O(n62103));   // verilog/coms.v(88[17:63])
    defparam i11_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1181 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[14][2] ), 
            .I2(Kp_23__N_1271), .I3(n6_adj_5492), .O(n60248));
    defparam i4_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1182 (.I0(n60248), .I1(\data_in_frame[16] [3]), 
            .I2(n62103), .I3(GND_net), .O(n55556));
    defparam i2_3_lut_adj_1182.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(\data_in_frame[18][2] ), .I1(\data_in_frame[18][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n28507));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(n55186), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60484));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[6][3] ), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[8] [3]), .O(n26));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1185 (.I0(n54872), .I1(n60607), .I2(n55163), 
            .I3(n60428), .O(n16_adj_5494));
    defparam i1_4_lut_adj_1185.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31847));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1186 (.I0(\data_in_frame[1] [6]), .I1(n28572), 
            .I2(\data_in_frame[8] [6]), .I3(n60176), .O(n24_adj_5495));
    defparam i9_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[4] [2]), .I1(n26), .I2(n20_adj_5496), 
            .I3(\data_in_frame[8] [4]), .O(n28_c));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[9] [6]), .I1(n28_c), .I2(n24_adj_5495), 
            .I3(n16_adj_5494), .O(n60791));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[6][5] ), .I1(Kp_23__N_1080), .I2(\data_in_frame[5][0] ), 
            .I3(Kp_23__N_875), .O(n28_adj_5497));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1187 (.I0(n60726), .I1(\data_in_frame[11] [6]), 
            .I2(n60287), .I3(n54597), .O(n26_adj_5498));
    defparam i10_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31844));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_4_lut_adj_1188 (.I0(n60791), .I1(n60467), .I2(n60562), 
            .I3(n60217), .O(n27_c));
    defparam i11_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1189 (.I0(n54746), .I1(n60484), .I2(n60208), 
            .I3(\data_in_frame[9] [0]), .O(n25_adj_5499));
    defparam i9_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n25_adj_5499), .I1(n27_c), .I2(n26_adj_5498), 
            .I3(n28_adj_5497), .O(n27251));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31841));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_71_i2_4_lut (.I0(\data_out_frame[8][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5][6] ), .C(clk16MHz), 
           .D(n31548));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5][7] ), .C(clk16MHz), 
           .D(n31551));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5486), .S(n59910));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_70_i2_4_lut (.I0(\data_out_frame[8][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31833));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_791_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5476), .S(n59909));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[18]_c [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28002));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31827));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31824));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31821));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_in_frame[14] [7]), .I1(n60659), 
            .I2(\data_in_frame[12] [5]), .I3(\data_in_frame[14] [5]), .O(n60374));
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_69_i2_4_lut (.I0(\data_out_frame[8][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_in_frame[19][2] ), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5504));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(n60374), .I1(n60235), .I2(n60759), 
            .I3(n6_adj_5504), .O(n60388));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31818));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1194 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[21]_c [2]), 
            .I2(\data_in_frame[21][3] ), .I3(n27264), .O(n60150));
    defparam i3_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1195 (.I0(n55712), .I1(n60726), .I2(\data_in_frame[12] [2]), 
            .I3(n55186), .O(n12_adj_5505));
    defparam i5_4_lut_adj_1195.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1196 (.I0(n55163), .I1(n12_adj_5505), .I2(\data_in_frame[14]_c [3]), 
            .I3(\data_in_frame[9] [6]), .O(n60190));
    defparam i6_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1197 (.I0(n54624), .I1(n60518), .I2(\data_in_frame[14] [4]), 
            .I3(GND_net), .O(n61729));
    defparam i2_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31815));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1198 (.I0(n61729), .I1(n60190), .I2(GND_net), 
            .I3(GND_net), .O(n55643));
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[12] [3]), .I1(n55712), 
            .I2(GND_net), .I3(GND_net), .O(n60235));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1200 (.I0(\data_in_frame[14] [6]), .I1(n28126), 
            .I2(\data_in_frame[12] [4]), .I3(n54626), .O(n54742));
    defparam i3_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(n54742), .I1(\data_in_frame[17][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n60649));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1202 (.I0(\data_in_frame[14] [5]), .I1(n28583), 
            .I2(n60235), .I3(\data_in_frame[12] [4]), .O(n54649));
    defparam i3_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31812));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31809));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_68_i2_4_lut (.I0(\data_out_frame[8][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1203 (.I0(\data_in_frame[19]_c [1]), .I1(n54649), 
            .I2(n60649), .I3(n6_adj_5507), .O(n60579));
    defparam i4_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1204 (.I0(n60224), .I1(\data_in_frame[15] [6]), 
            .I2(n28055), .I3(GND_net), .O(n60094));
    defparam i2_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1205 (.I0(\data_in_frame[13] [4]), .I1(n60094), 
            .I2(\data_in_frame[18][0] ), .I3(GND_net), .O(n60540));
    defparam i2_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17][7] ), 
            .I1(\data_in_frame[17][6] ), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1206 (.I0(\data_in_frame[20] [2]), .I1(n60540), 
            .I2(n62554), .I3(n4_adj_5474), .O(n60481));
    defparam i2_4_lut_adj_1206.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_67_i2_4_lut (.I0(\data_out_frame[8][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5508));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31806));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31803));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31800));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31794));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31791));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31788));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31785));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_66_i2_4_lut (.I0(\data_out_frame[8][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n64187));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31782));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_65_i2_4_lut (.I0(\data_out_frame[8][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31779));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1208 (.I0(n55482), .I1(n60646), .I2(n26045), 
            .I3(n64187), .O(n54624));
    defparam i1_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31776));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1209 (.I0(n28583), .I1(n54624), .I2(GND_net), 
            .I3(GND_net), .O(n54626));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31773));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31770));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n29831), 
            .D(n4947[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_in_frame[11] [6]), .I1(n26041), 
            .I2(GND_net), .I3(GND_net), .O(n60312));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(n55163), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60467));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n29831), 
            .D(n4947[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n29831), 
            .D(n4947[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31767));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(n28572), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n54746));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n29831), 
            .D(n4947[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60806));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60428));
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(n60167), .I1(n60428), .I2(\data_in_frame[9] [7]), 
            .I3(\data_in_frame[10] [1]), .O(n64067));
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i51639_4_lut (.I0(Kp_23__N_1067), .I1(n55710), .I2(n60051), 
            .I3(n55186), .O(n70909));
    defparam i51639_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64195));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n29831), 
            .D(n4947[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n29831), 
            .D(n4947[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n29831), 
            .D(n4947[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n29831), 
            .D(n4947[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n29831), 
            .D(n4947[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n29831), 
            .D(n4947[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n29831), 
            .D(n4947[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n29831), 
            .D(n4947[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n29831), 
            .D(n4947[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n29831), 
            .D(n4947[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n29831), 
            .D(n4947[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n29831), 
            .D(n4947[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n29831), 
            .D(n4947[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n29831), 
            .D(n4947[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n29831), 
            .D(n4947[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n29831), 
            .D(n4947[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n29831), 
            .D(n4947[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n29831), 
            .D(n4947[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6][0] ), .C(clk16MHz), 
           .D(n59122));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6][1] ), .C(clk16MHz), 
           .D(n31557));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6][2] ), .C(clk16MHz), 
           .D(n59126));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6][3] ), .C(clk16MHz), 
           .D(n59114));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6][4] ), .C(clk16MHz), 
           .D(n31566));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[11] [2]), .I3(GND_net), .O(n64197));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6][5] ), .C(clk16MHz), 
           .D(n59110));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1217 (.I0(n60559), .I1(n64197), .I2(n60806), 
            .I3(n64195), .O(n64203));
    defparam i1_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n29831), 
            .D(n4947[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6][6] ), .C(clk16MHz), 
           .D(n58986));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1218 (.I0(n54872), .I1(n70909), .I2(n60312), 
            .I3(n64067), .O(n64073));
    defparam i1_4_lut_adj_1218.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52057 (.I0(byte_transmit_counter[1]), 
            .I1(n64647), .I2(n64648), .I3(byte_transmit_counter[2]), .O(n71350));
    defparam byte_transmit_counter_1__bdd_4_lut_52057.LUT_INIT = 16'he4aa;
    SB_LUT4 n71350_bdd_4_lut (.I0(n71350), .I1(n64717), .I2(n64716), .I3(byte_transmit_counter[2]), 
            .O(n71353));
    defparam n71350_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1219 (.I0(n60518), .I1(n28386), .I2(n60720), 
            .I3(n64203), .O(n64209));
    defparam i1_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
           .D(n31576));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1220 (.I0(n64209), .I1(n60102), .I2(n64073), 
            .I3(n60769), .O(n27294));
    defparam i1_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n31583));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1271));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n31586));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n31625));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5513), .S(n59908));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1221 (.I0(n60559), .I1(n60584), .I2(\data_in_frame[8] [7]), 
            .I3(n60135), .O(n12_adj_5514));   // verilog/coms.v(18[27:29])
    defparam i5_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1222 (.I0(n36324), .I1(n12_adj_5514), .I2(n60723), 
            .I3(n24_adj_5515), .O(n28055));   // verilog/coms.v(18[27:29])
    defparam i6_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i15_2_lut (.I0(n54662), .I1(n28055), .I2(GND_net), .I3(GND_net), 
            .O(n58710));
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1223 (.I0(n60548), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[10] [3]), .I3(n60613), .O(n10_adj_5516));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1224 (.I0(n60105), .I1(n54602), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[13] [2]), .O(n28834));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31745));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1225 (.I0(\data_in_frame[9] [3]), .I1(n27843), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n28074));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31742));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31739));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n71700), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n29158), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2061), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2062), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n23276), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n58832), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2073), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n29161), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31736));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1226 (.I0(n28074), .I1(n60319), .I2(GND_net), 
            .I3(GND_net), .O(n54857));
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31733));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5517), .S(n59907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31730));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31727));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(\data_in_frame[17][3] ), .I1(n62185), 
            .I2(GND_net), .I3(GND_net), .O(n60800));
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h9999;
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31724));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1228 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [4]), 
            .I2(n60220), .I3(n28041), .O(n60720));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31721));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1229 (.I0(\data_in_frame[13] [0]), .I1(n28126), 
            .I2(\data_in_frame[15] [4]), .I3(Kp_23__N_1067), .O(n64061));
    defparam i1_3_lut_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31718));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31715));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(\data_in_frame[13] [0]), .I1(n28126), 
            .I2(n28834), .I3(GND_net), .O(n60319));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31712));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1196_9_lut (.I0(n59757), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n52659), .O(n59765)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_in_frame[15] [0]), .I1(n60720), 
            .I2(GND_net), .I3(GND_net), .O(n60659));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 add_1196_8_lut (.I0(n59757), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n52658), .O(n59761)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1232 (.I0(n55574), .I1(n60800), .I2(n60772), 
            .I3(n60662), .O(n28247));
    defparam i3_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31709));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_789_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n31688));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1233 (.I0(n58710), .I1(n28834), .I2(n60738), 
            .I3(n64173), .O(n64179));
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1234 (.I0(n60769), .I1(n64179), .I2(n64167), 
            .I3(n54857), .O(n54563));
    defparam i1_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31705));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n31691));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60701));
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60132));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n31694));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1237 (.I0(n60132), .I1(n60524), .I2(\data_in_frame[10] [7]), 
            .I3(n27956), .O(n12_adj_5521));
    defparam i5_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n31697));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1238 (.I0(n28134), .I1(n12_adj_5521), .I2(n60701), 
            .I3(\data_in_frame[12] [7]), .O(n62185));
    defparam i6_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1239 (.I0(\data_in_frame[12] [5]), .I1(n28583), 
            .I2(n28134), .I3(GND_net), .O(n28126));
    defparam i1_2_lut_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27810));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28366));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_CARRY add_1196_8 (.CI(n52658), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n52659));
    SB_LUT4 add_1196_7_lut (.I0(n59757), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n52657), .O(n59764)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n60105));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1085));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(n28529), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60220));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60587));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_CARRY add_1196_7 (.CI(n52657), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n52658));
    SB_LUT4 add_1196_6_lut (.I0(n59757), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n52656), .O(n59763)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1245 (.I0(n54662), .I1(n60587), .I2(n60220), 
            .I3(n27956), .O(n60738));
    defparam i3_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1246 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n27865));
    defparam i2_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1247 (.I0(\data_in_frame[8] [6]), .I1(n27865), 
            .I2(n28398), .I3(\data_in_frame[11] [2]), .O(n60224));
    defparam i3_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(n27956), .I1(n28041), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1249 (.I0(\data_in_frame[8] [5]), .I1(n60284), 
            .I2(\data_in_frame[6][3] ), .I3(Kp_23__N_872), .O(n27956));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(n27956), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60167));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60607));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1252 (.I0(\data_in_frame[7] [7]), .I1(n60293), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n27971));
    defparam i2_3_lut_adj_1252.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(n27971), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60631));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_CARRY add_1196_6 (.CI(n52656), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n52657));
    SB_LUT4 i3_4_lut_adj_1254 (.I0(n28490), .I1(n60631), .I2(n60337), 
            .I3(\data_in_frame[5][7] ), .O(n27992));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52048 (.I0(byte_transmit_counter[1]), 
            .I1(n64638), .I2(n64639), .I3(byte_transmit_counter[2]), .O(n71332));
    defparam byte_transmit_counter_1__bdd_4_lut_52048.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(n27992), .I1(n62335), .I2(GND_net), 
            .I3(GND_net), .O(n60646));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(n26041), .I1(n26045), .I2(GND_net), 
            .I3(GND_net), .O(n60251));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 n71332_bdd_4_lut (.I0(n71332), .I1(n64624), .I2(n64623), .I3(byte_transmit_counter[2]), 
            .O(n71335));
    defparam n71332_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_1196_5_lut (.I0(n59757), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n52655), .O(n59762)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_5_lut.LUT_INIT = 16'h8228;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2889), .D(n29032), 
            .S(n31014));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1196_5 (.CI(n52655), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n52656));
    SB_LUT4 i1_4_lut_adj_1257 (.I0(n64019), .I1(n7_adj_5523), .I2(Kp_23__N_1067), 
            .I3(n28386), .O(n64025));
    defparam i1_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1258 (.I0(n60251), .I1(n60646), .I2(n55565), 
            .I3(n64025), .O(n27211));
    defparam i1_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 add_1196_4_lut (.I0(n59757), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n52654), .O(n59760)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1196_4 (.CI(n52654), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n52655));
    SB_LUT4 i3_4_lut_adj_1259 (.I0(\data_in_frame[2][0] ), .I1(n60331), 
            .I2(\data_in_frame[4] [3]), .I3(n28463), .O(Kp_23__N_875));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\data_in_frame[6][4] ), .I1(Kp_23__N_875), 
            .I2(GND_net), .I3(GND_net), .O(n60284));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 add_1196_3_lut (.I0(n59757), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n52653), .O(n59759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1196_3 (.CI(n52653), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n52654));
    SB_LUT4 add_1196_2_lut (.I0(n59757), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n59758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1196_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1261 (.I0(Kp_23__N_1085), .I1(n28366), .I2(n27810), 
            .I3(\data_in_frame[9] [3]), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1262 (.I0(\data_in_frame[11] [1]), .I1(n27211), 
            .I2(n54872), .I3(GND_net), .O(n60102));
    defparam i1_3_lut_adj_1262.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1263 (.I0(n7), .I1(n60102), .I2(Kp_23__N_1080), 
            .I3(\data_in_frame[10] [7]), .O(n54662));
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 equal_2037_i7_2_lut (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5523));   // verilog/coms.v(239[9:81])
    defparam equal_2037_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_1196_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n52653));
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60051));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1265 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[13] [2]), .I3(GND_net), .O(n8_adj_5524));
    defparam i3_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1266 (.I0(n54662), .I1(n8_adj_5524), .I2(n61746), 
            .I3(n60224), .O(n62554));
    defparam i4_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1267 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n60738), .I3(\data_in_frame[13] [1]), .O(n55599));
    defparam i3_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(\data_in_frame[15] [3]), .I1(n62185), 
            .I2(\data_in_frame[17][4] ), .I3(GND_net), .O(n54740));
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5522), .S(n59906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5520), .S(n59905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5519), .S(n59904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5518), .S(n59833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5512), .S(n59903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5511), .S(n59902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8][1] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5510), .S(n59901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8][2] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5509), .S(n59900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8][3] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5508), .S(n59899));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8][4] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5506), .S(n59898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8][5] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5503), .S(n59897));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8][6] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5501), .S(n59896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8][7] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5500), .S(n59895));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5493), .S(n59894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5490), .S(n59893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5485), .S(n59892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5478), .S(n59891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5477), .S(n59890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5475), .S(n59889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5473), .S(n59888));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5472), .S(n59887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5468), .S(n59886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5466), .S(n59885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5464), .S(n59884));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5461), .S(n59883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5459), .S(n59882));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5458), .S(n59881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5456), .S(n59880));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5455), .S(n59879));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11][1] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5451), .S(n59878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11][2] ), .C(clk16MHz), 
            .E(n32669), .D(n2_adj_5450), .S(n31321));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11][3] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5449), .S(n59877));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11][4] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5448), .S(n59876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11][5] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5447), .S(n59875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11][6] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5446), .S(n59874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11][7] ), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5445), .S(n59873));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5444), .S(n59872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5443), .S(n59871));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5441), .S(n59870));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5439), .S(n59869));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5436), .S(n59868));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5432), .S(n59867));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5429), .S(n59866));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5422), .S(n59865));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5421), .S(n59864));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5419), .S(n59863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5416), .S(n59862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5413), .S(n59861));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5411), .S(n59860));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5410), .S(n59859));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5408), .S(n59834));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2889), .D(n13), .S(n59858));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n32691), .D(n2_adj_5407), .S(n31299));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5403), .S(n59857));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5397), .S(n59856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5395), .S(n59855));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5392), .S(n59854));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n31624));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5356), .S(n31294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n31623));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5355), .S(n59853));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n31622));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5351), .S(n59852));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n31621));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5348), .S(n59851));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n31620));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5343), .S(n59850));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n31619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5342), .S(n59849));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n31618));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5339), .S(n59848));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n31617));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5332), .S(n59847));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n31616));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n31615));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5318), .S(n59846));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n31614));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n31613));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n31612));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5316), .S(n59845));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n31611));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n31610));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n31609));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n32706), .D(n2_adj_5313), .S(n31284));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n31608));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n31607));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n31606));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n31605));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n31604));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n31603));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5525), .S(n59844));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n31602));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n31601));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n31600));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n31599));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n31598));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n31597));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5526), .S(n59843));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n31596));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n31595));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n31594));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5527), .S(n59842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n31590));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5528), .S(n59841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5529), .S(n59840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5530), .S(n59839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5531), .S(n31277));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5532), .S(n59838));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5533), .S(n59837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5534), .S(n59836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5535), .S(n59835));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1269 (.I0(n54563), .I1(\data_in_frame[19]_c [4]), 
            .I2(n28247), .I3(GND_net), .O(n55653));
    defparam i2_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5536), .S(n59831));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52035 (.I0(byte_transmit_counter[1]), 
            .I1(n64896), .I2(n64897), .I3(byte_transmit_counter[2]), .O(n71326));
    defparam byte_transmit_counter_1__bdd_4_lut_52035.LUT_INIT = 16'he4aa;
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2889), .D(n1_adj_5537), .S(n31004));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1270 (.I0(n54740), .I1(n55599), .I2(n62554), 
            .I3(\data_in_frame[17][5] ), .O(n62393));
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60135));   // verilog/coms.v(18[27:29])
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1272 (.I0(n28435), .I1(\data_in_frame[6][6] ), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[7] [0]), .O(n60208));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1273 (.I0(\data_in_frame[1] [7]), .I1(n60576), 
            .I2(n60176), .I3(n28435), .O(n36324));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2044__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n30058), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_2_lut_adj_1274 (.I0(n28296), .I1(n60173), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5538));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1275 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5][4] ), 
            .I2(n60111), .I3(n6_adj_5538), .O(n55163));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_869), 
            .I2(\data_in_frame[6][2] ), .I3(n28027), .O(n28529));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5539), .S(n59830));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1277 (.I0(n60208), .I1(n60584), .I2(GND_net), 
            .I3(GND_net), .O(n28398));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[2][4] ), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60122));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1279 (.I0(\data_in_frame[2][0] ), .I1(n28018), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[1] [4]), .O(n10_adj_5434));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 n71326_bdd_4_lut (.I0(n71326), .I1(n64603), .I2(n64602), .I3(byte_transmit_counter[2]), 
            .O(n71329));
    defparam n71326_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1280 (.I0(n28006), .I1(Kp_23__N_872), .I2(Kp_23__N_869), 
            .I3(\data_in_frame[8] [4]), .O(n28041));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1281 (.I0(\data_in_frame[5][1] ), .I1(\data_in_frame[5][0] ), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n14_adj_5540));
    defparam i5_3_lut_adj_1281.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1282 (.I0(n60122), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[2][5] ), .I3(n60079), .O(n15_adj_5541));
    defparam i6_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1283 (.I0(n15_adj_5541), .I1(\data_in_frame[2] [6]), 
            .I2(n14_adj_5540), .I3(\data_in_frame[4] [6]), .O(n28559));
    defparam i8_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5542), .S(n59829));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1284 (.I0(n28694), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[5][2] ), .I3(n60365), .O(n10_adj_5543));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1285 (.I0(n28296), .I1(n10_adj_5543), .I2(\data_in_frame[7] [4]), 
            .I3(GND_net), .O(n60217));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut_adj_1285.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(n60190), .I1(n60473), .I2(n28877), 
            .I3(GND_net), .O(n60275));
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52030 (.I0(byte_transmit_counter[1]), 
            .I1(n11), .I2(n12_adj_5544), .I3(byte_transmit_counter[2]), 
            .O(n71320));
    defparam byte_transmit_counter_1__bdd_4_lut_52030.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1287 (.I0(n27849), .I1(\data_in_frame[7] [6]), 
            .I2(n28009), .I3(GND_net), .O(n26045));
    defparam i2_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 select_791_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_791_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i4_4_lut_adj_1288 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_5545));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1288.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1289 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5546));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1289.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1290 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_5547));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1290.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1291 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5548));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1291.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1292 (.I0(n9_adj_5548), .I1(n11_adj_5547), .I2(n10_adj_5546), 
            .I3(n12_adj_5545), .O(n62747));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1292.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[5][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n60613));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60272));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[3]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60337));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28018));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(n60190), .I1(n60473), .I2(n60202), 
            .I3(GND_net), .O(n54264));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 select_791_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1298 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n60115));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1298.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n28490));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[0]), .O(n71518));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1300 (.I0(n28490), .I1(n60416), .I2(n60115), 
            .I3(\data_in_frame[1] [4]), .O(n28930));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[6][6] ), .I1(\data_in_frame[6][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5515));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_in_frame[5][5] ), .I1(n28009), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5549));
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(n61729), .I1(\data_in_frame[16] [6]), 
            .I2(n54649), .I3(GND_net), .O(n28877));
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1304 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3][3] ), 
            .I2(n27996), .I3(n6_adj_5549), .O(n60293));
    defparam i4_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1305 (.I0(\data_in_frame[14][2] ), .I1(n27251), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n60473));
    defparam i1_2_lut_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1306 (.I0(\data_in_frame[14][2] ), .I1(n27251), 
            .I2(\data_in_frame[11] [5]), .I3(n60508), .O(n60698));
    defparam i2_3_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2889), .D(n1_adj_5502), .S(n59758));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1307 (.I0(Kp_23__N_799), .I1(n54597), .I2(n60287), 
            .I3(n64047), .O(n55542));   // verilog/coms.v(88[17:28])
    defparam i1_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1308 (.I0(n55542), .I1(\data_in_frame[7] [7]), 
            .I2(n60293), .I3(GND_net), .O(n55482));
    defparam i2_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1309 (.I0(n27900), .I1(Kp_23__N_767), .I2(\data_in_frame[3]_c [1]), 
            .I3(n28296), .O(n14_adj_5550));   // verilog/coms.v(74[16:69])
    defparam i6_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1310 (.I0(\data_in_frame[0] [7]), .I1(n14_adj_5550), 
            .I2(n10_adj_5551), .I3(\data_in_frame[7] [3]), .O(n55186));   // verilog/coms.v(74[16:69])
    defparam i7_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1311 (.I0(n28027), .I1(n28930), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_c));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1312 (.I0(\data_in_frame[5][1] ), .I1(\data_in_frame[5][2] ), 
            .I2(\data_in_frame[4] [7]), .I3(GND_net), .O(n60199));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60576));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i7_2_lut (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[1][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n27996));   // verilog/coms.v(99[12:25])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[3][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n60079));
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n60176));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1316 (.I0(\data_in_frame[3][2] ), .I1(\data_in_frame[1][0] ), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1][1] ), .O(n60365));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 n71320_bdd_4_lut (.I0(n71320), .I1(n67645), .I2(n67644), .I3(byte_transmit_counter[2]), 
            .O(n71323));
    defparam n71320_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1317 (.I0(\data_in_frame[5][4] ), .I1(n60365), 
            .I2(\data_in_frame[5][5] ), .I3(GND_net), .O(n27849));
    defparam i2_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1318 (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[3]_c [4]), 
            .I2(\data_in_frame[1]_c [3]), .I3(GND_net), .O(n28009));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1318.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\data_in_frame[5][6] ), .I1(n28009), 
            .I2(GND_net), .I3(GND_net), .O(n60416));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1320 (.I0(\data_in_frame[3]_c [1]), .I1(n60545), 
            .I2(\data_in_frame[5] [3]), .I3(\data_in_frame[3][3] ), .O(n60173));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\data_in_frame[5][0] ), .I1(Kp_23__N_799), 
            .I2(GND_net), .I3(GND_net), .O(n28429));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1322 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2][5] ), .I3(GND_net), .O(n27900));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__7__I_0_4044_2_lut (.I0(\data_in_frame[0] [7]), 
            .I1(\data_in_frame[0] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_753));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_0__7__I_0_4044_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_33_lut  (.I0(n67576), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n53427), .O(n30148)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[6][3] ), .I1(\data_in_frame[6][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n28006));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60111));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1325 (.I0(\data_in_frame[5][7] ), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[4] [0]), .O(n64125));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_32_lut  (.I0(n67577), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n53426), .O(n30146)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_32  (.CI(n53426), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n53427));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_31_lut  (.I0(n67579), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n53425), .O(n30144)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_31  (.CI(n53425), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n53426));
    SB_LUT4 i1_4_lut_adj_1326 (.I0(n60576), .I1(n64129), .I2(n60199), 
            .I3(n64125), .O(n64133));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_30_lut  (.I0(n67580), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n53424), .O(n30142)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_30  (.CI(n53424), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n53425));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_29_lut  (.I0(n67581), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n53423), .O(n30140)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1327 (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[2][2] ), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[2][4] ), .O(n64147));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1328 (.I0(n28429), .I1(n60173), .I2(n60416), 
            .I3(n64133), .O(n64139));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1329 (.I0(n27849), .I1(n60142), .I2(n28435), 
            .I3(n64151), .O(n64157));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1330 (.I0(n28694), .I1(n64157), .I2(n64139), 
            .I3(n28296), .O(n54597));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60750));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_29  (.CI(n53423), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n53424));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_28_lut  (.I0(n67588), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n53422), .O(n30138)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_28  (.CI(n53422), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n53423));
    SB_LUT4 i6_4_lut_adj_1332 (.I0(n60750), .I1(n54597), .I2(n60111), 
            .I3(n60747), .O(n15_adj_5552));   // verilog/coms.v(81[16:27])
    defparam i6_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1333 (.I0(n15_adj_5552), .I1(n60296), .I2(n14_adj_5553), 
            .I3(n28435), .O(n62486));   // verilog/coms.v(81[16:27])
    defparam i8_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut (.I0(n28386), .I1(n62335), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n21_adj_5554));
    defparam i4_3_lut.LUT_INIT = 16'h4141;
    SB_LUT4 i10_4_lut_adj_1334 (.I0(n62747), .I1(n26041), .I2(n26045), 
            .I3(n62486), .O(n27_adj_5555));
    defparam i10_4_lut_adj_1334.LUT_INIT = 16'h0040;
    SB_LUT4 i9_3_lut (.I0(n4_c), .I1(n55186), .I2(n55482), .I3(GND_net), 
            .O(n26_adj_5556));
    defparam i9_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i45061_2_lut (.I0(n28559), .I1(n28041), .I2(GND_net), .I3(GND_net), 
            .O(n64318));
    defparam i45061_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45206_4_lut (.I0(n7), .I1(n28398), .I2(n28529), .I3(n55163), 
            .O(n64467));
    defparam i45206_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_27_lut  (.I0(n67591), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n53421), .O(n30136)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_27  (.CI(n53421), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n53422));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_26_lut  (.I0(n67592), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n53420), .O(n30134)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_26  (.CI(n53420), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n53421));
    SB_LUT4 i13513_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n31458));
    defparam i13513_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14_4_lut_adj_1335 (.I0(n27_adj_5555), .I1(n21_adj_5554), .I2(n27956), 
            .I3(n7_adj_5523), .O(n31_c));
    defparam i14_4_lut_adj_1335.LUT_INIT = 16'h0008;
    SB_LUT4 i16_4_lut (.I0(n31_c), .I1(n64467), .I2(n64318), .I3(n26_adj_5556), 
            .O(LED_N_3408));
    defparam i16_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_adj_1336 (.I0(\data_in_frame[21][4] ), .I1(\data_in_frame[18]_c [7]), 
            .I2(n60579), .I3(GND_net), .O(n7_adj_5557));
    defparam i2_3_lut_adj_1336.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1337 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[18][2] ), 
            .I2(n60481), .I3(GND_net), .O(n8_adj_5558));
    defparam i3_3_lut_adj_1337.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1338 (.I0(n60150), .I1(n60388), .I2(\data_in_frame[23] [4]), 
            .I3(GND_net), .O(n62764));
    defparam i2_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_LUT4 i45073_4_lut (.I0(\data_in_frame[22] [5]), .I1(n62747), .I2(n54773), 
            .I3(n55778), .O(n64331));
    defparam i45073_4_lut.LUT_INIT = 16'hdeed;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_25_lut  (.I0(n67595), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n53419), .O(n30132)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_25  (.CI(n53419), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n53420));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_24_lut  (.I0(n67596), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n53418), .O(n30130)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_24  (.CI(n53418), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n53419));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_23_lut  (.I0(n67601), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n53417), .O(n30128)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_23  (.CI(n53417), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n53418));
    SB_LUT4 n71518_bdd_4_lut (.I0(n71518), .I1(\data_out_frame[26] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[0]), 
            .O(n71521));
    defparam n71518_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1339 (.I0(n62103), .I1(n62764), .I2(n8_adj_5558), 
            .I3(\data_in_frame[22][4] ), .O(n64093));
    defparam i1_4_lut_adj_1339.LUT_INIT = 16'h4884;
    SB_LUT4 i3_4_lut_adj_1340 (.I0(\data_in_frame[22][6] ), .I1(n60458), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[20] [4]), .O(n62652));
    defparam i3_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1341 (.I0(n7_adj_5557), .I1(\data_in_frame[23] [5]), 
            .I2(\data_in_frame[21][3] ), .I3(n61855), .O(n62789));
    defparam i4_4_lut_adj_1341.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1342 (.I0(n62789), .I1(n62652), .I2(n64093), 
            .I3(n64331), .O(n64099));
    defparam i1_4_lut_adj_1342.LUT_INIT = 16'h0080;
    SB_LUT4 i4_4_lut_adj_1343 (.I0(n60257), .I1(\data_in_frame[22][1] ), 
            .I2(\data_in_frame[21] [7]), .I3(n60604), .O(n10_adj_5559));
    defparam i4_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_22_lut  (.I0(n67602), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n53416), .O(n30126)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_22  (.CI(n53416), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n53417));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_21_lut  (.I0(n67646), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n53415), .O(n30124)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_21  (.CI(n53415), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n53416));
    SB_LUT4 i1_4_lut_adj_1344 (.I0(n64099), .I1(\data_in_frame[22][0] ), 
            .I2(n8_adj_5442), .I3(\data_in_frame[19]_c [6]), .O(n64101));
    defparam i1_4_lut_adj_1344.LUT_INIT = 16'h8228;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_20_lut  (.I0(n67647), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n53414), .O(n30122)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_20  (.CI(n53414), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n53415));
    SB_LUT4 i1_4_lut_adj_1345 (.I0(\data_in_frame[17][6] ), .I1(n64101), 
            .I2(n10_adj_5559), .I3(\data_in_frame[20] [0]), .O(n64103));
    defparam i1_4_lut_adj_1345.LUT_INIT = 16'h4884;
    SB_LUT4 i3_4_lut_adj_1346 (.I0(\data_in_frame[23] [6]), .I1(\data_in_frame[21][4] ), 
            .I2(n61855), .I3(n60388), .O(n8_adj_5560));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1347 (.I0(n64103), .I1(n26003), .I2(n60260), 
            .I3(\data_in_frame[23] [7]), .O(n64105));
    defparam i1_4_lut_adj_1347.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1348 (.I0(n60512), .I1(n60579), .I2(\data_in_frame[23] [3]), 
            .I3(n60202), .O(n12_adj_5561));
    defparam i5_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1349 (.I0(n60202), .I1(n60512), .I2(\data_in_frame[18]_c [7]), 
            .I3(\data_in_frame[23] [1]), .O(n64249));
    defparam i1_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1350 (.I0(n60481), .I1(\data_in_frame[18][1] ), 
            .I2(\data_in_frame[22][3] ), .I3(n60682), .O(n10_adj_5562));
    defparam i4_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_19_lut  (.I0(n67648), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n53413), .O(n30120)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_19  (.CI(n53413), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n53414));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_18_lut  (.I0(n67649), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n53412), .O(n30118)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_18  (.CI(n53412), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n53413));
    SB_LUT4 i5_4_lut_adj_1351 (.I0(\data_in_frame[17][6] ), .I1(n60495), 
            .I2(n27873), .I3(\data_in_frame[22][2] ), .O(n12_adj_5563));
    defparam i5_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1352 (.I0(\data_in_frame[21][5] ), .I1(n64105), 
            .I2(n8_adj_5560), .I3(n26003), .O(n64107));
    defparam i1_4_lut_adj_1352.LUT_INIT = 16'h4884;
    SB_LUT4 i6_4_lut_adj_1353 (.I0(\data_in_frame[21][1] ), .I1(n12_adj_5561), 
            .I2(n60735), .I3(\data_in_frame[21]_c [2]), .O(n62338));
    defparam i6_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1354 (.I0(n27223), .I1(n12_adj_5563), .I2(n60682), 
            .I3(n54740), .O(n62155));
    defparam i6_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1355 (.I0(\data_in_frame[19][7] ), .I1(n10_adj_5562), 
            .I2(\data_in_frame[20] [1]), .I3(GND_net), .O(n62150));
    defparam i5_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1356 (.I0(n62150), .I1(n62155), .I2(n62338), 
            .I3(n64107), .O(n64113));
    defparam i1_4_lut_adj_1356.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1357 (.I0(n60601), .I1(n60443), .I2(n27264), 
            .I3(n64249), .O(n62272));
    defparam i1_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_17_lut  (.I0(n67650), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n53411), .O(n30116)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_17  (.CI(n53411), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n53412));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_16_lut  (.I0(n67651), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n53410), .O(n30114)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_16  (.CI(n53410), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n53411));
    SB_LUT4 i1_4_lut_adj_1358 (.I0(\data_in_frame[21][1] ), .I1(n64113), 
            .I2(n55671), .I3(\data_in_frame[23] [2]), .O(n64115));
    defparam i1_4_lut_adj_1358.LUT_INIT = 16'h4884;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n71512));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1359 (.I0(n62602), .I1(n55708), .I2(n60306), 
            .I3(\data_in_frame[22] [7]), .O(n64185));
    defparam i1_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1360 (.I0(n64185), .I1(n64115), .I2(n62272), 
            .I3(n55671), .O(n64119));
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'h0804;
    SB_LUT4 i1_4_lut_adj_1361 (.I0(n64119), .I1(n60443), .I2(n55671), 
            .I3(\data_in_frame[23] [0]), .O(Kp_23__N_612));
    defparam i1_4_lut_adj_1361.LUT_INIT = 16'h8228;
    SB_LUT4 i13514_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n31459));
    defparam i13514_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13515_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][0] ), 
            .I3(\Kp[0] ), .O(n31460));
    defparam i13515_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13516_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][0] ), 
            .I3(\Ki[0] ), .O(n31461));
    defparam i13516_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_15_lut  (.I0(n67659), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n53409), .O(n30112)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_15  (.CI(n53409), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n53410));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_14_lut  (.I0(n67671), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n53408), .O(n30110)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_14  (.CI(n53408), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n53409));
    SB_LUT4 n71512_bdd_4_lut (.I0(n71512), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n71515));
    defparam n71512_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14217_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n32162));
    defparam i14217_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14218_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n32163));
    defparam i14218_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14219_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n32164));
    defparam i14219_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51669_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_612), 
            .I2(LED_N_3408), .I3(Kp_23__N_1748), .O(n29831));
    defparam i51669_4_lut.LUT_INIT = 16'hc4a0;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5564), .S(n31269));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_13_lut  (.I0(n67672), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n53407), .O(n30108)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_13  (.CI(n53407), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n53408));
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [19]), .O(n44));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14220_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n32165));
    defparam i14220_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut_adj_1362 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [18]), .O(n42));   // verilog/coms.v(157[7:23])
    defparam i16_4_lut_adj_1362.LUT_INIT = 16'hfffe;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_12_lut  (.I0(n67673), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n53406), .O(n30106)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_12  (.CI(n53406), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n53407));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_11_lut  (.I0(n67676), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n53405), .O(n30104)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_11  (.CI(n53405), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n53406));
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [17]), .I3(\FRAME_MATCHER.i [8]), .O(n43));   // verilog/coms.v(157[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1363 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1363.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1364 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut_adj_1364.LUT_INIT = 16'hfffe;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_10_lut  (.I0(n67677), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n53404), .O(n30102)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_10  (.CI(n53404), .I0(n30361), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n53405));
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(157[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n69670), .I2(n67758), .I3(byte_transmit_counter_c[4]), 
            .O(n71506));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71506_bdd_4_lut (.I0(n71506), .I1(n71329), .I2(n71437), .I3(byte_transmit_counter_c[4]), 
            .O(tx_data[3]));
    defparam n71506_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52176 (.I0(byte_transmit_counter_c[3]), 
            .I1(n69637), .I2(n67745), .I3(byte_transmit_counter_c[4]), 
            .O(n71500));
    defparam byte_transmit_counter_3__bdd_4_lut_52176.LUT_INIT = 16'he4aa;
    SB_LUT4 n71500_bdd_4_lut (.I0(n71500), .I1(n71377), .I2(n71431), .I3(byte_transmit_counter_c[4]), 
            .O(tx_data[4]));
    defparam n71500_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52181 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71494));
    defparam byte_transmit_counter_0__bdd_4_lut_52181.LUT_INIT = 16'he4aa;
    SB_LUT4 n71494_bdd_4_lut (.I0(n71494), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71497));
    defparam n71494_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_9_lut  (.I0(n67678), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n53403), .O(n30100)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_9  (.CI(n53403), .I0(n30361), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n53404));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52166 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n71482));
    defparam byte_transmit_counter_0__bdd_4_lut_52166.LUT_INIT = 16'he4aa;
    SB_LUT4 n71482_bdd_4_lut (.I0(n71482), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n71485));
    defparam n71482_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52156 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n71476));
    defparam byte_transmit_counter_0__bdd_4_lut_52156.LUT_INIT = 16'he4aa;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_8_lut  (.I0(n67679), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n53402), .O(n30098)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_8  (.CI(n53402), .I0(n30361), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n53403));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_7_lut  (.I0(n67682), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n53401), .O(n30096)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_7  (.CI(n53401), .I0(n30361), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n53402));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_6_lut  (.I0(n67683), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n53400), .O(n30094)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_6  (.CI(n53400), .I0(n30361), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n53401));
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(157[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_5_lut  (.I0(n67689), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n53399), .O(n30092)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_5  (.CI(n53399), .I0(n30361), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n53400));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_4_lut  (.I0(n67690), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n53398), .O(n30090)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_4  (.CI(n53398), .I0(n30361), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n53399));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_3_lut  (.I0(n67691), .I1(n30361), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n53397), .O(n30088)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_3  (.CI(n53397), .I0(n30361), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n53398));
    SB_LUT4 \FRAME_MATCHER.i_2044_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2044_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2044_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n53397));
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [12]), .O(n45_c));   // verilog/coms.v(157[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1365 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5565), .I3(n60011), .O(n29032));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1365.LUT_INIT = 16'haaa8;
    SB_LUT4 i45353_3_lut (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64623));
    defparam i45353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14221_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n32166));
    defparam i14221_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i25_4_lut (.I0(n45_c), .I1(n50), .I2(n39), .I3(n40), .O(n27621));   // verilog/coms.v(157[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23756_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27621), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i23756_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2081));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71476_bdd_4_lut (.I0(n71476), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71479));
    defparam n71476_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14222_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n32167));
    defparam i14222_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52062 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11][6] ), 
            .I3(byte_transmit_counter[1]), .O(n71314));
    defparam byte_transmit_counter_0__bdd_4_lut_52062.LUT_INIT = 16'he4aa;
    SB_LUT4 i45354_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11][2] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64624));
    defparam i45354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45611_3_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64881));
    defparam i45611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45612_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11][5] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64882));
    defparam i45612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71314_bdd_4_lut (.I0(n71314), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8][6] ), .I3(byte_transmit_counter[1]), 
            .O(n71317));
    defparam n71314_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n31478));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i45369_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64639));
    defparam i45369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45315_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64585));
    defparam i45315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45314_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64584));
    defparam i45314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45368_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64638));
    defparam i45368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14223_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n32168));
    defparam i14223_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5566), .S(n59828));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17][0] ), .C(clk16MHz), 
           .D(n31954));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14224_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n32169));
    defparam i14224_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_3_lut_adj_1366 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[21] [6]), 
            .I2(n60782), .I3(GND_net), .O(n8_adj_5567));
    defparam i3_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_210_i3_4_lut (.I0(n54653), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5567), .I3(n60741), .O(n3_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i14225_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n32170));
    defparam i14225_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i17935_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n32171));
    defparam i17935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14227_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n32172));
    defparam i14227_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1367 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[22] [4]), 
            .I2(\data_out_frame[22] [3]), .I3(n55280), .O(n60634));
    defparam i1_4_lut_adj_1367.LUT_INIT = 16'h9669;
    SB_LUT4 i14228_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n32173));
    defparam i14228_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1368 (.I0(n54606), .I1(n54653), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n61872));
    defparam i2_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\data_out_frame[21] [6]), .I1(n54618), 
            .I2(GND_net), .I3(GND_net), .O(n60643));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1370 (.I0(n7_adj_5568), .I1(\data_out_frame[17] [5]), 
            .I2(n55614), .I3(n60775), .O(n55280));
    defparam i4_4_lut_adj_1370.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1371 (.I0(n55544), .I1(n55570), .I2(n55280), 
            .I3(GND_net), .O(n14_adj_5569));
    defparam i5_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1372 (.I0(n60643), .I1(n62106), .I2(n55641), 
            .I3(n60362), .O(n15_adj_5570));
    defparam i6_4_lut_adj_1372.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1373 (.I0(n15_adj_5570), .I1(\data_out_frame[22] [1]), 
            .I2(n14_adj_5569), .I3(n54636), .O(n62047));
    defparam i8_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n31957));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n31962));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17][3] ), .C(clk16MHz), 
           .D(n31965));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n31426));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n31429));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17][4] ), .C(clk16MHz), 
           .D(n31968));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17][5] ), .C(clk16MHz), 
           .D(n31971));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17][6] ), .C(clk16MHz), 
           .D(n31974));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17][7] ), .C(clk16MHz), 
           .D(n31977));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18][0] ), .C(clk16MHz), 
           .D(n59150));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18][1] ), .C(clk16MHz), 
           .D(n59148));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18][2] ), .C(clk16MHz), 
           .D(n59146));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18][3] ), .C(clk16MHz), 
           .D(n31990));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18][4] ), .C(clk16MHz), 
           .D(n59144));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n31996));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n59142));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18]_c [7]), .C(clk16MHz), 
           .D(n59064));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n31433));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n31437));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n59140));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19]_c [1]), .C(clk16MHz), 
           .D(n59106));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19][2] ), .C(clk16MHz), 
           .D(n59138));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19]_c [3]), .C(clk16MHz), 
           .D(n32437));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2][0] ), .C(clk16MHz), 
           .D(n31440));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19]_c [4]), .C(clk16MHz), 
           .D(n32435));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19]_c [5]), .C(clk16MHz), 
           .D(n59052));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19]_c [6]), .C(clk16MHz), 
           .D(n59118));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19][7] ), .C(clk16MHz), 
           .D(n59136));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n32038));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2][1] ), .C(clk16MHz), 
           .D(n31443));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32427));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1]_c [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n59316));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n59308));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n32418));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32415));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32412));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32409));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1374 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[22] [0]), 
            .I2(n54771), .I3(GND_net), .O(n55544));
    defparam i2_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32406));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32403));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32400));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32397));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n32041));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n59322));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n32048));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n32051));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n59214));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n32059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n32062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21][0] ), .C(clk16MHz), 
           .D(n32066));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21][1] ), .C(clk16MHz), 
           .D(n59050));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2][2] ), .C(clk16MHz), 
           .D(n31446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2][3] ), .C(clk16MHz), 
           .D(n31449));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21]_c [2]), .C(clk16MHz), 
           .D(n59046));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21][3] ), .C(clk16MHz), 
           .D(n32078));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2][4] ), .C(clk16MHz), 
           .D(n31452));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21][4] ), .C(clk16MHz), 
           .D(n32088));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2][5] ), .C(clk16MHz), 
           .D(n31455));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21][5] ), .C(clk16MHz), 
           .D(n32092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21]_c [6]), .C(clk16MHz), 
           .D(n59058));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n32098));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n59060));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22][0] ), .C(clk16MHz), 
           .D(n59062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22][1] ), .C(clk16MHz), 
           .D(n32108));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22][2] ), .C(clk16MHz), 
           .D(n32112));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22][3] ), .C(clk16MHz), 
           .D(n32115));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22][4] ), .C(clk16MHz), 
           .D(n32118));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n32351));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22][6] ), .C(clk16MHz), 
           .D(n32350));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n32349));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n32130));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n32133));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n59220));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n32140));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n32143));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n32146));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n32149));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n59230));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n31467));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n32334));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
           .D(n31482));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3]_c [1]), .C(clk16MHz), 
           .D(n31485));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n32307), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n32306), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n32305), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n32304), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n32303), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n32302), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n32301), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n32300), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n32299), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n32298), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n32297), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n32296), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n32295), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n32294), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n32293), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n32292), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n32291), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n32290), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n32289), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n32288), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n32287), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n32286), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n32285), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n32284), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n32283), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n32282), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n32281), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n32280), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n32279), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n32278), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n32277), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n32276), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n32275), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n32274), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n32273), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n32272), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n32271), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n32270), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n32269), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n32268), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n32267), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n32266), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n32265), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n32264), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n32263), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n32262), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n32261), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n32260), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n32259), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n32258), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n32257), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n32256), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n32255), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n32254), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n32253), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n32252), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n32251), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n32250), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n32249), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n32248), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n32247), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n32246), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n32245), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n32244), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n32243), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n32242), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n32241), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n32240), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n32239), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n32238), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n32237), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n32236), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n32235), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n32234), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n32233), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n32232), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
           .D(n31488));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n32229));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n32228));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n32227));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n32226));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n32225));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n32224));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n32223));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n32222));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n32221));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n32220));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n32219));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n32218));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n32217));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n32216));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n32215));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n32214));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n32213));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n32212));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n32211));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n32210));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n32209));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n32208));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n32207));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n32206));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n32205));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n32204));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n31465), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52171 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71173), .I2(n67746), .I3(byte_transmit_counter_c[4]), 
            .O(n71470));
    defparam byte_transmit_counter_3__bdd_4_lut_52171.LUT_INIT = 16'he4aa;
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n31464));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n31463));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n31462));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2889), .D(n2_adj_5571), .S(n59827));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n32203));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n32202));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n32201));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n32200));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n32199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n32198));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n32197));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n32196));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n32195));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n32194));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n32193));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n32192));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n32191));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n32190));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n32189));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n32188));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n32187));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n32186));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n32185));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n32184), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n32183), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n32182), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n32181), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n32180), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n32179), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n32178), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n32177), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n32176), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n32175), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n32174), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n32173), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n32172), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n32171), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n32170), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n32169), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n32168), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n32167), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n32166), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n32165), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n32164), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n32163), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n32162), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n31491));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3]_c [4]), .C(clk16MHz), 
           .D(n59294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3]_c [5]), .C(clk16MHz), 
           .D(n59298));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
           .D(n31500));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
           .D(n31503));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1375 (.I0(\data_out_frame[21] [7]), .I1(n55544), 
            .I2(\data_out_frame[21] [5]), .I3(GND_net), .O(n60424));
    defparam i2_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i14229_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n32174));
    defparam i14229_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n31461), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n31460), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1376 (.I0(n60782), .I1(n62106), .I2(\data_out_frame[23] [7]), 
            .I3(n55554), .O(n25812));
    defparam i3_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n31459), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n31458), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14230_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n32175));
    defparam i14230_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n31506));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1377 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60669));
    defparam i1_2_lut_adj_1377.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1378 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [1]), .I3(GND_net), .O(n60452));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_out_frame[20] [4]), .I1(n60452), 
            .I2(GND_net), .I3(GND_net), .O(n28707));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i13752_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n31697));
    defparam i13752_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n59304));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_2044__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n30088), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n30090), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n30092), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n30094), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n30096), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n30098), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n30100), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n30102), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n30104), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n30106), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n30108), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n30110), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n30112), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n30114), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n30116), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n30118), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n30120), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n30122), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n30124), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n30126), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n30128), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n30130), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n30132), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n30134), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n30136), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n30138), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n30140), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n30142), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n30144), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n30146), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2044__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n30148), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i3_4_lut_adj_1380 (.I0(n62354), .I1(n28707), .I2(n28330), 
            .I3(\data_out_frame[20] [5]), .O(n54936));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1380.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1381 (.I0(\data_out_frame[15] [3]), .I1(n60185), 
            .I2(n27799), .I3(GND_net), .O(n54771));
    defparam i2_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 i13749_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n31694));
    defparam i13749_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14231_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n32176));
    defparam i14231_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n31512));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1382 (.I0(n54771), .I1(\data_out_frame[19] [5]), 
            .I2(n62117), .I3(GND_net), .O(n55554));
    defparam i1_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n31515));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n31518));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n31521));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n31524));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n31527));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13746_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n31691));
    defparam i13746_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5][0] ), .C(clk16MHz), 
           .D(n31530));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13760_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n31705));
    defparam i13760_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5][1] ), .C(clk16MHz), 
           .D(n31533));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14232_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n32177));
    defparam i14232_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14233_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n32178));
    defparam i14233_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1383 (.I0(\data_out_frame[16] [3]), .I1(n54982), 
            .I2(n60241), .I3(GND_net), .O(n60478));
    defparam i1_3_lut_adj_1383.LUT_INIT = 16'h6969;
    SB_LUT4 i13743_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n31688));
    defparam i13743_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_789_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13680_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n31625));
    defparam i13680_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5][2] ), .C(clk16MHz), 
           .D(n31536));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1384 (.I0(n60625), .I1(n60182), .I2(\data_out_frame[11][1] ), 
            .I3(n60717), .O(n10_adj_5572));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i13641_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n31586));
    defparam i13641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13638_3_lut_4_lut (.I0(n167), .I1(n60032), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n31583));
    defparam i13638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1385 (.I0(n60230), .I1(n27799), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5573));
    defparam i1_2_lut_adj_1385.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1386 (.I0(\data_out_frame[17] [5]), .I1(n5_adj_5573), 
            .I2(\data_out_frame[15] [3]), .I3(n55614), .O(n54618));
    defparam i1_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 i14234_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n32179));
    defparam i14234_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_out_frame[19] [3]), .I1(n54618), 
            .I2(GND_net), .I3(GND_net), .O(n60345));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1388 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27913));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1388.LUT_INIT = 16'h6666;
    SB_LUT4 i16_4_lut_adj_1389 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(n54752), .I3(\data_out_frame[17] [2]), .O(n40_adj_5574));
    defparam i16_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1390 (.I0(n27913), .I1(\data_out_frame[18] [7]), 
            .I2(n60281), .I3(\data_out_frame[19] [4]), .O(n38));
    defparam i14_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1391 (.I0(n60345), .I1(\data_out_frame[19] [6]), 
            .I2(n60241), .I3(\data_out_frame[16] [5]), .O(n39_adj_5575));
    defparam i15_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1392 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[18] [2]), 
            .I2(n60637), .I3(n60054), .O(n37));
    defparam i13_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1393 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[17] [3]), 
            .I2(n60342), .I3(\data_out_frame[17] [6]), .O(n42_adj_5576));
    defparam i18_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 select_791_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n1_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39_adj_5575), .I2(n38), .I3(n40_adj_5574), 
            .O(n46));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1394 (.I0(n55614), .I1(n55303), .I2(n60145), 
            .I3(\data_out_frame[17] [1]), .O(n41_adj_5577));
    defparam i17_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut (.I0(n41_adj_5577), .I1(n46), .I2(n42_adj_5576), 
            .I3(GND_net), .O(n60679));
    defparam i23_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1395 (.I0(n60679), .I1(n60446), .I2(n28864), 
            .I3(n55719), .O(n13_adj_5578));
    defparam i5_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1396 (.I0(n13_adj_5578), .I1(n11_adj_5579), .I2(n62514), 
            .I3(n54578), .O(n62354));
    defparam i7_4_lut_adj_1396.LUT_INIT = 16'h9669;
    SB_LUT4 i14235_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n32180));
    defparam i14235_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14236_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n32181));
    defparam i14236_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1397 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[11][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5580));
    defparam i1_2_lut_adj_1397.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1398 (.I0(n60625), .I1(n60325), .I2(n60729), 
            .I3(n6_adj_5580), .O(n60230));
    defparam i4_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 n71470_bdd_4_lut (.I0(n71470), .I1(n71365), .I2(n7_adj_5581), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n71470_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1399 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60054));
    defparam i1_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i14237_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n32182));
    defparam i14237_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1400 (.I0(n60775), .I1(n60595), .I2(n60230), 
            .I3(n6_adj_5582), .O(n54636));
    defparam i4_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1401 (.I0(n55303), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60595));
    defparam i1_2_lut_adj_1401.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\data_out_frame[19] [7]), .I1(n60145), 
            .I2(GND_net), .I3(GND_net), .O(n60568));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h6666;
    SB_LUT4 i45051_3_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [6]), .I3(n28435), .O(n64308));   // verilog/coms.v(80[16:27])
    defparam i45051_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i2_3_lut_adj_1403 (.I0(n54638), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[15] [2]), .I3(GND_net), .O(n60185));
    defparam i2_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1404 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [5]), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1404.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1405 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(Kp_23__N_767), .I3(\data_in_frame[1][0] ), .O(n28296));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1406 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n60410), .I3(n6_c), .O(n55105));
    defparam i4_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1407 (.I0(\data_out_frame[18] [1]), .I1(n60352), 
            .I2(n55105), .I3(GND_net), .O(n55641));
    defparam i2_3_lut_adj_1407.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1408 (.I0(n60568), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[20] [0]), .I3(n60595), .O(n10_adj_5583));
    defparam i4_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1409 (.I0(n60185), .I1(n10_adj_5583), .I2(\data_out_frame[22] [2]), 
            .I3(GND_net), .O(n55690));
    defparam i5_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1410 (.I0(n28889), .I1(n60349), .I2(n37_adj_5584), 
            .I3(\data_out_frame[15] [7]), .O(n55645));
    defparam i3_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1411 (.I0(n28169), .I1(n60290), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n37_adj_5584));
    defparam i2_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_out_frame[13] [7]), .I1(n54789), 
            .I2(GND_net), .I3(GND_net), .O(n60349));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1413 (.I0(n60640), .I1(n60161), .I2(n28198), 
            .I3(\data_out_frame[11][7] ), .O(n18_adj_5585));
    defparam i7_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1414 (.I0(n27770), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5586));
    defparam i5_2_lut_adj_1414.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1415 (.I0(\data_out_frame[8][2] ), .I1(n18_adj_5585), 
            .I2(\data_out_frame[14] [1]), .I3(\data_out_frame[10] [4]), 
            .O(n20_adj_5587));
    defparam i9_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1416 (.I0(n60753), .I1(n20_adj_5587), .I2(n16_adj_5586), 
            .I3(n60349), .O(n62514));
    defparam i10_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1417 (.I0(n37_adj_5584), .I1(n45_adj_5588), .I2(n20_adj_5589), 
            .I3(GND_net), .O(n60322));
    defparam i2_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1418 (.I0(n55703), .I1(n60322), .I2(n62514), 
            .I3(\data_out_frame[16] [2]), .O(n55659));
    defparam i3_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1419 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [2]), 
            .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1419.LUT_INIT = 16'ha088;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_out_frame[9] [2]), .I1(n60729), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5590));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1421 (.I0(n1130), .I1(n28188), .I2(n60565), .I3(n6_adj_5590), 
            .O(n45_adj_5588));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1422 (.I0(\data_out_frame[6] [7]), .I1(n60328), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[4] [5]), .O(n12_adj_5591));
    defparam i5_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1423 (.I0(\data_out_frame[7] [1]), .I1(n12_adj_5591), 
            .I2(\data_out_frame[11][5] ), .I3(n60244), .O(n54789));
    defparam i6_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1424 (.I0(n54789), .I1(n45_adj_5588), .I2(GND_net), 
            .I3(GND_net), .O(n60410));
    defparam i1_2_lut_adj_1424.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\data_out_frame[16] [1]), .I1(n55645), 
            .I2(GND_net), .I3(GND_net), .O(n55703));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1426 (.I0(\data_out_frame[16] [0]), .I1(n1835), 
            .I2(n7_adj_5592), .I3(n8_adj_5593), .O(n60352));
    defparam i2_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\data_out_frame[18] [3]), .I1(n55659), 
            .I2(GND_net), .I3(GND_net), .O(n55770));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(\data_out_frame[20] [7]), .I1(n62354), 
            .I2(GND_net), .I3(GND_net), .O(n60076));
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1429 (.I0(\data_out_frame[20] [5]), .I1(n55776), 
            .I2(GND_net), .I3(GND_net), .O(n55625));
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h9999;
    SB_LUT4 i14238_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n32183));
    defparam i14238_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1430 (.I0(\data_out_frame[22] [1]), .I1(n55690), 
            .I2(n55627), .I3(n6_adj_5594), .O(n55550));
    defparam i4_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1431 (.I0(n55663), .I1(\data_out_frame[20] [0]), 
            .I2(n60449), .I3(n55554), .O(n55570));
    defparam i1_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1432 (.I0(\data_out_frame[21] [7]), .I1(n55570), 
            .I2(n55550), .I3(n55625), .O(n55739));
    defparam i3_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i14239_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n32184));
    defparam i14239_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1433 (.I0(n61872), .I1(n60635), .I2(GND_net), 
            .I3(GND_net), .O(n60464));
    defparam i1_2_lut_adj_1433.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5296));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(\data_out_frame[22] [4]), .I1(n55627), 
            .I2(GND_net), .I3(GND_net), .O(n60073));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h9999;
    SB_LUT4 i13520_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n31465));
    defparam i13520_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1435 (.I0(n60073), .I1(n60464), .I2(n62640), 
            .I3(n55739), .O(n12_adj_5595));
    defparam i5_4_lut_adj_1435.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_209_i3_4_lut (.I0(n62047), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5595), .I3(n8_adj_5596), .O(n3_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_209_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_791_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n1_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i18677_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n32232));
    defparam i18677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14288_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n32233));
    defparam i14288_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18710_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n32234));
    defparam i18710_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14290_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n32235));
    defparam i14290_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14291_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n32236));
    defparam i14291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(reset), .I1(n3491), .I2(GND_net), .I3(GND_net), 
            .O(n60002));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14292_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n32237));
    defparam i14292_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13649_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n31594));   // verilog/coms.v(130[12] 305[6])
    defparam i13649_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1437 (.I0(\data_out_frame[18] [3]), .I1(n55659), 
            .I2(n60352), .I3(\data_out_frame[20] [4]), .O(n55776));
    defparam i1_2_lut_3_lut_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1438 (.I0(\data_out_frame[18] [3]), .I1(n55659), 
            .I2(n60352), .I3(n54936), .O(n60362));
    defparam i1_2_lut_3_lut_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n39975));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'hdddd;
    SB_LUT4 i13533_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n31478));   // verilog/coms.v(130[12] 305[6])
    defparam i13533_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13650_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n31595));   // verilog/coms.v(130[12] 305[6])
    defparam i13650_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14293_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n32238));
    defparam i14293_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14294_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n32239));
    defparam i14294_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13651_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n31596));   // verilog/coms.v(130[12] 305[6])
    defparam i13651_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14295_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][7] ), 
            .I3(\Ki[7] ), .O(n32240));
    defparam i14295_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13652_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n31597));   // verilog/coms.v(130[12] 305[6])
    defparam i13652_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14296_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][6] ), 
            .I3(\Ki[6] ), .O(n32241));
    defparam i14296_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13653_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n31598));   // verilog/coms.v(130[12] 305[6])
    defparam i13653_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1440 (.I0(n28963), .I1(n54578), .I2(GND_net), 
            .I3(GND_net), .O(n55561));
    defparam i1_2_lut_adj_1440.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1441 (.I0(n61989), .I1(n28963), .I2(\data_out_frame[17] [0]), 
            .I3(GND_net), .O(n60342));
    defparam i2_3_lut_adj_1441.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1442 (.I0(\data_out_frame[19] [1]), .I1(n60616), 
            .I2(n28864), .I3(n60268), .O(n12_adj_5597));
    defparam i5_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1443 (.I0(\data_out_frame[18] [7]), .I1(n12_adj_5597), 
            .I2(\data_out_frame[19] [0]), .I3(n60342), .O(n60446));
    defparam i6_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i14297_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][5] ), 
            .I3(\Ki[5] ), .O(n32242));
    defparam i14297_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13654_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n31599));   // verilog/coms.v(130[12] 305[6])
    defparam i13654_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1444 (.I0(Kp_23__N_753), .I1(n60515), .I2(n60272), 
            .I3(\data_in_frame[0] [3]), .O(Kp_23__N_748));   // verilog/coms.v(73[16:62])
    defparam i3_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i14298_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][4] ), 
            .I3(\Ki[4] ), .O(n32243));
    defparam i14298_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1445 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n60211));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1445.LUT_INIT = 16'h6666;
    SB_LUT4 i13655_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n31600));   // verilog/coms.v(130[12] 305[6])
    defparam i13655_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(n54982), .I1(n60446), .I2(GND_net), 
            .I3(GND_net), .O(n28869));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1447 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60797));
    defparam i1_2_lut_adj_1447.LUT_INIT = 16'h6666;
    SB_LUT4 i45617_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64887));
    defparam i45617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1448 (.I0(\data_out_frame[17] [1]), .I1(n54585), 
            .I2(n60153), .I3(\data_out_frame[16] [7]), .O(n60490));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i45618_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64888));
    defparam i45618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45639_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64909));
    defparam i45639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45638_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64908));
    defparam i45638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1449 (.I0(n60521), .I1(n60809), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[10] [0]), .O(n10_adj_5598));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1450 (.I0(n60066), .I1(n10_adj_5598), .I2(\data_out_frame[12] [3]), 
            .I3(GND_net), .O(n28963));   // verilog/coms.v(77[16:27])
    defparam i5_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(n27770), .I1(\data_out_frame[8][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5599));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i13656_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n31601));   // verilog/coms.v(130[12] 305[6])
    defparam i13656_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13657_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n31602));   // verilog/coms.v(130[12] 305[6])
    defparam i13657_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1452 (.I0(n27774), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[5] [7]), .I3(n6_adj_5599), .O(n60530));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i13658_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n31603));   // verilog/coms.v(130[12] 305[6])
    defparam i13658_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14299_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n32244));
    defparam i14299_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(\data_out_frame[8][3] ), .I1(n28169), 
            .I2(GND_net), .I3(GND_net), .O(n60640));
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i45452_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64722));
    defparam i45452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45453_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64723));
    defparam i45453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1454 (.I0(n60711), .I1(n28524), .I2(n28620), 
            .I3(\data_out_frame[10] [7]), .O(n12_adj_5600));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i45351_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64621));
    defparam i45351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13659_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n31604));   // verilog/coms.v(130[12] 305[6])
    defparam i13659_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i45350_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64620));
    defparam i45350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45428_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64698));
    defparam i45428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45429_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64699));
    defparam i45429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45441_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64711));
    defparam i45441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45440_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64710));
    defparam i45440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1455 (.I0(\data_out_frame[10] [1]), .I1(n12_adj_5600), 
            .I2(\data_out_frame[10] [5]), .I3(n62456), .O(n62385));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 i45335_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64605));
    defparam i45335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13660_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n31605));   // verilog/coms.v(130[12] 305[6])
    defparam i13660_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_4_lut_adj_1456 (.I0(n61660), .I1(n60711), .I2(n28347), 
            .I3(n60530), .O(n12_adj_5601));
    defparam i5_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i45336_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64606));
    defparam i45336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45348_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64618));
    defparam i45348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_748), .I3(GND_net), .O(n55167));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i45347_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64617));
    defparam i45347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45641_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64911));
    defparam i45641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45642_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64912));
    defparam i45642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45633_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64903));
    defparam i45633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1458 (.I0(n27767), .I1(n12_adj_5601), .I2(n62385), 
            .I3(n60640), .O(n55614));
    defparam i6_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1459 (.I0(n60170), .I1(n28864), .I2(n60490), 
            .I3(\data_out_frame[19] [3]), .O(n55706));
    defparam i1_2_lut_3_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1460 (.I0(n60705), .I1(n1191), .I2(\data_out_frame[12] [6]), 
            .I3(n60708), .O(n10_adj_5602));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1461 (.I0(n60530), .I1(n10_adj_5602), .I2(\data_out_frame[8][2] ), 
            .I3(GND_net), .O(n54585));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i45632_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64902));
    defparam i45632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2][4] ), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n27907));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i13661_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n31606));   // verilog/coms.v(130[12] 305[6])
    defparam i13661_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13662_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n31607));   // verilog/coms.v(130[12] 305[6])
    defparam i13662_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13679_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n31624));   // verilog/coms.v(130[12] 305[6])
    defparam i13679_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1463 (.I0(\data_out_frame[21] [2]), .I1(n54982), 
            .I2(n60446), .I3(\data_out_frame[20] [7]), .O(n9));
    defparam i1_2_lut_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1464 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[4] [6]), .O(n28188));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1465 (.I0(n60708), .I1(\data_out_frame[10] [4]), 
            .I2(n1516), .I3(n60533), .O(n28198));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i13678_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n31623));   // verilog/coms.v(130[12] 305[6])
    defparam i13678_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13677_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n31622));   // verilog/coms.v(130[12] 305[6])
    defparam i13677_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13676_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n31621));   // verilog/coms.v(130[12] 305[6])
    defparam i13676_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13675_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n31620));   // verilog/coms.v(130[12] 305[6])
    defparam i13675_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1466 (.I0(n28198), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[12] [4]), 
            .O(n28864));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n59968));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1467 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26][1] ), 
            .O(n59967));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1467.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1468 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26][2] ), 
            .O(n59966));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1468.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1469 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n59965));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1469.LUT_INIT = 16'h5100;
    SB_LUT4 i3_4_lut_adj_1470 (.I0(\data_out_frame[15] [1]), .I1(n54638), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [2]), 
            .O(n60170));
    defparam i3_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i13674_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n31619));   // verilog/coms.v(130[12] 305[6])
    defparam i13674_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1471 (.I0(n60170), .I1(n28864), .I2(GND_net), 
            .I3(GND_net), .O(n28205));
    defparam i1_2_lut_adj_1471.LUT_INIT = 16'h6666;
    SB_LUT4 i48733_2_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67616));
    defparam i48733_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48690_2_lut (.I0(\data_out_frame[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67617));
    defparam i48690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5603));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_adj_5604));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45320_3_lut (.I0(\data_out_frame[8][1] ), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64590));
    defparam i45320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45321_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11][1] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64591));
    defparam i45321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1472 (.I0(\data_out_frame[17] [3]), .I1(n54585), 
            .I2(n55614), .I3(n60385), .O(n62117));
    defparam i3_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1473 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5295));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1473.LUT_INIT = 16'ha088;
    SB_LUT4 i45630_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64900));
    defparam i45630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45629_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64899));
    defparam i45629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5605));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48727_2_lut (.I0(\data_out_frame[3][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67615));
    defparam i48727_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5606));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i4_3_lut (.I0(\data_out_frame[4] [3]), 
            .I1(\data_out_frame[5] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_adj_5607));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12127_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30071));   // verilog/coms.v(109[34:55])
    defparam i12127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18632_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][2] ), 
            .I3(\Ki[2] ), .O(n32245));
    defparam i18632_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13673_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n31618));   // verilog/coms.v(130[12] 305[6])
    defparam i13673_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i45600_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64870));
    defparam i45600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45601_4_lut (.I0(n64870), .I1(n30071), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64871));
    defparam i45601_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45599_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64869));
    defparam i45599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13672_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n31617));   // verilog/coms.v(130[12] 305[6])
    defparam i13672_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i49495_2_lut (.I0(n71389), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67755));
    defparam i49495_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_789_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5294));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i49243_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67741));
    defparam i49243_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1474 (.I0(n62117), .I1(\data_out_frame[19] [4]), 
            .I2(n28205), .I3(GND_net), .O(n62106));
    defparam i2_3_lut_adj_1474.LUT_INIT = 16'h6969;
    SB_LUT4 i45393_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64663));
    defparam i45393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1475 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n59964));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1475.LUT_INIT = 16'h5100;
    SB_LUT4 i45394_4_lut (.I0(n64663), .I1(n67741), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n64664));
    defparam i45394_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i45392_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64662));
    defparam i45392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1476 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n59962));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1476.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1477 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n59963));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1477.LUT_INIT = 16'h5100;
    SB_LUT4 i18656_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5][1] ), 
            .I3(\Ki[1] ), .O(n32246));
    defparam i18656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1478 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n59970));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1478.LUT_INIT = 16'h5100;
    SB_LUT4 i4_4_lut_adj_1479 (.I0(\data_out_frame[21] [4]), .I1(n28963), 
            .I2(n60170), .I3(n6_adj_5608), .O(n54653));
    defparam i4_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i48965_2_lut (.I0(n71401), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67743));
    defparam i48965_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45435_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64705));
    defparam i45435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45436_4_lut (.I0(n64705), .I1(n30156), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n64706));
    defparam i45436_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i45434_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64704));
    defparam i45434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13671_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n31616));   // verilog/coms.v(130[12] 305[6])
    defparam i13671_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(\data_out_frame[21] [5]), .I1(n62106), 
            .I2(GND_net), .I3(GND_net), .O(n60391));
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h9999;
    SB_LUT4 i49026_2_lut (.I0(n71383), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67730));
    defparam i49026_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12083_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30026));   // verilog/coms.v(109[34:55])
    defparam i12083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45411_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64681));
    defparam i45411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45412_4_lut (.I0(n64681), .I1(n30026), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64682));
    defparam i45412_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45410_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64680));
    defparam i45410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1481 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n59956));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1481.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1482 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27][1] ), 
            .O(n59961));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1482.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1483 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n60565));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1483.LUT_INIT = 16'h6666;
    SB_LUT4 i49311_2_lut (.I0(n71515), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67742));
    defparam i49311_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12081_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30024));   // verilog/coms.v(109[34:55])
    defparam i12081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45408_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64678));
    defparam i45408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1484 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27][2] ), 
            .O(n59957));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1484.LUT_INIT = 16'h5100;
    SB_LUT4 select_789_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45409_4_lut (.I0(n64678), .I1(n30024), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64679));
    defparam i45409_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45407_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64677));
    defparam i45407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1485 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n59958));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1485.LUT_INIT = 16'h5100;
    SB_LUT4 i24203125_i1_3_lut (.I0(n71317), .I1(n71485), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_5609));
    defparam i24203125_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1486 (.I0(\data_out_frame[13] [5]), .I1(n28714), 
            .I2(n8_adj_5610), .I3(n60139), .O(n28889));
    defparam i1_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1487 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n60153));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1488 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n59955));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1488.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1489 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n59959));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1489.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(\data_out_frame[6] [1]), .I1(n27770), 
            .I2(GND_net), .I3(GND_net), .O(n27767));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[8][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n60573));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 i45644_3_lut (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64914));
    defparam i45644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1492 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n28714));
    defparam i2_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i11_3_lut_adj_1493 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n38_adj_5611));
    defparam i11_3_lut_adj_1493.LUT_INIT = 16'h9696;
    SB_LUT4 i18_4_lut_adj_1494 (.I0(\data_out_frame[4] [5]), .I1(n60196), 
            .I2(\data_out_frame[7] [6]), .I3(n28918), .O(n45_adj_5612));
    defparam i18_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i18921_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n32247));
    defparam i18921_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15_4_lut_adj_1495 (.I0(n60598), .I1(n60744), .I2(\data_out_frame[7] [5]), 
            .I3(\data_out_frame[9] [7]), .O(n42_adj_5613));
    defparam i15_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i45645_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11][4] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64915));
    defparam i45645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1496 (.I0(n3491), .I1(n161), .I2(\FRAME_MATCHER.i[0] ), 
            .I3(n1), .O(n144));
    defparam i3_4_lut_adj_1496.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1497 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n59960));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1497.LUT_INIT = 16'h5100;
    SB_LUT4 i17_4_lut_adj_1498 (.I0(n60062), .I1(n60108), .I2(n60573), 
            .I3(\data_out_frame[5] [4]), .O(n44_adj_5615));
    defparam i17_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n45_adj_5612), .I1(\data_out_frame[5] [5]), .I2(n38_adj_5611), 
            .I3(n27767), .O(n50_adj_5616));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i48969_2_lut (.I0(n10_adj_5617), .I1(n144), .I2(GND_net), 
            .I3(GND_net), .O(n67722));   // verilog/coms.v(94[13:20])
    defparam i48969_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i22131_4_lut (.I0(n163), .I1(n67722), .I2(rx_data[3]), .I3(\data_in_frame[14]_c [3]), 
            .O(n40004));   // verilog/coms.v(94[13:20])
    defparam i22131_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22132_3_lut (.I0(n40004), .I1(\data_in_frame[14]_c [3]), .I2(reset), 
            .I3(GND_net), .O(n31886));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14303_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n32248));
    defparam i14303_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14304_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][5] ), 
            .I3(\Kp[13] ), .O(n32249));
    defparam i14304_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1499 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n59969));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1499.LUT_INIT = 16'h5100;
    SB_LUT4 i21_4_lut (.I0(n28714), .I1(n42_adj_5613), .I2(\data_out_frame[9] [1]), 
            .I3(\data_out_frame[7] [2]), .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14305_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][4] ), 
            .I3(\Kp[12] ), .O(n32250));
    defparam i14305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13670_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n31615));   // verilog/coms.v(130[12] 305[6])
    defparam i13670_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22_4_lut_adj_1500 (.I0(n28524), .I1(n44_adj_5615), .I2(n32), 
            .I3(n1182), .O(n49));
    defparam i22_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i14306_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][3] ), 
            .I3(\Kp[11] ), .O(n32251));
    defparam i14306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[4] [7]), .I3(\data_out_frame[4] [4]), .O(n47));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13669_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n31614));   // verilog/coms.v(130[12] 305[6])
    defparam i13669_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14307_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][2] ), 
            .I3(\Kp[10] ), .O(n32252));
    defparam i14307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i26_4_lut (.I0(n47), .I1(n49), .I2(n48), .I3(n50_adj_5616), 
            .O(n62456));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1501 (.I0(\data_out_frame[13] [1]), .I1(n62456), 
            .I2(n28714), .I3(GND_net), .O(n60788));
    defparam i2_3_lut_adj_1501.LUT_INIT = 16'h6969;
    SB_LUT4 i14308_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][1] ), 
            .I3(\Kp[9] ), .O(n32253));
    defparam i14308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1502 (.I0(\data_in_frame[2][3] ), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n28435));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1502.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5589));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1504 (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[8][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n60182));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1504.LUT_INIT = 16'h6666;
    SB_LUT4 i13668_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n31613));   // verilog/coms.v(130[12] 305[6])
    defparam i13668_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13667_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n31612));   // verilog/coms.v(130[12] 305[6])
    defparam i13667_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1505 (.I0(n1191), .I1(\data_out_frame[12] [7]), 
            .I2(n60108), .I3(n60156), .O(n15_adj_5618));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1506 (.I0(n15_adj_5618), .I1(\data_out_frame[6] [0]), 
            .I2(n14_adj_5619), .I3(\data_out_frame[8][3] ), .O(n54638));   // verilog/coms.v(88[17:28])
    defparam i8_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1507 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60244));
    defparam i1_2_lut_adj_1507.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60717));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 i14309_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][0] ), 
            .I3(\Kp[8] ), .O(n32254));
    defparam i14309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1509 (.I0(\data_out_frame[8][4] ), .I1(n27774), 
            .I2(n60553), .I3(n6_adj_5620), .O(n60325));
    defparam i4_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i14310_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [7]), 
            .I3(\Kp[7] ), .O(n32255));
    defparam i14310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60637));
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i14311_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [6]), 
            .I3(\Kp[6] ), .O(n32256));
    defparam i14311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1511 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n60705));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1511.LUT_INIT = 16'h9696;
    SB_LUT4 i14312_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [5]), 
            .I3(\Kp[5] ), .O(n32257));
    defparam i14312_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1512 (.I0(\data_out_frame[8][6] ), .I1(n60156), 
            .I2(GND_net), .I3(GND_net), .O(n28769));
    defparam i1_2_lut_adj_1512.LUT_INIT = 16'h6666;
    SB_LUT4 i18819_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [4]), 
            .I3(\Kp[4] ), .O(n32258));
    defparam i18819_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1513 (.I0(\data_out_frame[4] [6]), .I1(n60214), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n28445));
    defparam i2_3_lut_adj_1513.LUT_INIT = 16'h9696;
    SB_LUT4 i14314_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][3] ), 
            .I3(\Kp[3] ), .O(n32259));
    defparam i14314_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60196));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27763));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14315_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][2] ), 
            .I3(\Kp[2] ), .O(n32260));
    defparam i14315_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5621));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1517 (.I0(n1191), .I1(n27763), .I2(n60316), .I3(n6_adj_5621), 
            .O(n60214));   // verilog/coms.v(74[16:62])
    defparam i4_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i18874_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [1]), 
            .I3(\Kp[1] ), .O(n32261));
    defparam i18874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1518 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n60156));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1518.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[8][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n60082));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1520 (.I0(n27774), .I1(n60156), .I2(\data_out_frame[8][5] ), 
            .I3(GND_net), .O(n28524));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1520.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60553));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1522 (.I0(n60214), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n60125));
    defparam i2_3_lut_adj_1522.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1523 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60598));
    defparam i1_2_lut_adj_1523.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1524 (.I0(n60139), .I1(n60556), .I2(\data_out_frame[13] [4]), 
            .I3(n28769), .O(n12_adj_5622));
    defparam i5_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1525 (.I0(\data_out_frame[11][2] ), .I1(n12_adj_5622), 
            .I2(n60598), .I3(\data_out_frame[8][7] ), .O(n55303));
    defparam i6_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60385));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1527 (.I0(n60125), .I1(n60553), .I2(n28524), 
            .I3(n60082), .O(n12_adj_5623));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1528 (.I0(\data_out_frame[11][2] ), .I1(n12_adj_5623), 
            .I2(n60714), .I3(n28445), .O(n62204));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i14317_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n32262));
    defparam i14317_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13666_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n31611));   // verilog/coms.v(130[12] 305[6])
    defparam i13666_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1529 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[16] [0]), 
            .I2(n62204), .I3(n55303), .O(n60381));
    defparam i1_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1530 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [5]), .I3(GND_net), .O(n60145));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1530.LUT_INIT = 16'h9696;
    SB_LUT4 i13665_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n31610));   // verilog/coms.v(130[12] 305[6])
    defparam i13665_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14318_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n32263));
    defparam i14318_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60556));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i13664_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n31609));   // verilog/coms.v(130[12] 305[6])
    defparam i13664_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13663_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n31608));   // verilog/coms.v(130[12] 305[6])
    defparam i13663_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1532 (.I0(\data_out_frame[7] [6]), .I1(n60778), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[12] [0]), .O(n60161));
    defparam i3_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i394_2_lut (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1182));   // verilog/coms.v(78[16:27])
    defparam i394_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1533 (.I0(n28188), .I1(\data_out_frame[11][6] ), 
            .I2(\data_out_frame[4] [7]), .I3(n6_adj_5624), .O(n60290));
    defparam i4_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1534 (.I0(\data_out_frame[14] [2]), .I1(n60610), 
            .I2(n60161), .I3(\data_out_frame[12] [1]), .O(n10_adj_5625));
    defparam i4_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i14319_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n32264));
    defparam i14319_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_3_lut_adj_1535 (.I0(n60290), .I1(n10_adj_5625), .I2(n1182), 
            .I3(GND_net), .O(n54578));
    defparam i5_3_lut_adj_1535.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60812));
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut_adj_1537 (.I0(\data_out_frame[6] [1]), .I1(n54578), 
            .I2(GND_net), .I3(GND_net), .O(n28_adj_5626));
    defparam i5_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i14320_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n32265));
    defparam i14320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15_4_lut_adj_1538 (.I0(n29000), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[11][5] ), .I3(\data_out_frame[4] [0]), .O(n38_adj_5627));
    defparam i15_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i14321_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n32266));
    defparam i14321_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13_4_lut_adj_1539 (.I0(n60705), .I1(n60637), .I2(n60744), 
            .I3(n60325), .O(n36));
    defparam i13_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1540 (.I0(n54638), .I1(n38_adj_5627), .I2(n28_adj_5626), 
            .I3(\data_out_frame[11][3] ), .O(n42_adj_5628));
    defparam i19_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1541 (.I0(\data_out_frame[14] [0]), .I1(n60788), 
            .I2(n55303), .I3(n60714), .O(n40_adj_5629));
    defparam i17_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1542 (.I0(n60675), .I1(n36), .I2(n60048), .I3(n60812), 
            .O(n41_adj_5630));
    defparam i18_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1543 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[14] [6]), 
            .I2(n20_adj_5589), .I3(\data_out_frame[11][7] ), .O(n39_adj_5631));
    defparam i16_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1544 (.I0(n39_adj_5631), .I1(n41_adj_5630), .I2(n40_adj_5629), 
            .I3(n42_adj_5628), .O(n62609));
    defparam i22_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i14322_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n32267));
    defparam i14322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1545 (.I0(n60153), .I1(n28889), .I2(n1835), .I3(n62609), 
            .O(n10_adj_5632));
    defparam i4_4_lut_adj_1545.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1546 (.I0(n60145), .I1(n60381), .I2(n10_adj_5632), 
            .I3(n60385), .O(n28303));
    defparam i1_4_lut_adj_1546.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1547 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n60044), .O(n30400));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1547.LUT_INIT = 16'hfffd;
    SB_LUT4 i14323_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n32268));
    defparam i14323_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1548 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[8][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n60753));
    defparam i1_2_lut_adj_1548.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60521));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1550 (.I0(n60066), .I1(n60527), .I2(GND_net), 
            .I3(GND_net), .O(n60048));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1550.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60533));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5633));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1553 (.I0(n60048), .I1(\data_out_frame[10] [1]), 
            .I2(n60521), .I3(n6_adj_5633), .O(n60281));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1554 (.I0(n60455), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [0]), .I3(n60533), .O(n10_adj_5634));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1555 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n60036), .O(n60042));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1555.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_1556 (.I0(n1516), .I1(n60281), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n1655));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1556.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1557 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n60778));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1557.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1558 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60675));
    defparam i1_2_lut_adj_1558.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1559 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28347));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1559.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1560 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n60164));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1561 (.I0(\data_out_frame[9] [5]), .I1(n60164), 
            .I2(\data_out_frame[4] [7]), .I3(\data_out_frame[5] [1]), .O(n28169));   // verilog/coms.v(76[16:34])
    defparam i3_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(\data_out_frame[10] [0]), .I1(n28169), 
            .I2(GND_net), .I3(GND_net), .O(n28620));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1563 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60316));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1563.LUT_INIT = 16'h6666;
    SB_LUT4 i14324_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n32269));
    defparam i14324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14325_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n32270));
    defparam i14325_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60527));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[11][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5635));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1566 (.I0(n60527), .I1(n60316), .I2(n60610), 
            .I3(n6_adj_5635), .O(n54752));   // verilog/coms.v(74[16:62])
    defparam i4_4_lut_adj_1566.LUT_INIT = 16'h6996;
    SB_LUT4 i14326_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n32271));
    defparam i14326_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1567 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60455));
    defparam i1_2_lut_adj_1567.LUT_INIT = 16'h6666;
    SB_LUT4 i14327_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n32272));
    defparam i14327_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1568 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n60036), .O(n60039));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1568.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52146 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71179), .I2(n67759), .I3(byte_transmit_counter_c[4]), 
            .O(n71464));
    defparam byte_transmit_counter_3__bdd_4_lut_52146.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1569 (.I0(\data_out_frame[16] [5]), .I1(n60268), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n28021));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1569.LUT_INIT = 16'h9696;
    SB_LUT4 i12212_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n30156));   // verilog/coms.v(109[34:55])
    defparam i12212_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut_adj_1570 (.I0(n60455), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[14] [3]), .I3(n54752), .O(n10_adj_5636));
    defparam i4_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 equal_297_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n8_adj_5637));   // verilog/coms.v(157[7:23])
    defparam equal_297_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1571 (.I0(n60616), .I1(n29000), .I2(n55719), 
            .I3(n28021), .O(n61989));
    defparam i3_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i14328_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n32273));
    defparam i14328_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n59220));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1572 (.I0(\data_in_frame[16] [5]), .I1(n61729), 
            .I2(n60190), .I3(n60278), .O(n64089));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1572.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1573 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n27595), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n4_adj_5638));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1573.LUT_INIT = 16'hfff4;
    SB_LUT4 i14329_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n32274));
    defparam i14329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1574 (.I0(n10_adj_6), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(GND_net), .O(n40142));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1574.LUT_INIT = 16'hfbfb;
    SB_LUT4 i4_4_lut_adj_1575 (.I0(\data_out_frame[21] [3]), .I1(n60268), 
            .I2(n60490), .I3(n6_adj_5640), .O(n54606));
    defparam i4_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1576 (.I0(n54689), .I1(n54606), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n61755));
    defparam i2_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 select_791_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1577 (.I0(\data_in_frame[9] [2]), .I1(n60208), 
            .I2(n60584), .I3(n28559), .O(n27843));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1578 (.I0(n61755), .I1(n54695), .I2(\data_out_frame[25] [7]), 
            .I3(GND_net), .O(n8_adj_5641));
    defparam i3_3_lut_adj_1578.LUT_INIT = 16'h6969;
    SB_LUT4 i13059_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n31004));   // verilog/coms.v(130[12] 305[6])
    defparam i13059_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_789_Select_208_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5641), .I3(\data_out_frame[23] [6]), 
            .O(n3_adj_5425));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_208_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1579 (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_5642), 
            .I2(reset), .I3(n86), .O(n30449));
    defparam i1_2_lut_3_lut_4_lut_adj_1579.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1580 (.I0(n30400), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[1]_c [2]), .O(n59316));
    defparam i1_4_lut_4_lut_4_lut_adj_1580.LUT_INIT = 16'hfe10;
    SB_LUT4 i14330_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n32275));
    defparam i14330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14331_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n32276));
    defparam i14331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14332_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n32277));
    defparam i14332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'ha088;
    SB_LUT4 i14333_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n32278));
    defparam i14333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1582 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [6]), 
            .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'ha088;
    SB_LUT4 i14334_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n32279));
    defparam i14334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1583 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [3]), 
            .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1583.LUT_INIT = 16'ha088;
    SB_LUT4 i14335_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n32280));
    defparam i14335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1584 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [2]), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1585 (.I0(n10_adj_5617), .I1(n152), .I2(GND_net), 
            .I3(GND_net), .O(n163));
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'heeee;
    SB_LUT4 i45045_2_lut_4_lut (.I0(control_mode[2]), .I1(n70677), .I2(PWMLimit[23]), 
            .I3(setpoint[23]), .O(n64302));
    defparam i45045_2_lut_4_lut.LUT_INIT = 16'heafe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1586 (.I0(n10_adj_6), .I1(n161), .I2(n3491), 
            .I3(n8_adj_5642), .O(n30366));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1586.LUT_INIT = 16'hffbf;
    SB_LUT4 i14336_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n32281));
    defparam i14336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14337_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n32282));
    defparam i14337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1587 (.I0(n10_adj_6), .I1(n161), .I2(n3491), 
            .I3(rx_data[7]), .O(n4_adj_5643));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1587.LUT_INIT = 16'h4000;
    SB_LUT4 select_789_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14338_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n32283));
    defparam i14338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [0]), 
            .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'ha088;
    SB_LUT4 i14339_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n32284));
    defparam i14339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n86), .I2(GND_net), .I3(GND_net), 
            .O(n80));
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i14340_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n32285));
    defparam i14340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14341_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n32286));
    defparam i14341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1589 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [3]), 
            .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1589.LUT_INIT = 16'ha088;
    SB_LUT4 i14342_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n32287));
    defparam i14342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1590 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [2]), 
            .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1590.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [1]), 
            .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1592 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n60026));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1592.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1593 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [0]), 
            .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1593.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14343_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n32288));
    defparam i14343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14344_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14]_c [3]), 
            .I3(deadband[19]), .O(n32289));
    defparam i14344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1594 (.I0(n10_adj_6), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n60017), .O(n30380));
    defparam i1_2_lut_3_lut_4_lut_adj_1594.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_4_lut (.I0(reset), .I1(n30400), .I2(\data_in_frame[1][1] ), 
            .I3(rx_data[1]), .O(n59308));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 select_789_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1595 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [4]), 
            .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1595.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51634_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[3]_c [5]), 
            .I2(n30416), .I3(GND_net), .O(n59298));   // verilog/coms.v(94[13:20])
    defparam i51634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51633_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[3]_c [4]), 
            .I2(n30416), .I3(GND_net), .O(n59294));   // verilog/coms.v(94[13:20])
    defparam i51633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14345_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][2] ), 
            .I3(deadband[18]), .O(n32290));
    defparam i14345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14346_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][1] ), 
            .I3(deadband[17]), .O(n32291));
    defparam i14346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18995_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21]_c [6]), 
            .I2(n24903), .I3(GND_net), .O(n32194));
    defparam i18995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19047_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21]_c [2]), 
            .I2(n24903), .I3(GND_net), .O(n32198));
    defparam i19047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14347_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14][0] ), 
            .I3(deadband[16]), .O(n32292));
    defparam i14347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71464_bdd_4_lut (.I0(n71464), .I1(n14_adj_5609), .I2(n7_adj_5644), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n71464_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [6]), 
            .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5571));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19048_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21][0] ), 
            .I2(n24903), .I3(GND_net), .O(n31464));
    defparam i19048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48734_2_lut (.I0(n71407), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67746));
    defparam i48734_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_789_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18821_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n24903), .I3(GND_net), .O(n32204));
    defparam i18821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18826_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1]_c [2]), 
            .I2(n24903), .I3(GND_net), .O(n32205));
    defparam i18826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18878_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n24877), .I3(GND_net), .O(n32219));
    defparam i18878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14348_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n32293));
    defparam i14348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18426_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n24877), .I3(GND_net), .O(n32223));
    defparam i18426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i167_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n167));
    defparam i167_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_789_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18431_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6][6] ), 
            .I2(n24877), .I3(GND_net), .O(n32224));
    defparam i18431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14349_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n32294));
    defparam i14349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14350_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n32295));
    defparam i14350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14351_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n32296));
    defparam i14351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_3_lut (.I0(LED_N_3408), .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2513 ), 
            .I3(GND_net), .O(n24877));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i14352_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n32297));
    defparam i14352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_3_lut_adj_1597 (.I0(Kp_23__N_612), .I1(reset), .I2(Kp_23__N_1748), 
            .I3(GND_net), .O(n24903));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut_adj_1597.LUT_INIT = 16'h2020;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52141 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71185), .I2(n67742), .I3(byte_transmit_counter_c[4]), 
            .O(n71458));
    defparam byte_transmit_counter_3__bdd_4_lut_52141.LUT_INIT = 16'he4aa;
    SB_LUT4 select_789_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14353_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n32298));
    defparam i14353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71458_bdd_4_lut (.I0(n71458), .I1(n71353), .I2(n7_adj_5645), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n71458_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1598 (.I0(n10), .I1(n60017), .I2(rx_data_ready), 
            .I3(\FRAME_MATCHER.rx_data_ready_prev ), .O(n30390));
    defparam i2_3_lut_4_lut_adj_1598.LUT_INIT = 16'hffef;
    SB_LUT4 select_789_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14354_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n32299));
    defparam i14354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_2_lut_adj_1599 (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n59757));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut_adj_1599.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_4_lut_adj_1600 (.I0(n55706), .I1(\data_out_frame[21] [5]), 
            .I2(n62106), .I3(n54653), .O(n54695));
    defparam i2_3_lut_4_lut_adj_1600.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1601 (.I0(\data_out_frame[21] [2]), .I1(n54982), 
            .I2(n60446), .I3(GND_net), .O(n54689));
    defparam i1_2_lut_3_lut_adj_1601.LUT_INIT = 16'h9696;
    SB_LUT4 i21_2_lut_4_lut (.I0(n1516), .I1(n60281), .I2(\data_out_frame[12] [4]), 
            .I3(\data_out_frame[14] [5]), .O(n29000));   // verilog/coms.v(100[12:26])
    defparam i21_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1602 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(n10_adj_5636), .I3(n60809), .O(n55719));
    defparam i5_3_lut_4_lut_adj_1602.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1603 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[10] [0]), 
            .I2(n28169), .I3(GND_net), .O(n60610));
    defparam i1_2_lut_3_lut_adj_1603.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1604 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(n60778), .I3(GND_net), .O(n60809));
    defparam i1_2_lut_3_lut_adj_1604.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1605 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[8][1] ), .I3(\data_out_frame[5] [3]), .O(n60066));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1605.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1606 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[9] [4]), .O(n6_adj_5624));
    defparam i1_2_lut_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1607 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n27774));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1608 (.I0(\data_out_frame[11][1] ), .I1(\data_out_frame[8][6] ), 
            .I2(n60156), .I3(GND_net), .O(n60714));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1608.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1609 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[9] [5]), .O(n60744));
    defparam i2_3_lut_4_lut_adj_1609.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1610 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[13] [2]), .I3(GND_net), .O(n6_adj_5620));
    defparam i1_2_lut_3_lut_adj_1610.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1611 (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[8][4] ), 
            .I2(\data_out_frame[8][5] ), .I3(GND_net), .O(n60108));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1611.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1612 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1));
    defparam i1_2_lut_adj_1612.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1613 (.I0(\data_out_frame[6] [6]), .I1(n60214), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n28918));
    defparam i1_2_lut_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1614 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[8][3] ), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[8][1] ), .O(n60062));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1614.LUT_INIT = 16'h6996;
    SB_LUT4 i14355_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n32300));
    defparam i14355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n60328));
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'h9696;
    SB_LUT4 i13540_3_lut (.I0(\data_in_frame[3]_c [1]), .I1(rx_data[1]), 
            .I2(n30416), .I3(GND_net), .O(n31485));   // verilog/coms.v(130[12] 305[6])
    defparam i13540_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i41707_3_lut (.I0(reset), .I1(n8_adj_5642), .I2(n60044), .I3(GND_net), 
            .O(n30416));
    defparam i41707_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5677_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1964), 
            .I2(n61882), .I3(n4452), .O(n23271));   // verilog/coms.v(148[4] 304[11])
    defparam i5677_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n23271), .I1(n1964), .I2(n24814), .I3(n4_adj_5638), 
            .O(n29161));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'hbbba;
    SB_LUT4 select_789_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2073));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14356_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n32301));
    defparam i14356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1617 (.I0(\data_out_frame[8][6] ), .I1(n60156), 
            .I2(n60788), .I3(\data_out_frame[12] [7]), .O(n61660));
    defparam i2_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 i45021_4_lut (.I0(n1964), .I1(n1967), .I2(n3303), .I3(n1970), 
            .O(n64276));   // verilog/coms.v(139[4] 141[7])
    defparam i45021_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i14357_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n32302));
    defparam i14357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_789_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1618 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1967), 
            .I2(n64276), .I3(n62294), .O(n58832));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1618.LUT_INIT = 16'hb3a0;
    SB_LUT4 i5682_4_lut (.I0(n1968), .I1(\FRAME_MATCHER.state[3] ), .I2(n1970), 
            .I3(n27595), .O(n23276));   // verilog/coms.v(148[4] 304[11])
    defparam i5682_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 select_789_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2062));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2061));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1619 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n6_adj_5646));   // verilog/coms.v(118[11:12])
    defparam i2_3_lut_adj_1619.LUT_INIT = 16'hecec;
    SB_LUT4 i18919_3_lut (.I0(n30414), .I1(rx_data[7]), .I2(\data_in_frame[2] [7]), 
            .I3(GND_net), .O(n32334));   // verilog/coms.v(94[13:20])
    defparam i18919_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13522_3_lut (.I0(\data_in_frame[2] [6]), .I1(rx_data[6]), .I2(n30414), 
            .I3(GND_net), .O(n31467));   // verilog/coms.v(130[12] 305[6])
    defparam i13522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23751_4_lut (.I0(n27491), .I1(\FRAME_MATCHER.i [31]), .I2(n6_adj_5646), 
            .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i23751_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 select_789_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1620 (.I0(\FRAME_MATCHER.i [4]), .I1(n27621), .I2(GND_net), 
            .I3(GND_net), .O(n27491));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1620.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n8_c));
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'hf7f7;
    SB_LUT4 i23754_4_lut (.I0(n27491), .I1(\FRAME_MATCHER.i [31]), .I2(n8_adj_5637), 
            .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i23754_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 select_789_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14358_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n32303));
    defparam i14358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14359_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n32304));
    defparam i14359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52136 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71191), .I2(n67730), .I3(byte_transmit_counter_c[4]), 
            .O(n71452));
    defparam byte_transmit_counter_3__bdd_4_lut_52136.LUT_INIT = 16'he4aa;
    SB_LUT4 n71452_bdd_4_lut (.I0(n71452), .I1(n71323), .I2(n7_adj_5647), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n71452_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52131 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71197), .I2(n67743), .I3(byte_transmit_counter_c[4]), 
            .O(n71446));
    defparam byte_transmit_counter_3__bdd_4_lut_52131.LUT_INIT = 16'he4aa;
    SB_LUT4 i22116_4_lut (.I0(n30362), .I1(n96), .I2(rx_data[7]), .I3(\data_in_frame[22] [7]), 
            .O(n39989));   // verilog/coms.v(94[13:20])
    defparam i22116_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22117_3_lut (.I0(n39989), .I1(\data_in_frame[22] [7]), .I2(reset), 
            .I3(GND_net), .O(n32349));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n24814));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(n10_adj_6), .I1(n144), .I2(GND_net), 
            .I3(GND_net), .O(n96));
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'h4444;
    SB_LUT4 i22146_4_lut (.I0(n30362), .I1(n96), .I2(rx_data[5]), .I3(\data_in_frame[22] [5]), 
            .O(n40019));   // verilog/coms.v(94[13:20])
    defparam i22146_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22147_3_lut (.I0(n40019), .I1(\data_in_frame[22] [5]), .I2(reset), 
            .I3(GND_net), .O(n32351));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(n27595), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n29711));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1623 (.I0(n4452), .I1(n29711), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n24814), .O(n61670));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1623.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_2_lut_adj_1624 (.I0(n10_adj_6), .I1(n152), .I2(GND_net), 
            .I3(GND_net), .O(n30362));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1624.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1625 (.I0(n8_c), .I1(\data_in_frame[21] [7]), 
            .I2(n30452), .I3(n4_adj_5643), .O(n59060));   // verilog/coms.v(94[13:20])
    defparam i13_4_lut_adj_1625.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n27610), .I1(n1970), .I2(n1968), .I3(n61670), 
            .O(n29158));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'hbaaa;
    SB_LUT4 i2_2_lut_adj_1627 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5648));
    defparam i2_2_lut_adj_1627.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1628 (.I0(n39975), .I1(\data_in_frame[21]_c [6]), 
            .I2(n30452), .I3(n4_adj_5649), .O(n59058));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1628.LUT_INIT = 16'hc5c0;
    SB_LUT4 select_789_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i6_4_lut_adj_1629 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5650));
    defparam i6_4_lut_adj_1629.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1630 (.I0(\data_in[3] [6]), .I1(n14_adj_5650), 
            .I2(n10_adj_5648), .I3(\data_in[2] [1]), .O(n27634));
    defparam i7_4_lut_adj_1630.LUT_INIT = 16'hfffd;
    SB_LUT4 i14360_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n32305));
    defparam i14360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_3_lut_adj_1631 (.I0(rx_data[2]), .I1(\data_in_frame[21]_c [2]), 
            .I2(n30452), .I3(GND_net), .O(n59046));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1631.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_adj_1632 (.I0(rx_data[1]), .I1(\data_in_frame[21][1] ), 
            .I2(n30452), .I3(GND_net), .O(n59050));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1632.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1633 (.I0(n27634), .I1(\data_in[3] [7]), .I2(n27521), 
            .I3(\data_in[1] [6]), .O(n20_adj_5651));
    defparam i8_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i14361_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n32306));
    defparam i14361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[25] [7]), 
            .I2(n25812), .I3(GND_net), .O(n8_adj_5596));
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1635 (.I0(\data_in[1] [3]), .I1(\data_in[2] [6]), 
            .I2(\data_in[0] [5]), .I3(\data_in[1] [2]), .O(n19_adj_5652));
    defparam i7_4_lut_adj_1635.LUT_INIT = 16'hdfff;
    SB_LUT4 n71446_bdd_4_lut (.I0(n71446), .I1(n71335), .I2(n7_adj_5653), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[2]));
    defparam n71446_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i45222_4_lut (.I0(\data_in[3] [2]), .I1(\data_in[2] [5]), .I2(\data_in[0] [1]), 
            .I3(\data_in[2] [0]), .O(n64483));
    defparam i45222_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1636 (.I0(n64483), .I1(n19_adj_5652), .I2(n20_adj_5651), 
            .I3(GND_net), .O(n1964));
    defparam i11_3_lut_adj_1636.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1637 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n62354), .I3(GND_net), .O(n6_adj_5594));
    defparam i1_2_lut_3_lut_adj_1637.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[13] [6]), .I1(n54789), .I2(n45_adj_5588), 
            .I3(GND_net), .O(n7_adj_5592));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14362_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n32307));
    defparam i14362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_3_lut_4_lut_adj_1638 (.I0(\data_out_frame[16] [1]), .I1(n55645), 
            .I2(\data_out_frame[18] [2]), .I3(n55303), .O(n8_adj_5593));
    defparam i3_3_lut_4_lut_adj_1638.LUT_INIT = 16'h9669;
    SB_LUT4 select_789_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i18879_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [1]), 
            .I3(\data_in_frame[19]_c [1]), .O(n4947[1]));
    defparam i18879_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i7_4_lut_adj_1639 (.I0(\data_in[2] [4]), .I1(\data_in[1] [5]), 
            .I2(n27634), .I3(n27684), .O(n18_adj_5654));
    defparam i7_4_lut_adj_1639.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1640 (.I0(\data_in[0] [6]), .I1(n18_adj_5654), 
            .I2(\data_in[3] [0]), .I3(n27658), .O(n20_adj_5655));
    defparam i9_4_lut_adj_1640.LUT_INIT = 16'hfffd;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52126 (.I0(byte_transmit_counter_c[3]), 
            .I1(n71203), .I2(n67755), .I3(byte_transmit_counter_c[4]), 
            .O(n71440));
    defparam byte_transmit_counter_3__bdd_4_lut_52126.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1641 (.I0(\data_out_frame[4] [6]), .I1(n60214), 
            .I2(\data_out_frame[7] [0]), .I3(n28918), .O(n60729));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1641.LUT_INIT = 16'h6996;
    SB_LUT4 n71440_bdd_4_lut (.I0(n71440), .I1(n71305), .I2(n7_adj_5656), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n71440_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_2_lut (.I0(\data_in[2] [2]), .I1(\data_in[1] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5657));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1642 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [0]), 
            .I2(n55105), .I3(GND_net), .O(n6_adj_5582));
    defparam i1_2_lut_3_lut_adj_1642.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1643 (.I0(n27770), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(\data_out_frame[10] [6]), .O(n60625));
    defparam i2_3_lut_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52186 (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5607), .I2(n5_adj_5606), .I3(byte_transmit_counter[2]), 
            .O(n71434));
    defparam byte_transmit_counter_1__bdd_4_lut_52186.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1089_i3_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][2] ), .I3(\data_in_frame[19][2] ), .O(n4947[2]));
    defparam mux_1089_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i5_3_lut_4_lut_adj_1644 (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[8][7] ), 
            .I2(n10_adj_5572), .I3(\data_out_frame[6] [6]), .O(n27799));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1645 (.I0(n54936), .I1(n60322), .I2(n60695), 
            .I3(\data_out_frame[18] [4]), .O(n60449));
    defparam i1_2_lut_4_lut_adj_1645.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1646 (.I0(\data_in_frame[19]_c [6]), .I1(n30366), 
            .I2(n30449), .I3(rx_data[6]), .O(n59118));
    defparam i12_4_lut_adj_1646.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14_4_lut_adj_1647 (.I0(\data_in_frame[19]_c [5]), .I1(n7_adj_5467), 
            .I2(n30449), .I3(n4_adj_5658), .O(n59052));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1647.LUT_INIT = 16'h3a0a;
    SB_LUT4 i10_4_lut_adj_1648 (.I0(n15_adj_5657), .I1(n20_adj_5655), .I2(\data_in[0] [3]), 
            .I3(\data_in[1] [4]), .O(n1967));
    defparam i10_4_lut_adj_1648.LUT_INIT = 16'hfeff;
    SB_LUT4 i22300_4_lut (.I0(n30366), .I1(n53), .I2(rx_data[4]), .I3(\data_in_frame[19]_c [4]), 
            .O(n40172));   // verilog/coms.v(94[13:20])
    defparam i22300_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22301_3_lut (.I0(n40172), .I1(\data_in_frame[19]_c [4]), .I2(reset), 
            .I3(GND_net), .O(n32435));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_adj_1649 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [7]), 
            .I2(n60145), .I3(GND_net), .O(n7_adj_5568));
    defparam i2_2_lut_3_lut_adj_1649.LUT_INIT = 16'h9696;
    SB_LUT4 i22285_4_lut (.I0(n30366), .I1(n53), .I2(rx_data[3]), .I3(\data_in_frame[19]_c [3]), 
            .O(n40157));   // verilog/coms.v(94[13:20])
    defparam i22285_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22286_3_lut (.I0(n40157), .I1(\data_in_frame[19]_c [3]), .I2(reset), 
            .I3(GND_net), .O(n32437));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1650 (.I0(\data_in_frame[19]_c [1]), .I1(n8_adj_5642), 
            .I2(n30449), .I3(rx_data[1]), .O(n59106));   // verilog/coms.v(94[13:20])
    defparam i13_4_lut_adj_1650.LUT_INIT = 16'h3a0a;
    SB_LUT4 i2_2_lut_4_lut_adj_1651 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(\FRAME_MATCHER.i_31__N_2512 ), 
            .O(n6_adj_5565));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i13069_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n31014));   // verilog/coms.v(130[12] 305[6])
    defparam i13069_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mux_1089_i4_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][3] ), .I3(\data_in_frame[19]_c [3]), .O(n4947[3]));
    defparam mux_1089_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i4_4_lut_adj_1652 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5659));
    defparam i4_4_lut_adj_1652.LUT_INIT = 16'hfdff;
    SB_LUT4 i11_3_lut_adj_1653 (.I0(\data_in_frame[18]_c [7]), .I1(rx_data[7]), 
            .I2(n30447), .I3(GND_net), .O(n59064));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1653.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_adj_1654 (.I0(\data_in[3] [4]), .I1(n10_adj_5659), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n27658));
    defparam i5_3_lut_adj_1654.LUT_INIT = 16'hdfdf;
    SB_LUT4 i3_4_lut_adj_1655 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n3491), .I3(n161), .O(n86));
    defparam i3_4_lut_adj_1655.LUT_INIT = 16'h2000;
    SB_LUT4 select_789_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i5_3_lut_4_lut_adj_1656 (.I0(\data_in_frame[6][4] ), .I1(\data_in_frame[0] [3]), 
            .I2(n60122), .I3(n60613), .O(n14_adj_5553));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1657 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5660));
    defparam i5_3_lut_adj_1657.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1658 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(n27900), .I3(n64147), .O(n64151));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i14017_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n62670), .I3(GND_net), .O(n31962));   // verilog/coms.v(130[12] 305[6])
    defparam i14017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14012_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n62670), .I3(GND_net), .O(n31957));   // verilog/coms.v(130[12] 305[6])
    defparam i14012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1089_i5_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3]_c [4]), .I3(\data_in_frame[19]_c [4]), 
            .O(n4947[4]));
    defparam mux_1089_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i6_4_lut_adj_1659 (.I0(\data_in[0] [6]), .I1(n27658), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5661));
    defparam i6_4_lut_adj_1659.LUT_INIT = 16'hfeff;
    SB_LUT4 i17074_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [5]), 
            .I3(\data_in_frame[19]_c [5]), .O(n4947[5]));
    defparam i17074_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i8_4_lut_adj_1660 (.I0(n15_adj_5661), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5660), .I3(\data_in[0] [3]), .O(n27521));
    defparam i8_4_lut_adj_1660.LUT_INIT = 16'hfbff;
    SB_LUT4 n71434_bdd_4_lut (.I0(n71434), .I1(n67615), .I2(n1_adj_5605), 
            .I3(byte_transmit_counter[2]), .O(n71437));
    defparam n71434_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1089_i20_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1]_c [3]), .I3(\data_in_frame[17][3] ), .O(n4947[19]));
    defparam mux_1089_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1089_i21_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17][4] ), .O(n4947[20]));
    defparam mux_1089_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52025 (.I0(byte_transmit_counter[1]), 
            .I1(n64899), .I2(n64900), .I3(byte_transmit_counter[2]), .O(n71302));
    defparam byte_transmit_counter_1__bdd_4_lut_52025.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1089_i22_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17][5] ), .O(n4947[21]));
    defparam mux_1089_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut_4_lut_adj_1661 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6][3] ), 
            .I2(\data_in_frame[6][2] ), .I3(\data_in_frame[6][1] ), .O(n60747));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5566));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1662 (.I0(\data_in_frame[0] [3]), .I1(n60122), 
            .I2(\data_in_frame[2][3] ), .I3(n60515), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1089_i23_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17][6] ), .O(n4947[22]));
    defparam mux_1089_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut_4_lut_adj_1663 (.I0(n40142), .I1(n3491), .I2(n8_adj_5637), 
            .I3(reset), .O(n62228));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1663.LUT_INIT = 16'hfffb;
    SB_LUT4 select_791_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_c));   // verilog/coms.v(148[4] 304[11])
    defparam select_791_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i6_4_lut_adj_1664 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5662));
    defparam i6_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1665 (.I0(n40142), .I1(n3491), .I2(reset), 
            .I3(n8_c), .O(n30452));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1665.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1666 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2][1] ), .I3(GND_net), .O(n60142));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1666.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1667 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5663));
    defparam i7_4_lut_adj_1667.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1668 (.I0(n40142), .I1(n3491), .I2(n7_adj_5467), 
            .I3(\FRAME_MATCHER.i[0] ), .O(n30368));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1668.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1669 (.I0(n40142), .I1(n3491), .I2(rx_data[5]), 
            .I3(\FRAME_MATCHER.i[0] ), .O(n4_adj_5658));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1669.LUT_INIT = 16'h4000;
    SB_LUT4 mux_1089_i24_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17][7] ), .O(n4947[23]));
    defparam mux_1089_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1670 (.I0(n40142), .I1(n3491), .I2(rx_data[6]), 
            .I3(\FRAME_MATCHER.i[0] ), .O(n4_adj_5649));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1670.LUT_INIT = 16'h4000;
    SB_LUT4 mux_1089_i1_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][0] ), .I3(\data_in_frame[19] [0]), .O(n4947[0]));
    defparam mux_1089_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_789_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5291));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1089_i8_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19][7] ), .O(n4947[7]));
    defparam mux_1089_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_3_lut_4_lut_adj_1671 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n60026), .I3(LED_c), .O(n29481));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1671.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1672 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3491));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1672.LUT_INIT = 16'hfefe;
    SB_LUT4 n71302_bdd_4_lut (.I0(n71302), .I1(n64591), .I2(n64590), .I3(byte_transmit_counter[2]), 
            .O(n71305));
    defparam n71302_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1089_i9_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][0] ), .I3(\data_in_frame[18][0] ), .O(n4947[8]));
    defparam mux_1089_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1089_i10_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][1] ), .I3(\data_in_frame[18][1] ), .O(n4947[9]));
    defparam mux_1089_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i48914_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67691));   // verilog/coms.v(158[12:15])
    defparam i48914_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48911_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67690));   // verilog/coms.v(158[12:15])
    defparam i48911_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_adj_1673 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n60545), .I3(n27996), .O(Kp_23__N_767));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i48892_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67689));   // verilog/coms.v(158[12:15])
    defparam i48892_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48876_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67683));   // verilog/coms.v(158[12:15])
    defparam i48876_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_1674 (.I0(n17_adj_5663), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5662), .I3(\data_in[2] [6]), .O(n27684));
    defparam i9_4_lut_adj_1674.LUT_INIT = 16'hfbff;
    SB_LUT4 i48856_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67682));   // verilog/coms.v(158[12:15])
    defparam i48856_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48842_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67679));   // verilog/coms.v(158[12:15])
    defparam i48842_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48841_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67678));   // verilog/coms.v(158[12:15])
    defparam i48841_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1675 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n27521), .O(n16_adj_5664));
    defparam i6_4_lut_adj_1675.LUT_INIT = 16'hffef;
    SB_LUT4 i48765_2_lut (.I0(n71413), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67745));
    defparam i48765_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50367_3_lut (.I0(n71497), .I1(n71299), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n69637));
    defparam i50367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49454_2_lut (.I0(n71419), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67758));
    defparam i49454_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1089_i11_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][2] ), .I3(\data_in_frame[18][2] ), .O(n4947[10]));
    defparam mux_1089_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1089_i12_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][3] ), .I3(\data_in_frame[18][3] ), .O(n4947[11]));
    defparam mux_1089_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i50400_3_lut (.I0(n71479), .I1(n71371), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n69670));
    defparam i50400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48833_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67677));   // verilog/coms.v(158[12:15])
    defparam i48833_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48838_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67676));   // verilog/coms.v(158[12:15])
    defparam i48838_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1089_i13_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][4] ), .I3(\data_in_frame[18][4] ), .O(n4947[12]));
    defparam mux_1089_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i48830_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67673));   // verilog/coms.v(158[12:15])
    defparam i48830_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48828_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67672));   // verilog/coms.v(158[12:15])
    defparam i48828_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1089_i14_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][5] ), .I3(\data_in_frame[18] [5]), .O(n4947[13]));
    defparam mux_1089_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_789_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5564));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48651_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67671));   // verilog/coms.v(158[12:15])
    defparam i48651_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1676 (.I0(n27684), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5665));
    defparam i7_4_lut_adj_1676.LUT_INIT = 16'hbfff;
    SB_LUT4 i49465_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67659));   // verilog/coms.v(158[12:15])
    defparam i49465_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1089_i15_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n4947[14]));
    defparam mux_1089_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i48808_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67651));   // verilog/coms.v(158[12:15])
    defparam i48808_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48807_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67650));   // verilog/coms.v(158[12:15])
    defparam i48807_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48806_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67649));   // verilog/coms.v(158[12:15])
    defparam i48806_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48805_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67648));   // verilog/coms.v(158[12:15])
    defparam i48805_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48804_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67647));   // verilog/coms.v(158[12:15])
    defparam i48804_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48906_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67646));   // verilog/coms.v(158[12:15])
    defparam i48906_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1677 (.I0(n64302), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(n15_adj_5666), .O(n16_adj_5667));
    defparam i7_4_lut_adj_1677.LUT_INIT = 16'h0100;
    SB_LUT4 i8_4_lut_adj_1678 (.I0(control_update), .I1(n16_adj_5667), .I2(n41374), 
            .I3(control_mode[3]), .O(n27538));
    defparam i8_4_lut_adj_1678.LUT_INIT = 16'h0008;
    SB_LUT4 i48703_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67602));   // verilog/coms.v(158[12:15])
    defparam i48703_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48711_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67601));   // verilog/coms.v(158[12:15])
    defparam i48711_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48693_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67596));   // verilog/coms.v(158[12:15])
    defparam i48693_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_1679 (.I0(n17_adj_5665), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5664), .I3(\data_in[3] [3]), .O(n1970));
    defparam i9_4_lut_adj_1679.LUT_INIT = 16'hfbff;
    SB_LUT4 i48694_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67595));   // verilog/coms.v(158[12:15])
    defparam i48694_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48675_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67592));   // verilog/coms.v(158[12:15])
    defparam i48675_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49487_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67591));   // verilog/coms.v(158[12:15])
    defparam i49487_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52117 (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5604), .I2(n5_adj_5603), .I3(byte_transmit_counter[2]), 
            .O(n71428));
    defparam byte_transmit_counter_1__bdd_4_lut_52117.LUT_INIT = 16'he4aa;
    SB_LUT4 i48770_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67588));   // verilog/coms.v(158[12:15])
    defparam i48770_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48632_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67581));   // verilog/coms.v(158[12:15])
    defparam i48632_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1680 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n60011));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1680.LUT_INIT = 16'heeee;
    SB_LUT4 i48631_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67580));   // verilog/coms.v(158[12:15])
    defparam i48631_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48860_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67579));   // verilog/coms.v(158[12:15])
    defparam i48860_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48626_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67577));   // verilog/coms.v(158[12:15])
    defparam i48626_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i18920_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[18]_c [7]), .O(n4947[15]));
    defparam i18920_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1089_i17_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][0] ), .I3(\data_in_frame[17][0] ), .O(n4947[16]));
    defparam mux_1089_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1681 (.I0(n61729), .I1(\data_in_frame[16] [6]), 
            .I2(n54742), .I3(\data_in_frame[17][0] ), .O(n60759));
    defparam i1_2_lut_3_lut_4_lut_adj_1681.LUT_INIT = 16'h9669;
    SB_LUT4 i19387_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[1][1] ), 
            .I3(\data_in_frame[17] [1]), .O(n4947[17]));
    defparam i19387_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52020 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71296));
    defparam byte_transmit_counter_0__bdd_4_lut_52020.LUT_INIT = 16'he4aa;
    SB_LUT4 i19388_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[1]_c [2]), 
            .I3(\data_in_frame[17] [2]), .O(n4947[18]));
    defparam i19388_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i48772_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67576));   // verilog/coms.v(158[12:15])
    defparam i48772_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12417_1_lut (.I0(n3491), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30361));   // verilog/coms.v(148[4] 304[11])
    defparam i12417_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i366_2_lut (.I0(n1967), .I1(n1964), .I2(GND_net), .I3(GND_net), 
            .O(n1968));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17066_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[19]_c [6]), .O(n4947[6]));
    defparam i17066_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_3_lut_4_lut_adj_1682 (.I0(\data_in_frame[6][6] ), .I1(\data_in_frame[6][5] ), 
            .I2(\data_in_frame[4] [5]), .I3(\data_in_frame[6][4] ), .O(n64047));   // verilog/coms.v(88[17:28])
    defparam i1_3_lut_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 i48875_2_lut (.I0(\data_out_frame[9] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67644));
    defparam i48875_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48907_2_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n67645));
    defparam i48907_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1683 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5668));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1683.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5669));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_4_lut_adj_1685 (.I0(\data_in_frame[6][0] ), .I1(\data_in_frame[6] [7]), 
            .I2(n28006), .I3(\data_in_frame[6][1] ), .O(n60287));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1685.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1686 (.I0(\data_in_frame[6][1] ), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [7]), .O(n60548));   // verilog/coms.v(18[27:29])
    defparam i2_3_lut_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_LUT4 n71296_bdd_4_lut (.I0(n71296), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71299));
    defparam n71296_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i24050_4_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5669), .I3(n4_adj_5668), .O(n41899));
    defparam i24050_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1_2_lut_4_lut_adj_1687 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [5]), 
            .I2(n61729), .I3(n60190), .O(n6_adj_5507));
    defparam i1_2_lut_4_lut_adj_1687.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1688 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(n60122), .I3(n28463), .O(n28432));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1688.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6][6] ), 
            .I2(\data_in_frame[6][5] ), .I3(GND_net), .O(n60296));   // verilog/coms.v(18[27:29])
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 n71428_bdd_4_lut (.I0(n71428), .I1(n67617), .I2(n67616), .I3(byte_transmit_counter[2]), 
            .O(n71431));
    defparam n71428_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n1968), .I1(n60011), .I2(n1970), .I3(\FRAME_MATCHER.i_31__N_2507 ), 
            .O(n5_adj_5670));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'heccc;
    SB_LUT4 i3_4_lut_adj_1691 (.I0(n5_adj_5670), .I1(n62599), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n71700));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1691.LUT_INIT = 16'hefee;
    SB_LUT4 i1_2_lut_3_lut_adj_1692 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n60562));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1693 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10] [7]), 
            .I2(n60524), .I3(n28041), .O(n61746));
    defparam i2_3_lut_4_lut_adj_1693.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1694 (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(n54662), .I3(\data_in_frame[11] [0]), .O(n60524));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1695 (.I0(\data_in_frame[6][5] ), .I1(\data_in_frame[6][4] ), 
            .I2(Kp_23__N_875), .I3(n36324), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1696 (.I0(n27956), .I1(\data_in_frame[9] [0]), 
            .I2(n27211), .I3(Kp_23__N_1080), .O(n54872));
    defparam i1_3_lut_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 i51785_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n41899), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i51785_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_4_lut_adj_1697 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n41899), .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n27595));
    defparam i1_3_lut_4_lut_adj_1697.LUT_INIT = 16'hef00;
    SB_LUT4 i2_3_lut_4_lut_adj_1698 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(\FRAME_MATCHER.i_31__N_2511 ), .I3(n41899), .O(n62599));
    defparam i2_3_lut_4_lut_adj_1698.LUT_INIT = 16'h1000;
    SB_LUT4 i13855_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n31800));
    defparam i13855_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14473_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[1][0] ), .O(n32418));
    defparam i14473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13858_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n31803));
    defparam i13858_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13861_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n31806));
    defparam i13861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13864_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n31809));
    defparam i13864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1699 (.I0(n60208), .I1(n60584), .I2(n28559), 
            .I3(GND_net), .O(n60309));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1699.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i12_3_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\data_out_frame[15] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12_adj_5544));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i11_3_lut (.I0(\data_out_frame[12] [0]), 
            .I1(\data_out_frame[13] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13867_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n31812));
    defparam i13867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14482_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n32427));
    defparam i14482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13492_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n31437));
    defparam i13492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1700 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n54662), .I3(n28055), .O(n55574));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1700.LUT_INIT = 16'h9669;
    SB_LUT4 i13488_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n31433));
    defparam i13488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13870_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n31815));
    defparam i13870_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13481_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n31426));
    defparam i13481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13484_3_lut_4_lut (.I0(n30400), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n31429));
    defparam i13484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[12] [5]), .I1(n28583), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[10] [6]), .O(n6_adj_5481));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5542));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13873_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n31818));
    defparam i13873_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1701 (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_5642), 
            .I2(n86), .I3(GND_net), .O(n53));
    defparam i1_2_lut_3_lut_adj_1701.LUT_INIT = 16'h1010;
    SB_LUT4 i13876_3_lut_4_lut (.I0(n8_adj_5642), .I1(n60036), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n31821));
    defparam i13876_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i45332_3_lut (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64602));
    defparam i45332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45333_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11][3] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64603));
    defparam i45333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1702 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_6));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_adj_1702.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12114_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3491), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n30058));   // verilog/coms.v(158[12:15])
    defparam i12114_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 select_1747_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_1747_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45627_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64897));
    defparam i45627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45626_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64896));
    defparam i45626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1703 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n27294), .I3(GND_net), .O(n54602));
    defparam i1_2_lut_3_lut_adj_1703.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1704 (.I0(\data_in_frame[5][6] ), .I1(n28009), 
            .I2(n10_adj_5516), .I3(n27971), .O(n28583));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 i14117_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n32062));
    defparam i14117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1705 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [2]), .I3(GND_net), .O(n60559));   // verilog/coms.v(18[27:29])
    defparam i1_2_lut_3_lut_adj_1705.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14114_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n32059));
    defparam i14114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(\data_in_frame[20] [5]), 
            .I3(rx_data[5]), .O(n59214));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i14106_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n32051));
    defparam i14106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1706 (.I0(n28572), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[12] [3]), .I3(\data_in_frame[12] [2]), .O(n60518));
    defparam i2_3_lut_4_lut_adj_1706.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1707 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n26041), .I3(n26045), .O(n28572));
    defparam i1_2_lut_4_lut_adj_1707.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1708 (.I0(n28930), .I1(n55163), .I2(\data_in_frame[9] [7]), 
            .I3(n27992), .O(n55710));
    defparam i2_3_lut_4_lut_adj_1708.LUT_INIT = 16'h6996;
    SB_LUT4 i14103_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n32048));
    defparam i14103_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n59322));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14096_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n32041));
    defparam i14096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14093_3_lut_4_lut (.I0(n30380), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n32038));
    defparam i14093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1709 (.I0(n28134), .I1(n28583), .I2(n54624), 
            .I3(GND_net), .O(n60769));
    defparam i1_2_lut_3_lut_adj_1709.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5527));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1710 (.I0(\data_in_frame[16] [5]), .I1(n61729), 
            .I2(n60190), .I3(GND_net), .O(n60763));
    defparam i1_2_lut_3_lut_adj_1710.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1711 (.I0(n28930), .I1(n60467), .I2(n27992), 
            .I3(\data_in_frame[10] [1]), .O(n55712));
    defparam i1_2_lut_4_lut_adj_1711.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n60726));
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1713 (.I0(\data_in_frame[18]_c [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n60275), .I3(GND_net), .O(n27264));
    defparam i1_2_lut_3_lut_adj_1713.LUT_INIT = 16'h9696;
    SB_LUT4 select_789_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1714 (.I0(\data_in_frame[18][2] ), .I1(\data_in_frame[18][4] ), 
            .I2(n55556), .I3(GND_net), .O(n60458));
    defparam i1_2_lut_3_lut_adj_1714.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1715 (.I0(n27251), .I1(n60619), .I2(\data_in_frame[14][0] ), 
            .I3(n28074), .O(n6_adj_5492));
    defparam i1_2_lut_4_lut_adj_1715.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1716 (.I0(\data_in_frame[18][3] ), .I1(n60368), 
            .I2(n10_adj_5489), .I3(Kp_23__N_1271), .O(n55778));
    defparam i1_2_lut_4_lut_adj_1716.LUT_INIT = 16'h9669;
    SB_LUT4 i14153_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n32098));
    defparam i14153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1717 (.I0(n55186), .I1(\data_in_frame[9] [4]), 
            .I2(n28386), .I3(\data_in_frame[9] [3]), .O(n60622));
    defparam i2_3_lut_4_lut_adj_1717.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[16] [0]), 
            .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_adj_1719 (.I0(n62393), .I1(n28247), .I2(n62554), 
            .I3(n60461), .O(n60257));
    defparam i1_2_lut_4_lut_adj_1719.LUT_INIT = 16'h6996;
    SB_LUT4 i14452_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n32397));
    defparam i14452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14455_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n32400));
    defparam i14455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14458_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n32403));
    defparam i14458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14461_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n32406));
    defparam i14461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14464_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n32409));
    defparam i14464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_2_lut (.I0(PWMLimit[22]), .I1(setpoint[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14467_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n32412));
    defparam i14467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14470_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60032), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n32415));
    defparam i14470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_2_lut_adj_1720 (.I0(PWMLimit[15]), .I1(setpoint[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i13_2_lut_adj_1720.LUT_INIT = 16'h6666;
    SB_LUT4 i17934_3_lut (.I0(n28), .I1(PWMLimit[14]), .I2(setpoint[14]), 
            .I3(GND_net), .O(n30));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i17934_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_adj_1721 (.I0(control_mode[1]), .I1(control_mode[0]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5666));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1721.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1722 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(n58710), .O(n60461));
    defparam i1_2_lut_4_lut_adj_1722.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1723 (.I0(\data_in_frame[17] [1]), .I1(n54563), 
            .I2(\data_in_frame[19]_c [3]), .I3(n62306), .O(n61855));
    defparam i2_3_lut_4_lut_adj_1723.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1724 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1964), .I3(n1967), .O(n27610));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1724.LUT_INIT = 16'h4000;
    SB_LUT4 i51632_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(\data_in_frame[23] [7]), 
            .I3(rx_data[7]), .O(n59230));
    defparam i51632_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1725 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[13] [7]), 
            .I2(n60698), .I3(GND_net), .O(n60202));
    defparam i1_2_lut_3_lut_adj_1725.LUT_INIT = 16'h9696;
    SB_LUT4 i14204_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n32149));
    defparam i14204_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14201_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n32146));
    defparam i14201_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14188_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n32133));
    defparam i14188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14195_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n32140));
    defparam i14195_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1726 (.I0(n28074), .I1(n60319), .I2(n60772), 
            .I3(GND_net), .O(n60765));
    defparam i1_2_lut_3_lut_adj_1726.LUT_INIT = 16'h9696;
    SB_LUT4 i14185_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n32130));
    defparam i14185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14198_3_lut_4_lut (.I0(n30370), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n32143));
    defparam i14198_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1727 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5674));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1727.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1728 (.I0(n1964), .I1(n4452), .I2(n1967), 
            .I3(n1970), .O(n61882));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1728.LUT_INIT = 16'h2000;
    SB_LUT4 i1_3_lut_4_lut_adj_1729 (.I0(n28908), .I1(n27873), .I2(n60817), 
            .I3(n55599), .O(n62783));
    defparam i1_3_lut_4_lut_adj_1729.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1964), .I1(n4452), .I2(n4_adj_5638), 
            .I3(\FRAME_MATCHER.i_31__N_2514 ), .O(n62294));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i2_3_lut_4_lut_adj_1730 (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_5467), 
            .I2(n80), .I3(\FRAME_MATCHER.i [5]), .O(n30447));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_4_lut_adj_1730.LUT_INIT = 16'h0010;
    SB_LUT4 i13955_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n31900));
    defparam i13955_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13958_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n31903));
    defparam i13958_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13964_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n31909));
    defparam i13964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1731 (.I0(\data_in_frame[19] [0]), .I1(n28753), 
            .I2(n64089), .I3(\data_in_frame[18][2] ), .O(n60601));
    defparam i1_2_lut_4_lut_adj_1731.LUT_INIT = 16'h6996;
    SB_LUT4 i13967_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n31912));
    defparam i13967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13970_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n31915));
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13973_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n31918));
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13976_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n31921));
    defparam i13976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13979_3_lut_4_lut (.I0(n167), .I1(n60036), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n31924));
    defparam i13979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_789_Select_212_i3_3_lut_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(n62047), .I2(\FRAME_MATCHER.state[3] ), .I3(n60487), .O(n3_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_212_i3_3_lut_4_lut.LUT_INIT = 16'h6090;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1732 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(Kp_23__N_1271), .I3(n27294), .O(n60772));
    defparam i1_2_lut_3_lut_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1733 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60515));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1733.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1734 (.I0(n60368), .I1(n10_adj_5489), .I2(\data_in_frame[13] [7]), 
            .I3(\data_in_frame[13] [6]), .O(n61984));
    defparam i5_3_lut_4_lut_adj_1734.LUT_INIT = 16'h6996;
    SB_LUT4 i13764_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n31709));
    defparam i13764_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13767_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n31712));
    defparam i13767_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12470_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_5467), 
            .I2(n60044), .I3(reset), .O(n30414));   // verilog/coms.v(157[7:23])
    defparam i12470_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13770_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n31715));
    defparam i13770_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13773_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n31718));
    defparam i13773_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13776_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n31721));
    defparam i13776_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13779_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n31724));
    defparam i13779_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13782_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n31727));
    defparam i13782_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13785_3_lut_4_lut (.I0(n8_adj_5637), .I1(n60036), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n31730));
    defparam i13785_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13582_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n31527));
    defparam i13582_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13579_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n31524));
    defparam i13579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13576_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n31521));
    defparam i13576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13573_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n31518));
    defparam i13573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1735 (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_5674), 
            .I2(n60002), .I3(n40142), .O(n62670));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_4_lut_adj_1735.LUT_INIT = 16'hfffd;
    SB_LUT4 i13567_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n31512));
    defparam i13567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut_adj_1736 (.I0(n30390), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n59304));
    defparam i11_4_lut_4_lut_adj_1736.LUT_INIT = 16'hfe10;
    SB_LUT4 i13561_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n31506));
    defparam i13561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13570_3_lut_4_lut (.I0(n30390), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n31515));
    defparam i13570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52151 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n71416));
    defparam byte_transmit_counter_0__bdd_4_lut_52151.LUT_INIT = 16'he4aa;
    SB_LUT4 n71416_bdd_4_lut (.I0(n71416), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71419));
    defparam n71416_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52102 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71410));
    defparam byte_transmit_counter_0__bdd_4_lut_52102.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(n28055), .I1(n60319), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n60662));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h9696;
    SB_LUT4 equal_302_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n8_adj_5642));   // verilog/coms.v(157[7:23])
    defparam equal_302_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1737 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[18][3] ), 
            .I2(n64089), .I3(\data_in_frame[18][2] ), .O(n60735));
    defparam i1_3_lut_4_lut_adj_1737.LUT_INIT = 16'h6996;
    SB_LUT4 n71410_bdd_4_lut (.I0(n71410), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71413));
    defparam n71410_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(n27971), .I3(\data_in_frame[8] [0]), .O(n20_adj_5496));   // verilog/coms.v(81[16:27])
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1738 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n3491), .O(n60017));
    defparam i1_2_lut_3_lut_4_lut_adj_1738.LUT_INIT = 16'hfbff;
    SB_LUT4 i13631_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n30423), 
            .I3(GND_net), .O(n31576));   // verilog/coms.v(130[12] 305[6])
    defparam i13631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1739 (.I0(\data_out_frame[16] [4]), .I1(n28303), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n60616));
    defparam i1_2_lut_3_lut_adj_1739.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1740 (.I0(\data_out_frame[16] [4]), .I1(n28303), 
            .I2(n60689), .I3(GND_net), .O(n6_adj_5640));
    defparam i1_2_lut_3_lut_adj_1740.LUT_INIT = 16'h9696;
    SB_LUT4 i45446_3_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64716));
    defparam i45446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45447_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11][7] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64717));
    defparam i45447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45378_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64648));
    defparam i45378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[16] [7]), 
            .I2(n60478), .I3(n60797), .O(n11_adj_5579));   // verilog/coms.v(100[12:26])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i45377_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64647));
    defparam i45377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1741 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [1]), .I3(n60355), .O(n60689));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1741.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1742 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n60036), .O(n60038));
    defparam i1_2_lut_3_lut_4_lut_adj_1742.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1743 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [3]), .I3(n60797), .O(n6_adj_5608));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1743.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64871), .I3(n64869), .O(n7_adj_5656));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64664), .I3(n64662), .O(n7_adj_5653));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64706), .I3(n64704), .O(n7_adj_5647));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_2_lut_3_lut_adj_1744 (.I0(n61872), .I1(n60635), .I2(\data_out_frame[25] [0]), 
            .I3(GND_net), .O(n6_adj_5423));
    defparam i2_2_lut_3_lut_adj_1744.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64682), .I3(n64680), .O(n7_adj_5645));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64880), .I3(n64878), .O(n7_adj_5581));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64679), .I3(n64677), .O(n7_adj_5644));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1745 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n60199), .O(n10_adj_5551));   // verilog/coms.v(99[12:25])
    defparam i2_2_lut_3_lut_4_lut_adj_1745.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1746 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(n54578), .I3(GND_net), .O(n60695));
    defparam i1_2_lut_3_lut_adj_1746.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1747 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n60268));
    defparam i1_2_lut_3_lut_adj_1747.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52097 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n71404));
    defparam byte_transmit_counter_0__bdd_4_lut_52097.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1748 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[10] [4]), 
            .O(n60711));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1748.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1749 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[8][2] ), .I3(n10_adj_5634), .O(n1516));   // verilog/coms.v(88[17:63])
    defparam i5_3_lut_4_lut_adj_1749.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1750 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n60565), .I3(n60082), .O(n8_adj_5610));   // verilog/coms.v(100[12:26])
    defparam i3_3_lut_4_lut_adj_1750.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1751 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n60217), .O(n26041));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1751.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1752 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n28429), .O(n60723));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1752.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut_adj_1753 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [0]), 
            .I2(n60164), .I3(GND_net), .O(n32));   // verilog/coms.v(77[16:43])
    defparam i5_2_lut_3_lut_adj_1753.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1754 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[11][3] ), .I3(\data_out_frame[4] [7]), .O(n60139));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1754.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1755 (.I0(\data_in_frame[1][0] ), .I1(Kp_23__N_767), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[3][0] ), .O(n28694));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1755.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1756 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[13] [0]), .I3(\data_out_frame[12] [6]), 
            .O(n14_adj_5619));   // verilog/coms.v(88[17:63])
    defparam i5_3_lut_4_lut_adj_1756.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1757 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n27770));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1757.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1758 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[3]_c [5]), .O(n64129));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1758.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1759 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(n60062), .O(n60708));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1759.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1760 (.I0(n55546), .I1(\data_out_frame[20] [5]), 
            .I2(n55776), .I3(GND_net), .O(n6_adj_5354));
    defparam i1_2_lut_3_lut_adj_1760.LUT_INIT = 16'h6969;
    SB_LUT4 i13591_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[2]), 
            .I3(\data_in_frame[5][2] ), .O(n31536));
    defparam i13591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1761 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[20] [4]), 
            .I2(n60452), .I3(GND_net), .O(n60692));
    defparam i1_2_lut_3_lut_adj_1761.LUT_INIT = 16'h9696;
    SB_LUT4 i13588_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[1]), 
            .I3(\data_in_frame[5][1] ), .O(n31533));
    defparam i13588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13585_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[0]), 
            .I3(\data_in_frame[5][0] ), .O(n31530));
    defparam i13585_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13606_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[7]), 
            .I3(\data_in_frame[5][7] ), .O(n31551));
    defparam i13606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13603_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[6]), 
            .I3(\data_in_frame[5][6] ), .O(n31548));
    defparam i13603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13600_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[5]), 
            .I3(\data_in_frame[5][5] ), .O(n31545));
    defparam i13600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71404_bdd_4_lut (.I0(n71404), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71407));
    defparam n71404_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13597_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[4]), 
            .I3(\data_in_frame[5][4] ), .O(n31542));
    defparam i13597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1762 (.I0(\data_out_frame[22] [7]), .I1(n41_adj_5577), 
            .I2(n46), .I3(n42_adj_5576), .O(n60672));
    defparam i1_2_lut_4_lut_adj_1762.LUT_INIT = 16'h6996;
    SB_LUT4 i13594_3_lut_4_lut (.I0(n8_c), .I1(n60032), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n31539));
    defparam i13594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1763 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2][2] ), .I3(GND_net), .O(n28463));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1763.LUT_INIT = 16'h9696;
    SB_LUT4 equal_2036_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5675));   // verilog/coms.v(169[9:87])
    defparam equal_2036_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1764 (.I0(n28205), .I1(n60490), .I2(n60345), 
            .I3(n60424), .O(n60782));
    defparam i2_3_lut_4_lut_adj_1764.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1765 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1][0] ), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n26037));
    defparam i1_3_lut_adj_1765.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1766 (.I0(n26037), .I1(n62747), .I2(n55167), 
            .I3(n27900), .O(n22_adj_5676));
    defparam i9_4_lut_adj_1766.LUT_INIT = 16'h0020;
    SB_LUT4 i7_4_lut_adj_1767 (.I0(\data_in_frame[2][0] ), .I1(n10_adj_5675), 
            .I2(n60211), .I3(\data_in_frame[1]_c [2]), .O(n20_adj_5677));
    defparam i7_4_lut_adj_1767.LUT_INIT = 16'h2100;
    SB_LUT4 i11_4_lut_adj_1768 (.I0(n28463), .I1(n22_adj_5676), .I2(n16_adj_5426), 
            .I3(n27907), .O(n24_adj_5678));
    defparam i11_4_lut_adj_1768.LUT_INIT = 16'h0040;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n64308), .I1(\data_in_frame[1]_c [3]), 
            .I2(n24_adj_5678), .I3(n20_adj_5677), .O(n6_adj_5679));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'h4000;
    SB_LUT4 i4_4_lut_adj_1770 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n6_adj_5679), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i4_4_lut_adj_1770.LUT_INIT = 16'h8000;
    SB_LUT4 select_789_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52010 (.I0(byte_transmit_counter[1]), 
            .I1(n64902), .I2(n64903), .I3(byte_transmit_counter[2]), .O(n71200));
    defparam byte_transmit_counter_1__bdd_4_lut_52010.LUT_INIT = 16'he4aa;
    SB_LUT4 n71200_bdd_4_lut (.I0(n71200), .I1(n64912), .I2(n64911), .I3(byte_transmit_counter[2]), 
            .O(n71203));
    defparam n71200_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51927 (.I0(byte_transmit_counter[1]), 
            .I1(n64617), .I2(n64618), .I3(byte_transmit_counter[2]), .O(n71194));
    defparam byte_transmit_counter_1__bdd_4_lut_51927.LUT_INIT = 16'he4aa;
    SB_LUT4 n71194_bdd_4_lut (.I0(n71194), .I1(n64606), .I2(n64605), .I3(byte_transmit_counter[2]), 
            .O(n71197));
    defparam n71194_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51922 (.I0(byte_transmit_counter[1]), 
            .I1(n64710), .I2(n64711), .I3(byte_transmit_counter[2]), .O(n71188));
    defparam byte_transmit_counter_1__bdd_4_lut_51922.LUT_INIT = 16'he4aa;
    SB_LUT4 n71188_bdd_4_lut (.I0(n71188), .I1(n64699), .I2(n64698), .I3(byte_transmit_counter[2]), 
            .O(n71191));
    defparam n71188_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51917 (.I0(byte_transmit_counter[1]), 
            .I1(n64620), .I2(n64621), .I3(byte_transmit_counter[2]), .O(n71182));
    defparam byte_transmit_counter_1__bdd_4_lut_51917.LUT_INIT = 16'he4aa;
    SB_LUT4 n71182_bdd_4_lut (.I0(n71182), .I1(n64723), .I2(n64722), .I3(byte_transmit_counter[2]), 
            .O(n71185));
    defparam n71182_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1771 (.I0(n161), .I1(n60002), .I2(n10_adj_5617), 
            .I3(GND_net), .O(n60036));
    defparam i1_2_lut_3_lut_adj_1771.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51912 (.I0(byte_transmit_counter[1]), 
            .I1(n64890), .I2(n64891), .I3(byte_transmit_counter[2]), .O(n71176));
    defparam byte_transmit_counter_1__bdd_4_lut_51912.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1772 (.I0(n161), .I1(n60002), .I2(n10), 
            .I3(GND_net), .O(n60032));
    defparam i1_2_lut_3_lut_adj_1772.LUT_INIT = 16'hfdfd;
    SB_LUT4 n71176_bdd_4_lut (.I0(n71176), .I1(n64615), .I2(n64614), .I3(byte_transmit_counter[2]), 
            .O(n71179));
    defparam n71176_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_314_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10));   // verilog/coms.v(158[12:15])
    defparam equal_314_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_306_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5617));   // verilog/coms.v(158[12:15])
    defparam equal_306_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1773 (.I0(\data_out_frame[20] [3]), .I1(n55641), 
            .I2(\data_out_frame[22] [5]), .I3(n55776), .O(n55665));
    defparam i1_2_lut_3_lut_4_lut_adj_1773.LUT_INIT = 16'h6996;
    SB_LUT4 i13905_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n31850));
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13908_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n31853));
    defparam i13908_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51907 (.I0(byte_transmit_counter[1]), 
            .I1(n64908), .I2(n64909), .I3(byte_transmit_counter[2]), .O(n71170));
    defparam byte_transmit_counter_1__bdd_4_lut_51907.LUT_INIT = 16'he4aa;
    SB_LUT4 n71170_bdd_4_lut (.I0(n71170), .I1(n64888), .I2(n64887), .I3(byte_transmit_counter[2]), 
            .O(n71173));
    defparam n71170_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13911_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n31856));
    defparam i13911_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13914_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n31859));
    defparam i13914_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13917_3_lut_4_lut (.I0(n8_c), .I1(n60036), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n31862));
    defparam i13917_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.n1(n1_adj_7), .tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data}), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), 
            .r_Clock_Count({r_Clock_Count}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n29824(n29824), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n59688(n59688), 
            .n31480(n31480), .tx_active(tx_active), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n63187(n63187), .n27(n27), .n32074(n32074), .n71705(n71705), 
            .n63177(n63177), .n5235(n5235), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), .n29(n29), .n23(n23_adj_8), 
            .n61652(n61652), .n6(n6), .n60832(n60832), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.n31953(n31953), .rx_data({rx_data}), .clk16MHz(clk16MHz), 
            .baudrate({baudrate}), .GND_net(GND_net), .n31945(n31945), 
            .n27632(n27632), .VCC_net(VCC_net), .\r_SM_Main[2] (\r_SM_Main[2]_adj_9 ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29(n29), .n23(n23_adj_8), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), 
            .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), .r_Clock_Count({r_Clock_Count_adj_22}), 
            .n31702(n31702), .\r_SM_Main[1] (\r_SM_Main[1]_adj_18 ), .n29821(n29821), 
            .r_Bit_Index({r_Bit_Index}), .n32083(n32083), .n55814(n55814), 
            .rx_data_ready(rx_data_ready), .n32231(n32231), .n32087(n32087), 
            .n32021(n32021), .n32020(n32020), .n31961(n31961), .n6(n6_adj_20), 
            .n5232(n5232), .n4(n4), .n59686(n59686), .n63199(n63199), 
            .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), .n4_adj_5(n4_adj_21), 
            .n63175(n63175), .n41584(n41584), .n29817(n29817), .n60834(n60834)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n1, tx_o, clk16MHz, tx_data, r_SM_Main, \r_SM_Main_2__N_3536[1] , 
            r_Clock_Count, GND_net, VCC_net, n29824, \r_Bit_Index[0] , 
            n59688, n31480, tx_active, \r_SM_Main_2__N_3545[0] , n63187, 
            n27, n32074, n71705, n63177, n5235, \o_Rx_DV_N_3488[12] , 
            \o_Rx_DV_N_3488[24] , n29, n23, n61652, n6, n60832, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    output n1;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    output [8:0]r_Clock_Count;
    input GND_net;
    input VCC_net;
    output n29824;
    output \r_Bit_Index[0] ;
    output n59688;
    input n31480;
    output tx_active;
    input \r_SM_Main_2__N_3545[0] ;
    input n63187;
    input n27;
    input n32074;
    input n71705;
    output n63177;
    input n5235;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n29;
    input n23;
    input n61652;
    output n6;
    output n60832;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n3, n24885;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n23908, n31164;
    wire [8:0]n41;
    
    wire n3_adj_5290;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n64671, n64672, n71344, n53506, n53505, n53504, n53503, 
        n53502, n53501, n53500, n53499, n64714, n64713, o_Tx_Serial_N_3598;
    wire [2:0]n460;
    
    wire n31147, n23907, n60976, n67713, n67710, n63155, n63161;
    
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n23908), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i51794_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3536[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n31164));
    defparam i51794_4_lut.LUT_INIT = 16'h1115;
    SB_DFFESR r_Clock_Count_2057__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5290), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n24885), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n64671), 
            .I2(n64672), .I3(r_Bit_Index[2]), .O(n71344));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 r_Clock_Count_2057_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n53506), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2057_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n53505), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_9 (.CI(n53505), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n53506));
    SB_LUT4 r_Clock_Count_2057_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n53504), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_8 (.CI(n53504), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n53505));
    SB_LUT4 r_Clock_Count_2057_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n53503), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_7 (.CI(n53503), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n53504));
    SB_LUT4 r_Clock_Count_2057_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n53502), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_6 (.CI(n53502), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n53503));
    SB_LUT4 r_Clock_Count_2057_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n53501), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_5 (.CI(n53501), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n53502));
    SB_LUT4 r_Clock_Count_2057_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n53500), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_4 (.CI(n53500), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n53501));
    SB_LUT4 r_Clock_Count_2057_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n53499), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_3 (.CI(n53499), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n53500));
    SB_LUT4 r_Clock_Count_2057_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2057_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2057_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n53499));
    SB_LUT4 n71344_bdd_4_lut (.I0(n71344), .I1(n64714), .I2(n64713), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3598));
    defparam n71344_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_2057__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2057__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n31164));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n29824), 
            .D(n460[1]), .R(n31147));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n29824), 
            .D(n460[2]), .R(n31147));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59688));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n31480));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i6298_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n63187), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n23907));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i6298_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i6299_3_lut (.I0(n23907), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n23908));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i6299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41754_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n60976));
    defparam i41754_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3598), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i45443_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64713));
    defparam i45443_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n32074));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n71705));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i45444_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64714));
    defparam i45444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45402_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64672));
    defparam i45402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45401_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64671));
    defparam i45401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51896_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n29824));
    defparam i51896_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i1_3_lut_4_lut (.I0(n59688), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n63177));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i49388_3_lut (.I0(n5235), .I1(\o_Rx_DV_N_3488[12] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n67713));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49388_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i49385_4_lut (.I0(n67713), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67710));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49385_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n67710), .I1(n61652), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5290));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n24885));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n61652), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i2340_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2340_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i41617_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n60832));
    defparam i41617_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5235), .I2(n59688), 
            .I3(GND_net), .O(n63155));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), .I3(n63155), 
            .O(n63161));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1083 (.I0(n63161), .I1(n60976), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n31147));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'h0323;
    SB_LUT4 i2333_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2333_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n31953, rx_data, clk16MHz, baudrate, GND_net, n31945, 
            n27632, VCC_net, \r_SM_Main[2] , r_Rx_Data, RX_N_2, \o_Rx_DV_N_3488[24] , 
            n27, n29, n23, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , r_Clock_Count, n31702, 
            \r_SM_Main[1] , n29821, r_Bit_Index, n32083, n55814, rx_data_ready, 
            n32231, n32087, n32021, n32020, n31961, n6, n5232, 
            n4, n59686, n63199, \r_SM_Main_2__N_3446[1] , n4_adj_5, 
            n63175, n41584, n29817, n60834) /* synthesis syn_module_defined=1 */ ;
    input n31953;
    output [7:0]rx_data;
    input clk16MHz;
    input [31:0]baudrate;
    input GND_net;
    input n31945;
    output n27632;
    input VCC_net;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n29;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output [7:0]r_Clock_Count;
    input n31702;
    output \r_SM_Main[1] ;
    output n29821;
    output [2:0]r_Bit_Index;
    input n32083;
    input n55814;
    output rx_data_ready;
    input n32231;
    input n32087;
    input n32021;
    input n32020;
    input n31961;
    output n6;
    input n5232;
    output n4;
    output n59686;
    input n63199;
    input \r_SM_Main_2__N_3446[1] ;
    output n4_adj_5;
    output n63175;
    output n41584;
    output n29817;
    output n60834;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n3165, n19;
    wire [23:0]n8272;
    
    wire n2952, n1459, n53256, n3061;
    wire [23:0]n8298;
    wire [23:0]n294;
    
    wire n3166, n70618, n1262, n70490, n3062, n3167, n2240;
    wire [23:0]n8116;
    
    wire n2366;
    wire [23:0]n8142;
    
    wire n2489, n3063, n3168, n3055, n3160, n13, n21, n2488, 
        n23_c, n2484, n31, n53257, n2953, n1460, n53255, n15, 
        n17, n2954, n1011, n53254, n1838;
    wire [23:0]n8038;
    
    wire n1973, n60868, n60872, n2955, n856, n53253, n2956, n698, 
        n53252, n2957, n858, n53251, n29_c, n63995, n63991, n3159, 
        n31_adj_5020;
    wire [23:0]n8064;
    
    wire n2105;
    wire [23:0]n8090;
    
    wire n2234, n63997, n63845, n63993, n27751, n2360, n68082, 
        n2483, n63905, n63773, n64541, n64569, n60900, n63771, 
        n63769, n64573, n11, n9, n3171, n69094, n27739, n61130, 
        n2490, n19_adj_5021, n69830, n23_adj_5022, n21_adj_5023, n69826, 
        n27_c, n25, n68086, n3172, n6_c, n70378, n25_adj_5024, 
        n68523, n14, n37, n32, n70379;
    wire [23:0]n8168;
    
    wire n2603, n803, n9628, n23826, n46, n35, n33, n68070, 
        n12, n68065, n70730, n29_adj_5025, n27_adj_5026, n68516, 
        n70233, n8, n70380, n37_adj_5027, n35_adj_5028, n33_adj_5029, 
        n70338, n70381, n68113, n69070, n10, n69852, n70231, n70167, 
        n70875, n70372, n2491, n18, n41, n70155, n43, n70156, 
        n70895, n3155, n70896, n27648;
    wire [23:0]n8194;
    
    wire n2720, n3154, n70888, n3153, n70661, n60874, n33_adj_5030, 
        n3152, n70662, n3151, n48, n1415;
    wire [23:0]n7960;
    
    wire n1559, n68519, n69489;
    wire [23:0]n7986;
    
    wire n1700, n24, n26, n63395, n70703, n2713, n63069, n2845, 
        n63073, n538, n61122, n64485, n45, n69158, n63423, n64413, 
        n64489, n63623, n64561, n22, n30, n70769, n2353, n63063, 
        n20, n68514, n70633, n70634, n70468, n39, n69491, n64445, 
        n64549, n68014, n70911, n63635, n64531, n48_adj_5031, n962, 
        n70217;
    wire [23:0]n8246;
    
    wire n2827, n3084, n53250, n2828, n2977, n53249, n69156, n2829, 
        n2867, n53248, n70219, n2830, n2754, n53247, n2831, n2638, 
        n53246, n70882, n63071, n2832, n2519, n53245, n2833, n2397, 
        n53244, n27742, n2834, n2272, n53243, n2612, n2729;
    wire [23:0]n8220;
    
    wire n2843, n2938, n3046, n2946, n3054, n2939, n3047, n2941, 
        n3049, n2940, n3048, n2944, n3052, n35_adj_5032, n2945, 
        n3053, n33_adj_5033, n70822, n1831, n63059, n1977, n64503, 
        n2943, n3051, n37_adj_5034, n2947, n2948, n3056, n27_adj_5035, 
        n29_adj_5036, n2949, n3057, n44, n959, n9799, n23869, 
        n46_adj_5037, n1111, n2950, n3058, n44_adj_5038, n23_adj_5039, 
        n25_adj_5040, n44_adj_5041, n2942, n3050, n39_adj_5042, n3064, 
        n3065, n11_adj_5043, n2951, n3059, n13_adj_5044, n21_adj_5045, 
        n3060, n15_adj_5046, n17_adj_5047, n19_adj_5048, n1112, n31_adj_5049, 
        n68188;
    wire [23:0]n7908;
    
    wire n1261, n69251, n69886, n69880, n68192, n2835, n2144, 
        n53242, n2836, n2013, n53241, n1113, n43_adj_5050, n2714, 
        n2837, n1879, n53240, n2838, n1742, n53239, n2839, n1602, 
        n53238, n3066, n8_adj_5051, n70101, n2840, n53237, n70102, 
        n2841, n53236, n2842, n53235, n53234, n16, n34, n68171, 
        n14_adj_5052, n68167, n70728, n69202, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n2844, n53233, n10_adj_5053, n70107, r_Rx_Data_R, n70108, 
        n1116, n38, n68206, n69227, n53232, n40, n42, n61126;
    wire [23:0]n7934;
    
    wire n1408, n12_adj_5054, n20_adj_5055, n69200, n70248, n70873, 
        n68806, n70615, n33_adj_5056, n69848, n70897, n53231, n53230, 
        n70616, n2715, n53229, n2716, n53228, n2717, n53227, n70898, 
        n2718, n53226, n70892, n70886, n2719, n53225, n69850, 
        n53224, n2721, n53223, n2722, n53222, n2232, n2358, n52683, 
        n1267, n1414, n2723, n53221, n52682, n63051, n2724, n53220, 
        n2481, n2725, n53219, n2601, n2726, n53218, n2727, n53217, 
        n34_adj_5058, n2728, n53216, n53215, n2730, n53214, n70761, 
        n2596, n63067, n1558, n53213, n52681, n63107, n2597, n53212, 
        n2598, n53211, n52680;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n52679, n63105, n2599, n53210, n1699, n52678, n63103, 
        n2600, n53209, n52677, n53208, n2602, n53207, n41_adj_5061, 
        n70189, n27736, n43_adj_5062, n70190, n39_adj_5063, n68773, 
        n69678, n36, n38_adj_5064, n53206;
    wire [23:0]n8012;
    
    wire n1837, n52676, n63101, n37_adj_5065, n39_adj_5066, n2604, 
        n53205, n52675, n63099, n41_adj_5067, n2605, n53204, n2606, 
        n53203, n52674, n63049, n2607, n53202, n2608, n53201, 
        n45_adj_5068, n69116, n52673, n63097, n1972, n2609, n53200, 
        n2610, n53199, n31_adj_5069, n2611, n53198, n2104, n43_adj_5070, 
        n52672, n53197, n63847, n61134, n2476, n53196, n52671, 
        n2233, n2477, n53195, n52670, n2478, n53194, n2479, n53193, 
        n2359, n52669, n2482, n2480, n53192, n70203, n53191, n52668, 
        n53190, n61158, n53189, n53188, n52667, n2485, n53187, 
        n2486, n53186, n52666, n2487, n53185, n53184, n53183, 
        n52665, n53182, n53181, n63065, n61138, n53180, n2354, 
        n53179, n52664, n2355, n53178, n2356, n53177, n2357, n53176, 
        n35_adj_5071, n961, n23867, n68022, n48_adj_5072, n804, 
        n53175, n1701, n32_adj_5073, n39_adj_5074, n70181, n41_adj_5075, 
        n70182, n37_adj_5076, n68730, n69654, n34_adj_5077, n70207, 
        n53174, n43_adj_5078, n69121, n70483, n1694, n70484, n1693, 
        n48_adj_5079, n63889, n63875, n63877, n63865, n63821, n27715, 
        n1841, n1976, n2108, n2237, n2363, n27_adj_5080, n52663, 
        n53173, n2361, n53172, n2362, n53171, n53170, n1560, n1839, 
        n2364, n53169, n2365, n53168, n1974, n2106, n2235, n53167, 
        n63903, n63009, n63007, n63893, n2367, n53166, n61142, 
        n2227, n53165, n2228, n53164, n17_adj_5081, n2229, n53163, 
        n23_adj_5082, n21_adj_5083, n19_adj_5084, n68493, n29_adj_5085, 
        n27_adj_5086, n25_adj_5087, n68480, n35_adj_5088, n33_adj_5089, 
        n31_adj_5090, n70334, n16_adj_5091, n2230, n53162, n2231, 
        n53161, n52662, n53160, n53159, n53158, n53157, n2236, 
        n53156, n2109, n42_adj_5092, n960, n53155, n2238, n53154, 
        n2239, n53153, n53152, n63061, n61146, n2098, n53151, 
        n29_adj_5093, n2099, n53150, n42_adj_5094, n2100, n53149, 
        n2101, n53148, n2102, n53147, n41_adj_5095, n15_adj_5096, 
        n41_adj_5097, n1263, n39_adj_5098, n2103, n53146, n53145, 
        n37_adj_5099, n35_adj_5100, n39_adj_5101, n37_adj_5102, n53144, 
        n53143, n52661, n1410, n29_adj_5103, n39_adj_5104, n70151, 
        n31_adj_5105, n2107, n53142, n53141, n52660, n35_adj_5106, 
        n1554, n35_adj_5107, n23_adj_5108, n21_adj_5109, n19_adj_5110, 
        n68333, n1695, n53140, n23_adj_5111, n29_adj_5112, n25_adj_5113, 
        n2110, n27_adj_5114, n13_adj_5115, n15_adj_5116, n1966, n53139, 
        n33_adj_5117, n1967, n53138, n17_adj_5118, n1833, n31_adj_5119, 
        n19_adj_5120, n21_adj_5121, n1968, n53137, n61968, n33_adj_5122, 
        n68272, n1969, n53136, n1970, n53135, n69317, n69926, 
        n1971, n53134, n69922, n68276, n53133, n53132, n10_adj_5123, 
        n17_adj_5124, n69375;
    wire [7:0]n1;
    
    wire n29942, n31162, n41_adj_5126, n70152, n70121, n70122, n71701, 
        n18_adj_5127, n36_adj_5128, n68262, n53131, n3_adj_5129, n1975, 
        n53130, n53129, n53128, n68489, n69449, n53127, n16_adj_5130, 
        n68258, n70649, n1832, n53126, n69190, n69950, n37_adj_5131, 
        n35_adj_5132, n25_adj_5133, n69944, n1836, n37_adj_5134, n22_adj_5135, 
        n70220, n43_adj_5136, n69168, n53125, n20_adj_5137, n28, 
        n18_adj_5138, n68476, n70635, n70636, n70464, n37_adj_5139, 
        n69455, n1834, n53124, n70461, n69166, n70760, n31_adj_5140, 
        n29_adj_5141, n63797, n63601, n63621, n14_adj_5142, n22_adj_5143, 
        n12_adj_5144, n68292, n70647, n68335, n70648, n70434, n1835, 
        n53123, n63849, n63891, n37_adj_5145, n25_adj_5146, n23_adj_5147, 
        n21_adj_5148, n68397, n53122, n19_adj_5149, n17_adj_5150, 
        n69431, n69978, n27_adj_5151, n69972, n68399, n14_adj_5152, 
        n70145, n53121, n53120, n39_adj_5153, n70292, n53119, n1840, 
        n53118, n53117, n70833, n69188, n43_adj_5154, n61155, n12_adj_5162, 
        n70893, n70894, n70141, n53467, n41_adj_5163, n31_adj_5164, 
        n33_adj_5165, n35_adj_5166, n39_adj_5167, n70146, n22_adj_5168, 
        n45_adj_5169, n40_adj_5170, n43_adj_5171, n41_adj_5172, n68387, 
        n20_adj_5173, n68381, n70222, n69178, n18_adj_5174, n26_adj_5175, 
        n29_adj_5176, n68707, n53466, n53465, n53464, n53463, n53462, 
        n53461, n16_adj_5177, n68415, n70637, n64527, n64529, n53106, 
        n53105, n53104, n1696, n53103, n20_adj_5178, n38_adj_5179, 
        n32_adj_5180, n40_adj_5181, n28_adj_5182, n1697, n53102, n70142, 
        n70177, n70178, n1698, n53101, n68686, n53100, n53099, 
        n68323, n30_adj_5183, n68683, n70613, n18_adj_5184, n68321, 
        n70607, n69124, n70821, n69184, n53098, n41_adj_5185, n39_adj_5186, 
        n29_adj_5187, n16_adj_5188, n24_adj_5189, n31_adj_5190, n14_adj_5191, 
        n68349, n70639, n33_adj_5192, n1702, n70640;
    wire [2:0]n479;
    
    wire n31149, n70456, n27_adj_5193, n70310, n68670, n70819, n69182, 
        n30_adj_5194, n38_adj_5195, n70881, n26_adj_5196, n70175, 
        n1552, n53097, n1553, n53096, n1557, n70176, n68653, n28_adj_5197, 
        n68650, n70625, n69126, n70825, n70826, n70767, n48_adj_5198, 
        n23_adj_5199, n25_adj_5200, n805, n42_adj_5201, n43_adj_5202, 
        n33_adj_5203, n27_adj_5204, n21_adj_5205, n68561, n41_adj_5206, 
        n39_adj_5207, n68556, n37_adj_5208, n70497, n23_adj_5209, 
        n29_adj_5210, n27_adj_5211, n25_adj_5212, n68602, n20_adj_5213, 
        n26_adj_5214, n28_adj_5215, n35_adj_5216, n31_adj_5217, n68594, 
        n24_adj_5218, n32_adj_5219, n22_adj_5220, n68552, n70631, 
        n22_adj_5221, n70632, n70472, n70498, n28_adj_5222, n30_adj_5223, 
        n70344, n68558, n70726, n69152, n70823, n1115, n1265, 
        n70638, n70460, n70824, n53095, n1555, n53094, n70322, 
        n70701, n1412, n1556, n69176, n53093, n53092, n53091, 
        n53090, n53089, n64363, n48_adj_5224, n53088, n1409, n53087, 
        n53086, n1411, n53085, n53084, n1413, n53083, n53082, 
        n53081, n63057, n61164, n53080, n26_adj_5225, n34_adj_5226, 
        n53079, n53078, n1264, n53077, n53076, n1266, n53075, 
        n53074, n63055, n61168, n53073, n63627, n64447, n53072, 
        n53071, n1114, n53070, n53069, n53068, n63053, n61172, 
        n24_adj_5227, n68592, n70629;
    wire [23:0]n8324;
    
    wire n3186, n53314, n3082, n53313, n3188, n53312, n53311, 
        n53310, n3156, n53309, n3157, n53308, n3158, n53307, n53306, 
        n53305, n3161, n53304, n3162, n53303, n3163, n53302, n3164, 
        n53301, n53300, n53299, n53298, n53297, n3169, n53296, 
        n3170, n53295, n53294, n53293, n63077, n53292, n61114, 
        n53291, n53290, n53289, n53288, n53287, n53286, n53285, 
        n53284, n53283, n53282, n53281, n53280, n53279, n53278, 
        n53277, n53276, n53275, n53274, n53273, n53272, n53271, 
        n70630, n63075, n61118, n53270, n53269, n53268, n53267, 
        n53266, n53265, n53264, n53263, n53262, n53261, n63785, 
        n3_adj_5229, n63789, n53260, n53259, n5, n67700, n63793, 
        n59720, n67706, n8_adj_5230, n67697, n67703, n53258, n64431, 
        n64553, n2, n10015, n70474, n70350, n68600, n70386, n69146, 
        n31_adj_5231, n29_adj_5232, n33_adj_5233, n35_adj_5234, n39_adj_5235, 
        n37_adj_5236, n41_adj_5237, n63895, n63625, n63629, n63631, 
        n70611, n63633, n63637, n41626, n41624, n23812, n9792, 
        n70612, n28_adj_5238, n68621, n30_adj_5239, n59971, n14_adj_5240, 
        n15_adj_5241, n43_adj_5242, n27748, n67642, n67639, n67636, 
        n63131, n63137, n63897, n64473, n63807, n61175, n42_adj_5244, 
        n63775, n70491, n67685, n70492, n48_adj_5245, n63833, n63835, 
        n27700, n37_adj_5246, n41_adj_5247, n39_adj_5248, n67656, 
        n67653, n63765, n63743, n63843, n46_adj_5249, n48_adj_5250, 
        n27694, n32_adj_5251, n64475, n70183, n70184, n68753, n69662, 
        n34_adj_5252, n70205, n69118, n70485, n40_adj_5253, n70486, 
        n63167, n63173, n41_adj_5254, n39_adj_5255, n33_adj_5256, 
        n35_adj_5257, n37_adj_5258, n29_adj_5259, n31_adj_5260, n23_adj_5261, 
        n25_adj_5262, n45_adj_5263, n7, n9_adj_5264, n17_adj_5265, 
        n19_adj_5266, n21_adj_5267, n43_adj_5268, n70765, n27724, 
        n11_adj_5269, n13_adj_5270, n15_adj_5271, n27_adj_5272, n67971, 
        n67979, n16_adj_5273, n41_adj_5274, n67936, n8_adj_5275, n24_adj_5276, 
        n3274, n68025, n69019, n69007, n70431, n69772, n70673, 
        n12_adj_5277, n4_adj_5278, n70366, n70367, n67955, n10_adj_5279, 
        n30_adj_5280, n36_adj_5281, n67961, n70732, n70243, n70877, 
        n70878, n38_adj_5282, n40_adj_5283, n6_adj_5284, n68788, n70617, 
        n70370, n70371, n67941, n69854, n70241, n70814, n67943, 
        n70521, n40_adj_5285, n63029, n3253, n70523, n63037, n64493, 
        n64419, n62985, n64525, n62075, n63339, n63357, n27_adj_5286, 
        n68642, n64563, n38_adj_5287, n61643, n61149, n63647, n26_adj_5288, 
        n70171, n70172, n68630, n70627, n69134, n70827, n70828, 
        n63649, n64337, n48_adj_5289, n63899, n63691, n67620, n63907, 
        n67621;
    
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n31953));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2761_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n53256), 
            .O(n8272[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n31945));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8298[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51220_3_lut (.I0(n70618), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n70490));   // verilog/uart_rx.v(119[33:55])
    defparam i51220_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8298[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8116[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8142[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8298[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8298[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2761_8 (.CI(n53256), .I0(n2952), .I1(n1459), .CO(n53257));
    SB_LUT4 add_2761_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n53255), 
            .O(n8272[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_7 (.CI(n53255), .I0(n2953), .I1(n1460), .CO(n53256));
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2761_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n53254), 
            .O(n8272[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_6 (.CI(n53254), .I0(n2954), .I1(n1011), .CO(n53255));
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8038[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i534_3_lut (.I0(n60868), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n60872));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 add_2761_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n53253), 
            .O(n8272[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_5 (.CI(n53253), .I0(n2955), .I1(n856), .CO(n53254));
    SB_LUT4 add_2761_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n53252), 
            .O(n8272[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_4 (.CI(n53252), .I0(n2956), .I1(n698), .CO(n53253));
    SB_LUT4 add_2761_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n53251), 
            .O(n8272[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_3 (.CI(n53251), .I0(n2957), .I1(n858), .CO(n53252));
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63995));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_994 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63991));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8064[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8090[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n63995), .I1(n63997), .I2(n63845), .I3(n63993), 
            .O(n27751));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8116[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48812_4_lut (.I0(n29_c), .I1(n17), .I2(n15), .I3(n13), 
            .O(n68082));
    defparam i48812_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8142[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45308_4_lut (.I0(n63905), .I1(baudrate[20]), .I2(n63773), 
            .I3(n64541), .O(n64569));
    defparam i45308_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51677_4_lut (.I0(n60900), .I1(n63771), .I2(n64569), .I3(n63769), 
            .O(n64573));
    defparam i51677_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i49824_4_lut (.I0(n11), .I1(n9), .I2(n3171), .I3(baudrate[2]), 
            .O(n69094));
    defparam i49824_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i41907_1_lut (.I0(n27739), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61130));
    defparam i41907_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50560_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n69094), 
            .O(n69830));
    defparam i50560_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50556_4_lut (.I0(n23_adj_5022), .I1(n21_adj_5023), .I2(n19), 
            .I3(n69830), .O(n69826));
    defparam i50556_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48816_4_lut (.I0(n29_c), .I1(n27_c), .I2(n25), .I3(n69826), 
            .O(n68086));
    defparam i48816_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51108_3_lut (.I0(n6_c), .I1(baudrate[13]), .I2(n29_c), .I3(GND_net), 
            .O(n70378));   // verilog/uart_rx.v(119[33:55])
    defparam i51108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49253_4_lut (.I0(n25_adj_5024), .I1(n23_c), .I2(n21), .I3(n19_adj_5021), 
            .O(n68523));
    defparam i49253_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14), .I1(baudrate[17]), 
            .I2(n37), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51109_3_lut (.I0(n70378), .I1(baudrate[14]), .I2(n31_adj_5020), 
            .I3(GND_net), .O(n70379));   // verilog/uart_rx.v(119[33:55])
    defparam i51109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8168[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4048_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9628), .I3(n23826), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i4048_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 i48800_4_lut (.I0(n35), .I1(n33), .I2(n31_adj_5020), .I3(n68082), 
            .O(n68070));
    defparam i48800_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51460_4_lut (.I0(n32), .I1(n12), .I2(n37), .I3(n68065), 
            .O(n70730));   // verilog/uart_rx.v(119[33:55])
    defparam i51460_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49246_4_lut (.I0(n31), .I1(n29_adj_5025), .I2(n27_adj_5026), 
            .I3(n68523), .O(n68516));
    defparam i49246_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50963_3_lut (.I0(n70379), .I1(baudrate[15]), .I2(n33), .I3(GND_net), 
            .O(n70233));   // verilog/uart_rx.v(119[33:55])
    defparam i50963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51110_3_lut (.I0(n8), .I1(baudrate[10]), .I2(n23_adj_5022), 
            .I3(GND_net), .O(n70380));   // verilog/uart_rx.v(119[33:55])
    defparam i51110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51068_4_lut (.I0(n37_adj_5027), .I1(n35_adj_5028), .I2(n33_adj_5029), 
            .I3(n68516), .O(n70338));
    defparam i51068_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51111_3_lut (.I0(n70380), .I1(baudrate[11]), .I2(n25), .I3(GND_net), 
            .O(n70381));   // verilog/uart_rx.v(119[33:55])
    defparam i51111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49800_4_lut (.I0(n25), .I1(n23_adj_5022), .I2(n21_adj_5023), 
            .I3(n68113), .O(n69070));
    defparam i49800_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50582_3_lut (.I0(n10), .I1(baudrate[9]), .I2(n21_adj_5023), 
            .I3(GND_net), .O(n69852));   // verilog/uart_rx.v(119[33:55])
    defparam i50582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50961_3_lut (.I0(n70381), .I1(baudrate[12]), .I2(n27_c), 
            .I3(GND_net), .O(n70231));   // verilog/uart_rx.v(119[33:55])
    defparam i50961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50897_4_lut (.I0(n35), .I1(n33), .I2(n31_adj_5020), .I3(n68086), 
            .O(n70167));
    defparam i50897_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51605_4_lut (.I0(n70233), .I1(n70730), .I2(n37), .I3(n68070), 
            .O(n70875));   // verilog/uart_rx.v(119[33:55])
    defparam i51605_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51102_4_lut (.I0(n70231), .I1(n69852), .I2(n27_c), .I3(n69070), 
            .O(n70372));   // verilog/uart_rx.v(119[33:55])
    defparam i51102_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50885_3_lut (.I0(n18), .I1(baudrate[13]), .I2(n41), .I3(GND_net), 
            .O(n70155));   // verilog/uart_rx.v(119[33:55])
    defparam i50885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50886_3_lut (.I0(n70155), .I1(baudrate[14]), .I2(n43), .I3(GND_net), 
            .O(n70156));   // verilog/uart_rx.v(119[33:55])
    defparam i50886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51625_4_lut (.I0(n70372), .I1(n70875), .I2(n37), .I3(n70167), 
            .O(n70895));   // verilog/uart_rx.v(119[33:55])
    defparam i51625_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51626_3_lut (.I0(n70895), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n70896));   // verilog/uart_rx.v(119[33:55])
    defparam i51626_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51766_3_lut (.I0(n27648), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n27632));   // verilog/uart_rx.v(119[33:55])
    defparam i51766_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8194[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51618_3_lut (.I0(n70896), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n70888));   // verilog/uart_rx.v(119[33:55])
    defparam i51618_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51391_3_lut (.I0(n70888), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n70661));   // verilog/uart_rx.v(119[33:55])
    defparam i51391_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i639_4_lut (.I0(n60872), .I1(n294[19]), .I2(n46), .I3(baudrate[4]), 
            .O(n60874));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51392_3_lut (.I0(n70661), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n70662));   // verilog/uart_rx.v(119[33:55])
    defparam i51392_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50969_3_lut (.I0(n70662), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i50969_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7960[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50219_4_lut (.I0(n43), .I1(n41), .I2(n29_adj_5025), .I3(n68519), 
            .O(n69489));
    defparam i50219_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7986[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24), .I1(baudrate[7]), 
            .I2(n29_adj_5025), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_995 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n63395));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut (.I0(n70703), .I1(baudrate[18]), .I2(n2713), 
            .I3(n63069), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 add_2761_2_lut (.I0(n61122), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i45224_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n64485));
    defparam i45224_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51864_2_lut_4_lut (.I0(n70703), .I1(baudrate[18]), .I2(n2713), 
            .I3(n27739), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i51864_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i49888_3_lut (.I0(n70156), .I1(baudrate[15]), .I2(n45), .I3(GND_net), 
            .O(n69158));   // verilog/uart_rx.v(119[33:55])
    defparam i49888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_996 (.I0(n60900), .I1(n63395), .I2(n63991), .I3(baudrate[16]), 
            .O(n63423));
    defparam i1_4_lut_adj_996.LUT_INIT = 16'h0004;
    SB_LUT4 i45300_4_lut (.I0(n64485), .I1(n64413), .I2(n64489), .I3(n63623), 
            .O(n64561));
    defparam i45300_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22), .I1(baudrate[9]), 
            .I2(n33_adj_5029), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_997 (.I0(n70769), .I1(baudrate[15]), .I2(n2353), 
            .I3(n63063), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_997.LUT_INIT = 16'h7100;
    SB_LUT4 i51363_4_lut (.I0(n30), .I1(n20), .I2(n33_adj_5029), .I3(n68514), 
            .O(n70633));   // verilog/uart_rx.v(119[33:55])
    defparam i51363_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51364_3_lut (.I0(n70633), .I1(baudrate[10]), .I2(n35_adj_5028), 
            .I3(GND_net), .O(n70634));   // verilog/uart_rx.v(119[33:55])
    defparam i51364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51198_3_lut (.I0(n70634), .I1(baudrate[11]), .I2(n37_adj_5027), 
            .I3(GND_net), .O(n70468));   // verilog/uart_rx.v(119[33:55])
    defparam i51198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50221_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n70338), 
            .O(n69491));
    defparam i50221_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51804_2_lut_4_lut (.I0(n70769), .I1(baudrate[15]), .I2(n2353), 
            .I3(n64445), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i51804_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51641_4_lut (.I0(n64549), .I1(n68014), .I2(n64561), .I3(n63423), 
            .O(n70911));
    defparam i51641_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63635), .I1(n64531), .I2(baudrate[0]), 
            .I3(n48_adj_5031), .O(n962));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i50947_4_lut (.I0(n69158), .I1(n26), .I2(n45), .I3(n69489), 
            .O(n70217));   // verilog/uart_rx.v(119[33:55])
    defparam i50947_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2761_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53251));
    SB_LUT4 add_2760_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n53250), 
            .O(n8246[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2760_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n53249), 
            .O(n8246[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49886_3_lut (.I0(n70468), .I1(baudrate[12]), .I2(n39), .I3(GND_net), 
            .O(n69156));   // verilog/uart_rx.v(119[33:55])
    defparam i49886_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2760_20 (.CI(n53249), .I0(n2828), .I1(n2977), .CO(n53250));
    SB_LUT4 add_2760_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n53248), 
            .O(n8246[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_19 (.CI(n53248), .I0(n2829), .I1(n2867), .CO(n53249));
    SB_LUT4 i50949_4_lut (.I0(n69156), .I1(n70217), .I2(n45), .I3(n69491), 
            .O(n70219));   // verilog/uart_rx.v(119[33:55])
    defparam i50949_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2760_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n53247), 
            .O(n8246[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_18 (.CI(n53247), .I0(n2830), .I1(n2754), .CO(n53248));
    SB_LUT4 add_2760_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n53246), 
            .O(n8246[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_998 (.I0(n70882), .I1(baudrate[19]), .I2(n2827), 
            .I3(n63071), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_998.LUT_INIT = 16'h7100;
    SB_CARRY add_2760_17 (.CI(n53246), .I0(n2831), .I1(n2638), .CO(n53247));
    SB_LUT4 add_2760_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n53245), 
            .O(n8246[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_16 (.CI(n53245), .I0(n2832), .I1(n2519), .CO(n53246));
    SB_LUT4 add_2760_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n53244), 
            .O(n8246[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_15 (.CI(n53244), .I0(n2833), .I1(n2397), .CO(n53245));
    SB_LUT4 i51869_2_lut_4_lut (.I0(n70882), .I1(baudrate[19]), .I2(n2827), 
            .I3(n27742), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i51869_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2760_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n53243), 
            .O(n8246[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8194[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8220[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8272[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8272[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8272[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8272[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8272[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8272[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8272[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_999 (.I0(n70822), .I1(baudrate[11]), .I2(n1831), 
            .I3(n63059), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_999.LUT_INIT = 16'h7100;
    SB_LUT4 i51712_2_lut_4_lut (.I0(n70822), .I1(baudrate[11]), .I2(n1831), 
            .I3(n64503), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i51712_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8272[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8272[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8272[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8272[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i535_4_lut (.I0(n70911), .I1(n44), .I2(n294[20]), .I3(baudrate[2]), 
            .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_CARRY add_2760_14 (.CI(n53243), .I0(n2834), .I1(n2272), .CO(n53244));
    SB_LUT4 i4219_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9799), .I3(n23869), 
            .O(n46_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam i4219_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i742_4_lut (.I0(n60874), .I1(n294[18]), .I2(n46_adj_5037), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8272[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4041_2_lut (.I0(n23826), .I1(n9628), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam i4041_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5038), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4212_2_lut (.I0(n23869), .I1(n9799), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam i4212_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8272[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8272[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8272[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8272[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8272[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8272[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8272[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8272[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5041), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48918_4_lut (.I0(n31_adj_5049), .I1(n19_adj_5048), .I2(n17_adj_5047), 
            .I3(n15_adj_5046), .O(n68188));
    defparam i48918_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7908[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49981_4_lut (.I0(n13_adj_5044), .I1(n11_adj_5043), .I2(n3065), 
            .I3(baudrate[2]), .O(n69251));
    defparam i49981_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50616_4_lut (.I0(n19_adj_5048), .I1(n17_adj_5047), .I2(n15_adj_5046), 
            .I3(n69251), .O(n69886));
    defparam i50616_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50610_4_lut (.I0(n25_adj_5040), .I1(n23_adj_5039), .I2(n21_adj_5045), 
            .I3(n69886), .O(n69880));
    defparam i50610_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48922_4_lut (.I0(n31_adj_5049), .I1(n29_adj_5036), .I2(n27_adj_5035), 
            .I3(n69880), .O(n68192));
    defparam i48922_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2760_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n53242), 
            .O(n8246[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_13 (.CI(n53242), .I0(n2835), .I1(n2144), .CO(n53243));
    SB_LUT4 add_2760_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n53241), 
            .O(n8246[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8220[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2760_12 (.CI(n53241), .I0(n2836), .I1(n2013), .CO(n53242));
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8220[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2760_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n53240), 
            .O(n8246[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_11 (.CI(n53240), .I0(n2837), .I1(n1879), .CO(n53241));
    SB_LUT4 add_2760_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n53239), 
            .O(n8246[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_10 (.CI(n53239), .I0(n2838), .I1(n1742), .CO(n53240));
    SB_LUT4 add_2760_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n53238), 
            .O(n8246[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_9 (.CI(n53238), .I0(n2839), .I1(n1602), .CO(n53239));
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50831_3_lut (.I0(n8_adj_5051), .I1(baudrate[13]), .I2(n31_adj_5049), 
            .I3(GND_net), .O(n70101));   // verilog/uart_rx.v(119[33:55])
    defparam i50831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2760_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n53237), 
            .O(n8246[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50832_3_lut (.I0(n70101), .I1(baudrate[14]), .I2(n33_adj_5033), 
            .I3(GND_net), .O(n70102));   // verilog/uart_rx.v(119[33:55])
    defparam i50832_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2760_8 (.CI(n53237), .I0(n2840), .I1(n1459), .CO(n53238));
    SB_LUT4 add_2760_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n53236), 
            .O(n8246[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_7 (.CI(n53236), .I0(n2841), .I1(n1460), .CO(n53237));
    SB_LUT4 add_2760_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n53235), 
            .O(n8246[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2760_6 (.CI(n53235), .I0(n2842), .I1(n1011), .CO(n53236));
    SB_LUT4 add_2760_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n53234), 
            .O(n8246[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16), .I1(baudrate[17]), 
            .I2(n39_adj_5042), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48901_4_lut (.I0(n37_adj_5034), .I1(n35_adj_5032), .I2(n33_adj_5033), 
            .I3(n68188), .O(n68171));
    defparam i48901_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2760_5 (.CI(n53234), .I0(n2843), .I1(n856), .CO(n53235));
    SB_LUT4 i51458_4_lut (.I0(n34), .I1(n14_adj_5052), .I2(n39_adj_5042), 
            .I3(n68167), .O(n70728));   // verilog/uart_rx.v(119[33:55])
    defparam i51458_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49932_3_lut (.I0(n70102), .I1(baudrate[15]), .I2(n35_adj_5032), 
            .I3(GND_net), .O(n69202));   // verilog/uart_rx.v(119[33:55])
    defparam i49932_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2760_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n53233), 
            .O(n8246[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50837_3_lut (.I0(n10_adj_5053), .I1(baudrate[10]), .I2(n25_adj_5040), 
            .I3(GND_net), .O(n70107));   // verilog/uart_rx.v(119[33:55])
    defparam i50837_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2760_4 (.CI(n53233), .I0(n2844), .I1(n698), .CO(n53234));
    SB_LUT4 i50838_3_lut (.I0(n70107), .I1(baudrate[11]), .I2(n27_adj_5035), 
            .I3(GND_net), .O(n70108));   // verilog/uart_rx.v(119[33:55])
    defparam i50838_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49957_4_lut (.I0(n27_adj_5035), .I1(n25_adj_5040), .I2(n23_adj_5039), 
            .I3(n68206), .O(n69227));
    defparam i49957_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2760_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n53232), 
            .O(n8246[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40), .I1(baudrate[4]), .I2(n43_adj_5050), 
            .I3(GND_net), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2760_3 (.CI(n53232), .I0(n2845), .I1(n858), .CO(n53233));
    SB_LUT4 add_2760_2_lut (.I0(n61126), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2760_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2760_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53232));
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7934[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8220[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5054), .I1(baudrate[9]), 
            .I2(n23_adj_5039), .I3(GND_net), .O(n20_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49930_3_lut (.I0(n70108), .I1(baudrate[12]), .I2(n29_adj_5036), 
            .I3(GND_net), .O(n69200));   // verilog/uart_rx.v(119[33:55])
    defparam i49930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50978_4_lut (.I0(n37_adj_5034), .I1(n35_adj_5032), .I2(n33_adj_5033), 
            .I3(n68192), .O(n70248));
    defparam i50978_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51603_4_lut (.I0(n69202), .I1(n70728), .I2(n39_adj_5042), 
            .I3(n68171), .O(n70873));   // verilog/uart_rx.v(119[33:55])
    defparam i51603_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51345_4_lut (.I0(n42), .I1(n38), .I2(n43_adj_5050), .I3(n68806), 
            .O(n70615));   // verilog/uart_rx.v(119[33:55])
    defparam i51345_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50578_4_lut (.I0(n69200), .I1(n20_adj_5055), .I2(n29_adj_5036), 
            .I3(n69227), .O(n69848));   // verilog/uart_rx.v(119[33:55])
    defparam i50578_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51627_4_lut (.I0(n69848), .I1(n70873), .I2(n39_adj_5042), 
            .I3(n70248), .O(n70897));   // verilog/uart_rx.v(119[33:55])
    defparam i51627_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2759_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n53231), 
            .O(n8220[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2759_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n53230), 
            .O(n8220[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_19 (.CI(n53230), .I0(n2714), .I1(n2867), .CO(n53231));
    SB_LUT4 i51346_3_lut (.I0(n70615), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n70616));   // verilog/uart_rx.v(119[33:55])
    defparam i51346_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2759_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n53229), 
            .O(n8220[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_18 (.CI(n53229), .I0(n2715), .I1(n2754), .CO(n53230));
    SB_LUT4 add_2759_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n53228), 
            .O(n8220[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_17 (.CI(n53228), .I0(n2716), .I1(n2638), .CO(n53229));
    SB_LUT4 add_2759_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n53227), 
            .O(n8220[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_16 (.CI(n53227), .I0(n2717), .I1(n2519), .CO(n53228));
    SB_LUT4 i51628_3_lut (.I0(n70897), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n70898));   // verilog/uart_rx.v(119[33:55])
    defparam i51628_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2759_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n53226), 
            .O(n8220[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1000 (.I0(n70892), .I1(baudrate[20]), .I2(n2938), 
            .I3(n63073), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1000.LUT_INIT = 16'h7100;
    SB_LUT4 i51616_3_lut (.I0(n70898), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n70886));   // verilog/uart_rx.v(119[33:55])
    defparam i51616_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2759_15 (.CI(n53226), .I0(n2718), .I1(n2397), .CO(n53227));
    SB_LUT4 add_2759_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n53225), 
            .O(n8220[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50580_3_lut (.I0(n70886), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n69850));   // verilog/uart_rx.v(119[33:55])
    defparam i50580_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2759_14 (.CI(n53225), .I0(n2719), .I1(n2272), .CO(n53226));
    SB_LUT4 add_2759_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n53224), 
            .O(n8220[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_13 (.CI(n53224), .I0(n2720), .I1(n2144), .CO(n53225));
    SB_LUT4 i51877_2_lut_4_lut (.I0(n70892), .I1(baudrate[20]), .I2(n2938), 
            .I3(n64541), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i51877_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2759_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n53223), 
            .O(n8220[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_12 (.CI(n53223), .I0(n2721), .I1(n2013), .CO(n53224));
    SB_LUT4 add_2759_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n53222), 
            .O(n8220[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8116[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n52683), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_11 (.CI(n53222), .I0(n2722), .I1(n1879), .CO(n53223));
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7934[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2759_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n53221), 
            .O(n8220[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_10 (.CI(n53221), .I0(n2723), .I1(n1742), .CO(n53222));
    SB_LUT4 sub_38_add_2_25_lut (.I0(n63051), .I1(n27632), .I2(VCC_net), 
            .I3(n52682), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2759_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n53220), 
            .O(n8220[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8142[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_25 (.CI(n52682), .I0(n27632), .I1(VCC_net), 
            .CO(n52683));
    SB_CARRY add_2759_9 (.CI(n53220), .I0(n2724), .I1(n1602), .CO(n53221));
    SB_LUT4 add_2759_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n53219), 
            .O(n8220[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8168[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8194[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2759_8 (.CI(n53219), .I0(n2725), .I1(n1459), .CO(n53220));
    SB_LUT4 add_2759_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n53218), 
            .O(n8220[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_7 (.CI(n53218), .I0(n2726), .I1(n1460), .CO(n53219));
    SB_LUT4 add_2759_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n53217), 
            .O(n8220[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2759_6 (.CI(n53217), .I0(n2727), .I1(n1011), .CO(n53218));
    SB_LUT4 add_2759_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n53216), 
            .O(n8220[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_5 (.CI(n53216), .I0(n2728), .I1(n856), .CO(n53217));
    SB_LUT4 add_2759_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n53215), 
            .O(n8220[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_4 (.CI(n53215), .I0(n2729), .I1(n698), .CO(n53216));
    SB_LUT4 add_2759_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n53214), 
            .O(n8220[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2759_3 (.CI(n53214), .I0(n2730), .I1(n858), .CO(n53215));
    SB_LUT4 i1_2_lut_4_lut_adj_1001 (.I0(n70761), .I1(baudrate[17]), .I2(n2596), 
            .I3(n63067), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1001.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7960[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2759_2_lut (.I0(n61130), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2759_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2759_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53214));
    SB_LUT4 add_2758_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n53213), 
            .O(n8194[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n63107), .I1(n64573), .I2(VCC_net), 
            .I3(n52681), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_24 (.CI(n52681), .I0(n64573), .I1(VCC_net), 
            .CO(n52682));
    SB_LUT4 add_2758_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n53212), 
            .O(n8194[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_18 (.CI(n53212), .I0(n2597), .I1(n2754), .CO(n53213));
    SB_LUT4 add_2758_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n53211), 
            .O(n8194[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_17 (.CI(n53211), .I0(n2598), .I1(n2638), .CO(n53212));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n52680), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n52680), .I0(n294[21]), .I1(VCC_net), 
            .CO(n52681));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n63105), .I1(n294[20]), .I2(VCC_net), 
            .I3(n52679), .O(n63107)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2758_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n53210), 
            .O(n8194[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7986[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_22 (.CI(n52679), .I0(n294[20]), .I1(VCC_net), 
            .CO(n52680));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n63103), .I1(n294[19]), .I2(VCC_net), 
            .I3(n52678), .O(n63105)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2758_16 (.CI(n53210), .I0(n2599), .I1(n2519), .CO(n53211));
    SB_LUT4 add_2758_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n53209), 
            .O(n8194[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_21 (.CI(n52678), .I0(n294[19]), .I1(VCC_net), 
            .CO(n52679));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n52677), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_15 (.CI(n53209), .I0(n2600), .I1(n2397), .CO(n53210));
    SB_LUT4 add_2758_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n53208), 
            .O(n8194[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_14 (.CI(n53208), .I0(n2601), .I1(n2272), .CO(n53209));
    SB_LUT4 add_2758_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n53207), 
            .O(n8194[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_13 (.CI(n53207), .I0(n2602), .I1(n2144), .CO(n53208));
    SB_LUT4 i50919_3_lut (.I0(n34_adj_5058), .I1(baudrate[5]), .I2(n41_adj_5061), 
            .I3(GND_net), .O(n70189));   // verilog/uart_rx.v(119[33:55])
    defparam i50919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51814_2_lut_4_lut (.I0(n70761), .I1(baudrate[17]), .I2(n2596), 
            .I3(n27736), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i51814_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8220[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50920_3_lut (.I0(n70189), .I1(baudrate[6]), .I2(n43_adj_5062), 
            .I3(GND_net), .O(n70190));   // verilog/uart_rx.v(119[33:55])
    defparam i50920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50408_4_lut (.I0(n43_adj_5062), .I1(n41_adj_5061), .I2(n39_adj_5063), 
            .I3(n68773), .O(n69678));
    defparam i50408_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8220[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39_adj_5063), 
            .I3(GND_net), .O(n38_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n53206), 
            .O(n8194[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n52677), .I0(n294[18]), .I1(VCC_net), 
            .CO(n52678));
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8012[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_19_lut (.I0(n63101), .I1(n294[17]), .I2(VCC_net), 
            .I3(n52676), .O(n63103)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2758_12 (.CI(n53206), .I0(n2603), .I1(n2013), .CO(n53207));
    SB_CARRY sub_38_add_2_19 (.CI(n52676), .I0(n294[17]), .I1(VCC_net), 
            .CO(n52677));
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8220[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2758_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n53205), 
            .O(n8194[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_11 (.CI(n53205), .I0(n2604), .I1(n1879), .CO(n53206));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n63099), .I1(n294[16]), .I2(VCC_net), 
            .I3(n52675), .O(n63101)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_18 (.CI(n52675), .I0(n294[16]), .I1(VCC_net), 
            .CO(n52676));
    SB_LUT4 add_2758_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n53204), 
            .O(n8194[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_10 (.CI(n53204), .I0(n2605), .I1(n1742), .CO(n53205));
    SB_LUT4 add_2758_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n53203), 
            .O(n8194[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n63049), .I1(n294[15]), .I2(VCC_net), 
            .I3(n52674), .O(n63051)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2758_9 (.CI(n53203), .I0(n2606), .I1(n1602), .CO(n53204));
    SB_LUT4 add_2758_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n53202), 
            .O(n8194[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_8 (.CI(n53202), .I0(n2607), .I1(n1459), .CO(n53203));
    SB_LUT4 add_2758_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n53201), 
            .O(n8194[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_17 (.CI(n52674), .I0(n294[15]), .I1(VCC_net), 
            .CO(n52675));
    SB_LUT4 i49846_3_lut (.I0(n70190), .I1(baudrate[7]), .I2(n45_adj_5068), 
            .I3(GND_net), .O(n69116));   // verilog/uart_rx.v(119[33:55])
    defparam i49846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n63097), .I1(n294[14]), .I2(VCC_net), 
            .I3(n52673), .O(n63099)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8038[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2758_7 (.CI(n53201), .I0(n2608), .I1(n1460), .CO(n53202));
    SB_LUT4 add_2758_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n53200), 
            .O(n8194[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_6 (.CI(n53200), .I0(n2609), .I1(n1011), .CO(n53201));
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8220[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n53199), 
            .O(n8194[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_5 (.CI(n53199), .I0(n2610), .I1(n856), .CO(n53200));
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8220[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n53198), 
            .O(n8194[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_16 (.CI(n52673), .I0(n294[14]), .I1(VCC_net), 
            .CO(n52674));
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8064[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n52672), .O(n63097)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2758_4 (.CI(n53198), .I0(n2611), .I1(n698), .CO(n53199));
    SB_LUT4 add_2758_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n53197), 
            .O(n8194[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_3 (.CI(n53197), .I0(n2612), .I1(n858), .CO(n53198));
    SB_LUT4 i1_2_lut_adj_1002 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n63847));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'heeee;
    SB_LUT4 add_2758_2_lut (.I0(n61134), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2758_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53197));
    SB_LUT4 add_2757_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n53196), 
            .O(n8168[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n52672), .I0(n294[13]), .I1(VCC_net), 
            .CO(n52673));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n52671), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_14 (.CI(n52671), .I0(n294[12]), .I1(VCC_net), 
            .CO(n52672));
    SB_LUT4 i1_2_lut_adj_1003 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n63845));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8090[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2757_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n53195), 
            .O(n8168[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_17 (.CI(n53195), .I0(n2477), .I1(n2638), .CO(n53196));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n52670), .O(n63049)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n52670), .I0(n294[11]), .I1(VCC_net), 
            .CO(n52671));
    SB_LUT4 add_2757_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n53194), 
            .O(n8168[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_16 (.CI(n53194), .I0(n2478), .I1(n2519), .CO(n53195));
    SB_LUT4 add_2757_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n53193), 
            .O(n8168[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8116[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n52669), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8142[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2757_15 (.CI(n53193), .I0(n2479), .I1(n2397), .CO(n53194));
    SB_LUT4 add_2757_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n53192), 
            .O(n8168[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50933_4_lut (.I0(n69116), .I1(n38_adj_5064), .I2(n45_adj_5068), 
            .I3(n69678), .O(n70203));   // verilog/uart_rx.v(119[33:55])
    defparam i50933_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2757_14 (.CI(n53192), .I0(n2480), .I1(n2272), .CO(n53193));
    SB_LUT4 add_2757_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n53191), 
            .O(n8168[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_13 (.CI(n53191), .I0(n2481), .I1(n2144), .CO(n53192));
    SB_CARRY sub_38_add_2_12 (.CI(n52669), .I0(n294[10]), .I1(VCC_net), 
            .CO(n52670));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n52668), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n53190), 
            .O(n8168[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23828_rep_4_2_lut (.I0(n7986[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61158));   // verilog/uart_rx.v(119[33:55])
    defparam i23828_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_38_add_2_11 (.CI(n52668), .I0(n294[9]), .I1(VCC_net), 
            .CO(n52669));
    SB_CARRY add_2757_12 (.CI(n53190), .I0(n2482), .I1(n2013), .CO(n53191));
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8168[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2757_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n53189), 
            .O(n8168[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_11 (.CI(n53189), .I0(n2483), .I1(n1879), .CO(n53190));
    SB_LUT4 add_2757_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n53188), 
            .O(n8168[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n52667), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n52667), .I0(n294[8]), .I1(VCC_net), 
            .CO(n52668));
    SB_CARRY add_2757_10 (.CI(n53188), .I0(n2484), .I1(n1742), .CO(n53189));
    SB_LUT4 add_2757_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n53187), 
            .O(n8168[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_9 (.CI(n53187), .I0(n2485), .I1(n1602), .CO(n53188));
    SB_LUT4 add_2757_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n53186), 
            .O(n8168[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n52666), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_8 (.CI(n53186), .I0(n2486), .I1(n1459), .CO(n53187));
    SB_LUT4 add_2757_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n53185), 
            .O(n8168[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_7 (.CI(n53185), .I0(n2487), .I1(n1460), .CO(n53186));
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8194[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2757_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n53184), 
            .O(n8168[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n52666), .I0(n294[7]), .I1(VCC_net), 
            .CO(n52667));
    SB_CARRY add_2757_6 (.CI(n53184), .I0(n2488), .I1(n1011), .CO(n53185));
    SB_LUT4 add_2757_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n53183), 
            .O(n8168[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n52665), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_5 (.CI(n53183), .I0(n2489), .I1(n856), .CO(n53184));
    SB_LUT4 add_2757_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n53182), 
            .O(n8168[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_4 (.CI(n53182), .I0(n2490), .I1(n698), .CO(n53183));
    SB_LUT4 add_2757_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n53181), 
            .O(n8168[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_3 (.CI(n53181), .I0(n2491), .I1(n858), .CO(n53182));
    SB_CARRY sub_38_add_2_8 (.CI(n52665), .I0(n294[6]), .I1(VCC_net), 
            .CO(n52666));
    SB_LUT4 add_2757_2_lut (.I0(n61138), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2757_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53181));
    SB_LUT4 add_2756_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n53180), 
            .O(n8142[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2756_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n53179), 
            .O(n8142[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n52664), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_16 (.CI(n53179), .I0(n2354), .I1(n2519), .CO(n53180));
    SB_LUT4 add_2756_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n53178), 
            .O(n8142[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_15 (.CI(n53178), .I0(n2355), .I1(n2397), .CO(n53179));
    SB_CARRY sub_38_add_2_7 (.CI(n52664), .I0(n294[5]), .I1(VCC_net), 
            .CO(n52665));
    SB_LUT4 add_2756_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n53177), 
            .O(n8142[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_14 (.CI(n53177), .I0(n2356), .I1(n2272), .CO(n53178));
    SB_LUT4 add_2756_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n53176), 
            .O(n8142[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_13 (.CI(n53176), .I0(n2357), .I1(n2144), .CO(n53177));
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6261_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n23867));   // verilog/uart_rx.v(119[33:55])
    defparam i6261_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i49415_4_lut (.I0(n27648), .I1(n68022), .I2(n48_adj_5072), 
            .I3(baudrate[0]), .O(n804));
    defparam i49415_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 add_2756_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n53175), 
            .O(n8142[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n61158), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2756_12 (.CI(n53175), .I0(n2358), .I1(n2013), .CO(n53176));
    SB_LUT4 i50911_3_lut (.I0(n32_adj_5073), .I1(baudrate[6]), .I2(n39_adj_5074), 
            .I3(GND_net), .O(n70181));   // verilog/uart_rx.v(119[33:55])
    defparam i50911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50912_3_lut (.I0(n70181), .I1(baudrate[7]), .I2(n41_adj_5075), 
            .I3(GND_net), .O(n70182));   // verilog/uart_rx.v(119[33:55])
    defparam i50912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50384_4_lut (.I0(n41_adj_5075), .I1(n39_adj_5074), .I2(n37_adj_5076), 
            .I3(n68730), .O(n69654));
    defparam i50384_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50937_3_lut (.I0(n34_adj_5077), .I1(baudrate[5]), .I2(n37_adj_5076), 
            .I3(GND_net), .O(n70207));   // verilog/uart_rx.v(119[33:55])
    defparam i50937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8246[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2756_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n53174), 
            .O(n8142[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49851_3_lut (.I0(n70182), .I1(baudrate[8]), .I2(n43_adj_5078), 
            .I3(GND_net), .O(n69121));   // verilog/uart_rx.v(119[33:55])
    defparam i49851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51213_4_lut (.I0(n69121), .I1(n70207), .I2(n43_adj_5078), 
            .I3(n69654), .O(n70483));   // verilog/uart_rx.v(119[33:55])
    defparam i51213_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51214_3_lut (.I0(n70483), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n70484));   // verilog/uart_rx.v(119[33:55])
    defparam i51214_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8220[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n70484), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8246[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(n63889), .I1(n63845), .I2(n63847), 
            .I3(baudrate[11]), .O(n63875));
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1005 (.I0(n63875), .I1(n63877), .I2(n63865), 
            .I3(n63821), .O(n27715));
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n27715), .I1(n48_adj_5079), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8038[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8064[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8246[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8090[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8116[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8142[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8168[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8194[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8220[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n52663), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_11 (.CI(n53174), .I0(n2359), .I1(n1879), .CO(n53175));
    SB_LUT4 add_2756_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n53173), 
            .O(n8142[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_10 (.CI(n53173), .I0(n2360), .I1(n1742), .CO(n53174));
    SB_LUT4 add_2756_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n53172), 
            .O(n8142[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_9 (.CI(n53172), .I0(n2361), .I1(n1602), .CO(n53173));
    SB_LUT4 add_2756_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n53171), 
            .O(n8142[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_8 (.CI(n53171), .I0(n2362), .I1(n1459), .CO(n53172));
    SB_LUT4 add_2756_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n53170), 
            .O(n8142[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7986[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8012[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_7 (.CI(n53170), .I0(n2363), .I1(n1460), .CO(n53171));
    SB_LUT4 add_2756_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n53169), 
            .O(n8142[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_6 (.CI(n53169), .I0(n2364), .I1(n1011), .CO(n53170));
    SB_LUT4 add_2756_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n53168), 
            .O(n8142[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8038[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8064[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8090[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8116[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_5 (.CI(n53168), .I0(n2365), .I1(n856), .CO(n53169));
    SB_LUT4 add_2756_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n53167), 
            .O(n8142[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8142[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(n63903), .I1(n63009), .I2(n63007), 
            .I3(n63893), .O(n27736));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_CARRY add_2756_4 (.CI(n53167), .I0(n2366), .I1(n698), .CO(n53168));
    SB_LUT4 add_2756_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n53166), 
            .O(n8142[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_3 (.CI(n53166), .I0(n2367), .I1(n858), .CO(n53167));
    SB_LUT4 add_2756_2_lut (.I0(n61142), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2756_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53166));
    SB_CARRY sub_38_add_2_6 (.CI(n52663), .I0(n294[4]), .I1(VCC_net), 
            .CO(n52664));
    SB_LUT4 add_2755_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n53165), 
            .O(n8116[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2755_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n53164), 
            .O(n8116[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_15 (.CI(n53164), .I0(n2228), .I1(n2397), .CO(n53165));
    SB_LUT4 add_2755_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n53163), 
            .O(n8116[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_14 (.CI(n53163), .I0(n2229), .I1(n2272), .CO(n53164));
    SB_LUT4 i49223_4_lut (.I0(n23_adj_5082), .I1(n21_adj_5083), .I2(n19_adj_5084), 
            .I3(n17_adj_5081), .O(n68493));
    defparam i49223_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49210_4_lut (.I0(n29_adj_5085), .I1(n27_adj_5086), .I2(n25_adj_5087), 
            .I3(n68493), .O(n68480));
    defparam i49210_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51064_4_lut (.I0(n35_adj_5088), .I1(n33_adj_5089), .I2(n31_adj_5090), 
            .I3(n68480), .O(n70334));
    defparam i51064_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2755_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n53162), 
            .O(n8116[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_13 (.CI(n53162), .I0(n2230), .I1(n2144), .CO(n53163));
    SB_LUT4 add_2755_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n53161), 
            .O(n8116[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n52662), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_12 (.CI(n53161), .I0(n2231), .I1(n2013), .CO(n53162));
    SB_LUT4 add_2755_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n53160), 
            .O(n8116[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_11 (.CI(n53160), .I0(n2232), .I1(n1879), .CO(n53161));
    SB_LUT4 add_2755_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n53159), 
            .O(n8116[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_10 (.CI(n53159), .I0(n2233), .I1(n1742), .CO(n53160));
    SB_LUT4 add_2755_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n53158), 
            .O(n8116[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_9 (.CI(n53158), .I0(n2234), .I1(n1602), .CO(n53159));
    SB_LUT4 add_2755_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n53157), 
            .O(n8116[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_8 (.CI(n53157), .I0(n2235), .I1(n1459), .CO(n53158));
    SB_LUT4 add_2755_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n53156), 
            .O(n8116[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8064[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2755_7 (.CI(n53156), .I0(n2236), .I1(n1460), .CO(n53157));
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5092), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 add_2755_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n53155), 
            .O(n8116[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_6 (.CI(n53155), .I0(n2237), .I1(n1011), .CO(n53156));
    SB_LUT4 add_2755_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n53154), 
            .O(n8116[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8090[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2755_5 (.CI(n53154), .I0(n2238), .I1(n856), .CO(n53155));
    SB_LUT4 add_2755_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n53153), 
            .O(n8116[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_4 (.CI(n53153), .I0(n2239), .I1(n698), .CO(n53154));
    SB_LUT4 add_2755_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n53152), 
            .O(n8116[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_3 (.CI(n53152), .I0(n2240), .I1(n858), .CO(n53153));
    SB_LUT4 add_2755_2_lut (.I0(n61146), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8220[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2755_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53152));
    SB_LUT4 add_2754_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n53151), 
            .O(n8090[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n53150), 
            .O(n8090[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8246[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_13 (.CI(n53150), .I0(n2099), .I1(n2272), .CO(n53151));
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8246[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5094), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8246[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n53149), 
            .O(n8090[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_12 (.CI(n53149), .I0(n2100), .I1(n2144), .CO(n53150));
    SB_LUT4 add_2754_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n53148), 
            .O(n8090[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8116[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_11 (.CI(n53148), .I0(n2101), .I1(n2013), .CO(n53149));
    SB_LUT4 add_2754_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n53147), 
            .O(n8090[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8246[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8246[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7908[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8246[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_10 (.CI(n53147), .I0(n2102), .I1(n1879), .CO(n53148));
    SB_LUT4 add_2754_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n53146), 
            .O(n8090[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_9 (.CI(n53146), .I0(n2103), .I1(n1742), .CO(n53147));
    SB_LUT4 add_2754_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n53145), 
            .O(n8090[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8246[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8246[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_8 (.CI(n53145), .I0(n2104), .I1(n1602), .CO(n53146));
    SB_LUT4 add_2754_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n53144), 
            .O(n8090[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_7 (.CI(n53144), .I0(n2105), .I1(n1459), .CO(n53145));
    SB_CARRY sub_38_add_2_5 (.CI(n52662), .I0(n294[3]), .I1(VCC_net), 
            .CO(n52663));
    SB_LUT4 add_2754_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n53143), 
            .O(n8090[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n52661), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8246[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8246[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7934[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50881_3_lut (.I0(n16_adj_5091), .I1(baudrate[13]), .I2(n39_adj_5104), 
            .I3(GND_net), .O(n70151));   // verilog/uart_rx.v(119[33:55])
    defparam i50881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_6 (.CI(n53143), .I0(n2106), .I1(n1460), .CO(n53144));
    SB_CARRY sub_38_add_2_4 (.CI(n52661), .I0(n294[2]), .I1(VCC_net), 
            .CO(n52662));
    SB_LUT4 add_2754_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n53142), 
            .O(n8090[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_5 (.CI(n53142), .I0(n2107), .I1(n1011), .CO(n53143));
    SB_LUT4 add_2754_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n53141), 
            .O(n8090[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_4 (.CI(n53141), .I0(n2108), .I1(n856), .CO(n53142));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n52660), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8246[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8246[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7960[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49063_4_lut (.I0(n35_adj_5107), .I1(n23_adj_5108), .I2(n21_adj_5109), 
            .I3(n19_adj_5110), .O(n68333));
    defparam i49063_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7986[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8246[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_3 (.CI(n52660), .I0(n294[1]), .I1(VCC_net), 
            .CO(n52661));
    SB_LUT4 add_2754_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n53140), 
            .O(n8090[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_3 (.CI(n53140), .I0(n2109), .I1(n698), .CO(n53141));
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8090[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n53140));
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8246[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2753_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n53139), 
            .O(n8064[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n53138), 
            .O(n8064[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2753_13 (.CI(n53138), .I0(n1967), .I1(n2144), .CO(n53139));
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8012[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n53137), 
            .O(n8064[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_12 (.CI(n53137), .I0(n1968), .I1(n2013), .CO(n53138));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n61968), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49002_4_lut (.I0(n33_adj_5117), .I1(n21_adj_5121), .I2(n19_adj_5120), 
            .I3(n17_adj_5118), .O(n68272));
    defparam i49002_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2753_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n53136), 
            .O(n8064[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_11 (.CI(n53136), .I0(n1969), .I1(n1879), .CO(n53137));
    SB_LUT4 add_2753_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n53135), 
            .O(n8064[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50047_4_lut (.I0(n15_adj_5116), .I1(n13_adj_5115), .I2(n2956), 
            .I3(baudrate[2]), .O(n69317));
    defparam i50047_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50656_4_lut (.I0(n21_adj_5121), .I1(n19_adj_5120), .I2(n17_adj_5118), 
            .I3(n69317), .O(n69926));
    defparam i50656_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2753_10 (.CI(n53135), .I0(n1970), .I1(n1742), .CO(n53136));
    SB_LUT4 add_2753_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n53134), 
            .O(n8064[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50652_4_lut (.I0(n27_adj_5114), .I1(n25_adj_5113), .I2(n23_adj_5111), 
            .I3(n69926), .O(n69922));
    defparam i50652_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n61968), .I1(GND_net), 
            .CO(n52660));
    SB_LUT4 i49006_4_lut (.I0(n33_adj_5117), .I1(n31_adj_5105), .I2(n29_adj_5103), 
            .I3(n69922), .O(n68276));
    defparam i49006_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2753_9 (.CI(n53134), .I0(n1971), .I1(n1602), .CO(n53135));
    SB_LUT4 add_2753_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n53133), 
            .O(n8064[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_8 (.CI(n53133), .I0(n1972), .I1(n1459), .CO(n53134));
    SB_LUT4 add_2753_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n53132), 
            .O(n8064[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_7 (.CI(n53132), .I0(n1973), .I1(n1460), .CO(n53133));
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50105_4_lut (.I0(n17_adj_5124), .I1(n15_adj_5096), .I2(n2844), 
            .I3(baudrate[2]), .O(n69375));
    defparam i50105_4_lut.LUT_INIT = 16'heffe;
    SB_DFFESR r_Clock_Count_2054__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n29942), .D(n1[0]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i50882_3_lut (.I0(n70151), .I1(baudrate[14]), .I2(n41_adj_5126), 
            .I3(GND_net), .O(n70152));   // verilog/uart_rx.v(119[33:55])
    defparam i50882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50851_3_lut (.I0(n10_adj_5123), .I1(baudrate[13]), .I2(n33_adj_5117), 
            .I3(GND_net), .O(n70121));   // verilog/uart_rx.v(119[33:55])
    defparam i50851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50852_3_lut (.I0(n70121), .I1(baudrate[14]), .I2(n35_adj_5100), 
            .I3(GND_net), .O(n70122));   // verilog/uart_rx.v(119[33:55])
    defparam i50852_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n31702));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8038[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n71701));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5127), .I1(baudrate[17]), 
            .I2(n41_adj_5097), .I3(GND_net), .O(n36_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48992_4_lut (.I0(n39_adj_5101), .I1(n37_adj_5099), .I2(n35_adj_5100), 
            .I3(n68272), .O(n68262));
    defparam i48992_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2753_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n53131), 
            .O(n8064[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_5129), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2753_6 (.CI(n53131), .I0(n1974), .I1(n1011), .CO(n53132));
    SB_LUT4 add_2753_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n53130), 
            .O(n8064[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_5 (.CI(n53130), .I0(n1975), .I1(n856), .CO(n53131));
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8064[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2753_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n53129), 
            .O(n8064[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_4 (.CI(n53129), .I0(n1976), .I1(n698), .CO(n53130));
    SB_LUT4 add_2753_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n53128), 
            .O(n8064[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_3 (.CI(n53128), .I0(n1977), .I1(n858), .CO(n53129));
    SB_LUT4 i50179_4_lut (.I0(n41_adj_5126), .I1(n39_adj_5104), .I2(n27_adj_5086), 
            .I3(n68489), .O(n69449));
    defparam i50179_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2753_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8064[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53128));
    SB_LUT4 add_2752_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n53127), 
            .O(n8038[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51379_4_lut (.I0(n36_adj_5128), .I1(n16_adj_5130), .I2(n41_adj_5097), 
            .I3(n68258), .O(n70649));   // verilog/uart_rx.v(119[33:55])
    defparam i51379_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2752_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n53126), 
            .O(n8038[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49920_3_lut (.I0(n70122), .I1(baudrate[15]), .I2(n37_adj_5099), 
            .I3(GND_net), .O(n69190));   // verilog/uart_rx.v(119[33:55])
    defparam i49920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50680_4_lut (.I0(n23_adj_5108), .I1(n21_adj_5109), .I2(n19_adj_5110), 
            .I3(n69375), .O(n69950));
    defparam i50680_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50674_4_lut (.I0(n29_adj_5093), .I1(n27_adj_5080), .I2(n25_adj_5133), 
            .I3(n69950), .O(n69944));
    defparam i50674_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2752_12 (.CI(n53126), .I0(n1832), .I1(n2013), .CO(n53127));
    SB_LUT4 i50950_3_lut (.I0(n22_adj_5135), .I1(baudrate[7]), .I2(n27_adj_5086), 
            .I3(GND_net), .O(n70220));   // verilog/uart_rx.v(119[33:55])
    defparam i50950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49898_3_lut (.I0(n70152), .I1(baudrate[15]), .I2(n43_adj_5136), 
            .I3(GND_net), .O(n69168));   // verilog/uart_rx.v(119[33:55])
    defparam i49898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n53125), 
            .O(n8038[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8090[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_11 (.CI(n53125), .I0(n1833), .I1(n1879), .CO(n53126));
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5137), .I1(baudrate[9]), 
            .I2(n31_adj_5090), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51365_4_lut (.I0(n28), .I1(n18_adj_5138), .I2(n31_adj_5090), 
            .I3(n68476), .O(n70635));   // verilog/uart_rx.v(119[33:55])
    defparam i51365_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51366_3_lut (.I0(n70635), .I1(baudrate[10]), .I2(n33_adj_5089), 
            .I3(GND_net), .O(n70636));   // verilog/uart_rx.v(119[33:55])
    defparam i51366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51194_3_lut (.I0(n70636), .I1(baudrate[11]), .I2(n35_adj_5088), 
            .I3(GND_net), .O(n70464));   // verilog/uart_rx.v(119[33:55])
    defparam i51194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50185_4_lut (.I0(n41_adj_5126), .I1(n39_adj_5104), .I2(n37_adj_5139), 
            .I3(n70334), .O(n69455));
    defparam i50185_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2752_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n53124), 
            .O(n8038[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51191_4_lut (.I0(n69168), .I1(n70220), .I2(n43_adj_5136), 
            .I3(n69449), .O(n70461));   // verilog/uart_rx.v(119[33:55])
    defparam i51191_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49896_3_lut (.I0(n70464), .I1(baudrate[12]), .I2(n37_adj_5139), 
            .I3(GND_net), .O(n69166));   // verilog/uart_rx.v(119[33:55])
    defparam i49896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51490_4_lut (.I0(n69166), .I1(n70461), .I2(n43_adj_5136), 
            .I3(n69455), .O(n70760));   // verilog/uart_rx.v(119[33:55])
    defparam i51490_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51491_3_lut (.I0(n70760), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n70761));   // verilog/uart_rx.v(119[33:55])
    defparam i51491_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8168[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8194[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8116[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(n63889), .I1(n63797), .I2(n63601), 
            .I3(baudrate[19]), .O(n63621));
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5142), .I1(baudrate[9]), 
            .I2(n25_adj_5113), .I3(GND_net), .O(n22_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51377_4_lut (.I0(n22_adj_5143), .I1(n12_adj_5144), .I2(n25_adj_5113), 
            .I3(n68292), .O(n70647));   // verilog/uart_rx.v(119[33:55])
    defparam i51377_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49065_4_lut (.I0(n35_adj_5107), .I1(n33_adj_5056), .I2(n31_adj_5069), 
            .I3(n69944), .O(n68335));
    defparam i49065_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2752_10 (.CI(n53124), .I0(n1834), .I1(n1742), .CO(n53125));
    SB_LUT4 i51378_3_lut (.I0(n70647), .I1(baudrate[10]), .I2(n27_adj_5114), 
            .I3(GND_net), .O(n70648));   // verilog/uart_rx.v(119[33:55])
    defparam i51378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51164_3_lut (.I0(n70648), .I1(baudrate[11]), .I2(n29_adj_5103), 
            .I3(GND_net), .O(n70434));   // verilog/uart_rx.v(119[33:55])
    defparam i51164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n53123), 
            .O(n8038[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(n63621), .I1(n63849), .I2(n63891), 
            .I3(n63847), .O(n27739));
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'hfffe;
    SB_LUT4 i49127_4_lut (.I0(n37_adj_5145), .I1(n25_adj_5146), .I2(n23_adj_5147), 
            .I3(n21_adj_5148), .O(n68397));
    defparam i49127_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2752_9 (.CI(n53123), .I0(n1835), .I1(n1602), .CO(n53124));
    SB_LUT4 add_2752_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n53122), 
            .O(n8038[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50161_4_lut (.I0(n19_adj_5149), .I1(n17_adj_5150), .I2(n2729), 
            .I3(baudrate[2]), .O(n69431));
    defparam i50161_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50708_4_lut (.I0(n25_adj_5146), .I1(n23_adj_5147), .I2(n21_adj_5148), 
            .I3(n69431), .O(n69978));
    defparam i50708_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50702_4_lut (.I0(n31_adj_5140), .I1(n29_adj_5141), .I2(n27_adj_5151), 
            .I3(n69978), .O(n69972));
    defparam i50702_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49129_4_lut (.I0(n37_adj_5145), .I1(n35_adj_5071), .I2(n33_adj_5030), 
            .I3(n69972), .O(n68399));
    defparam i49129_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50875_3_lut (.I0(n14_adj_5152), .I1(baudrate[13]), .I2(n37_adj_5145), 
            .I3(GND_net), .O(n70145));   // verilog/uart_rx.v(119[33:55])
    defparam i50875_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_8 (.CI(n53122), .I0(n1836), .I1(n1459), .CO(n53123));
    SB_LUT4 add_2752_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n53121), 
            .O(n8038[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_7 (.CI(n53121), .I0(n1837), .I1(n1460), .CO(n53122));
    SB_LUT4 add_2752_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n53120), 
            .O(n8038[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51022_4_lut (.I0(n39_adj_5101), .I1(n37_adj_5099), .I2(n35_adj_5100), 
            .I3(n68276), .O(n70292));
    defparam i51022_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2752_6 (.CI(n53120), .I0(n1838), .I1(n1011), .CO(n53121));
    SB_LUT4 add_2752_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n53119), 
            .O(n8038[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_5 (.CI(n53119), .I0(n1839), .I1(n856), .CO(n53120));
    SB_LUT4 add_2752_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n53118), 
            .O(n8038[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_4 (.CI(n53118), .I0(n1840), .I1(n698), .CO(n53119));
    SB_LUT4 add_2752_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n53117), 
            .O(n8038[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51563_4_lut (.I0(n69190), .I1(n70649), .I2(n41_adj_5097), 
            .I3(n68262), .O(n70833));   // verilog/uart_rx.v(119[33:55])
    defparam i51563_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49918_3_lut (.I0(n70434), .I1(baudrate[12]), .I2(n31_adj_5105), 
            .I3(GND_net), .O(n69188));   // verilog/uart_rx.v(119[33:55])
    defparam i49918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Clock_Count_2054__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n29942), .D(n1[7]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n29942), .D(n1[6]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n29942), .D(n1[5]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n29942), .D(n1[4]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n29942), .D(n1[3]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n29942), .D(n1[2]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2054__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n29942), .D(n1[1]), .R(n31162));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8142[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_3 (.CI(n53117), .I0(n1841), .I1(n858), .CO(n53118));
    SB_LUT4 add_2752_2_lut (.I0(n61155), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2752_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53117));
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51623_4_lut (.I0(n69188), .I1(n70833), .I2(n41_adj_5097), 
            .I3(n70292), .O(n70893));   // verilog/uart_rx.v(119[33:55])
    defparam i51623_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51624_3_lut (.I0(n70893), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n70894));   // verilog/uart_rx.v(119[33:55])
    defparam i51624_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50871_3_lut (.I0(n12_adj_5162), .I1(baudrate[13]), .I2(n35_adj_5107), 
            .I3(GND_net), .O(n70141));   // verilog/uart_rx.v(119[33:55])
    defparam i50871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8168[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2054_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n53467), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51622_3_lut (.I0(n70894), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n70892));   // verilog/uart_rx.v(119[33:55])
    defparam i51622_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50876_3_lut (.I0(n70145), .I1(baudrate[14]), .I2(n39_adj_5167), 
            .I3(GND_net), .O(n70146));   // verilog/uart_rx.v(119[33:55])
    defparam i50876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5168), .I1(baudrate[17]), 
            .I2(n45_adj_5169), .I3(GND_net), .O(n40_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49117_4_lut (.I0(n43_adj_5171), .I1(n41_adj_5172), .I2(n39_adj_5167), 
            .I3(n68397), .O(n68387));
    defparam i49117_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50952_4_lut (.I0(n40_adj_5170), .I1(n20_adj_5173), .I2(n45_adj_5169), 
            .I3(n68381), .O(n70222));   // verilog/uart_rx.v(119[33:55])
    defparam i50952_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49908_3_lut (.I0(n70146), .I1(baudrate[15]), .I2(n41_adj_5172), 
            .I3(GND_net), .O(n69178));   // verilog/uart_rx.v(119[33:55])
    defparam i49908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5174), .I1(baudrate[9]), 
            .I2(n29_adj_5141), .I3(GND_net), .O(n26_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49437_4_lut (.I0(n35_adj_5166), .I1(n33_adj_5165), .I2(n31_adj_5164), 
            .I3(n29_adj_5176), .O(n68707));
    defparam i49437_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 r_Clock_Count_2054_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n53466), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_8 (.CI(n53466), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n53467));
    SB_LUT4 r_Clock_Count_2054_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n53465), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_7 (.CI(n53465), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n53466));
    SB_LUT4 r_Clock_Count_2054_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n53464), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_6 (.CI(n53464), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n53465));
    SB_LUT4 r_Clock_Count_2054_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n53463), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_5 (.CI(n53463), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n53464));
    SB_LUT4 r_Clock_Count_2054_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n53462), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_4 (.CI(n53462), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n53463));
    SB_LUT4 r_Clock_Count_2054_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n53461), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_3 (.CI(n53461), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n53462));
    SB_LUT4 i51367_4_lut (.I0(n26_adj_5175), .I1(n16_adj_5177), .I2(n29_adj_5141), 
            .I3(n68415), .O(n70637));   // verilog/uart_rx.v(119[33:55])
    defparam i51367_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 r_Clock_Count_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n53461));
    SB_LUT4 i45268_2_lut (.I0(baudrate[8]), .I1(n64527), .I2(GND_net), 
            .I3(GND_net), .O(n64529));
    defparam i45268_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2751_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n53106), 
            .O(n8012[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2751_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n53105), 
            .O(n8012[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_10 (.CI(n53105), .I0(n1694), .I1(n1879), .CO(n53106));
    SB_LUT4 add_2751_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n53104), 
            .O(n8012[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_9 (.CI(n53104), .I0(n1695), .I1(n1742), .CO(n53105));
    SB_LUT4 add_2751_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n53103), 
            .O(n8012[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_8 (.CI(n53103), .I0(n1696), .I1(n1602), .CO(n53104));
    SB_LUT4 i1_2_lut_adj_1009 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n63635));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5178), .I1(baudrate[17]), 
            .I2(n43_adj_5070), .I3(GND_net), .O(n38_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5180), .I1(baudrate[9]), 
            .I2(n43_adj_5154), .I3(GND_net), .O(n40_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2751_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n53102), 
            .O(n8012[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_7 (.CI(n53102), .I0(n1697), .I1(n1459), .CO(n53103));
    SB_LUT4 i50872_3_lut (.I0(n70141), .I1(baudrate[14]), .I2(n37_adj_5065), 
            .I3(GND_net), .O(n70142));   // verilog/uart_rx.v(119[33:55])
    defparam i50872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50907_3_lut (.I0(n28_adj_5182), .I1(baudrate[5]), .I2(n35_adj_5166), 
            .I3(GND_net), .O(n70177));   // verilog/uart_rx.v(119[33:55])
    defparam i50907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50908_3_lut (.I0(n70177), .I1(baudrate[6]), .I2(n37_adj_5134), 
            .I3(GND_net), .O(n70178));   // verilog/uart_rx.v(119[33:55])
    defparam i50908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n53101), 
            .O(n8012[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_6 (.CI(n53101), .I0(n1698), .I1(n1460), .CO(n53102));
    SB_LUT4 i49416_4_lut (.I0(n41_adj_5163), .I1(n39_adj_5153), .I2(n37_adj_5134), 
            .I3(n68707), .O(n68686));
    defparam i49416_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2751_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n53100), 
            .O(n8012[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_5 (.CI(n53100), .I0(n1699), .I1(n1011), .CO(n53101));
    SB_LUT4 add_2751_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n53099), 
            .O(n8012[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49053_4_lut (.I0(n41_adj_5067), .I1(n39_adj_5066), .I2(n37_adj_5065), 
            .I3(n68333), .O(n68323));
    defparam i49053_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51343_4_lut (.I0(n40_adj_5181), .I1(n30_adj_5183), .I2(n43_adj_5154), 
            .I3(n68683), .O(n70613));   // verilog/uart_rx.v(119[33:55])
    defparam i51343_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51337_4_lut (.I0(n38_adj_5179), .I1(n18_adj_5184), .I2(n43_adj_5070), 
            .I3(n68321), .O(n70607));   // verilog/uart_rx.v(119[33:55])
    defparam i51337_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49854_3_lut (.I0(n70178), .I1(baudrate[7]), .I2(n39_adj_5153), 
            .I3(GND_net), .O(n69124));   // verilog/uart_rx.v(119[33:55])
    defparam i49854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51551_4_lut (.I0(n69124), .I1(n70613), .I2(n43_adj_5154), 
            .I3(n68686), .O(n70821));   // verilog/uart_rx.v(119[33:55])
    defparam i51551_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2751_4 (.CI(n53099), .I0(n1700), .I1(n856), .CO(n53100));
    SB_LUT4 i51552_3_lut (.I0(n70821), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n70822));   // verilog/uart_rx.v(119[33:55])
    defparam i51552_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49914_3_lut (.I0(n70142), .I1(baudrate[15]), .I2(n39_adj_5066), 
            .I3(GND_net), .O(n69184));   // verilog/uart_rx.v(119[33:55])
    defparam i49914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n53098), 
            .O(n8012[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_3 (.CI(n53098), .I0(n1701), .I1(n698), .CO(n53099));
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5188), .I1(baudrate[9]), 
            .I2(n27_adj_5080), .I3(GND_net), .O(n24_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51369_4_lut (.I0(n24_adj_5189), .I1(n14_adj_5191), .I2(n27_adj_5080), 
            .I3(n68349), .O(n70639));   // verilog/uart_rx.v(119[33:55])
    defparam i51369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8012[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51370_3_lut (.I0(n70639), .I1(baudrate[10]), .I2(n29_adj_5093), 
            .I3(GND_net), .O(n70640));   // verilog/uart_rx.v(119[33:55])
    defparam i51370_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n29821), 
            .D(n479[1]), .R(n31149));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i51186_3_lut (.I0(n70640), .I1(baudrate[11]), .I2(n31_adj_5069), 
            .I3(GND_net), .O(n70456));   // verilog/uart_rx.v(119[33:55])
    defparam i51186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51040_4_lut (.I0(n41_adj_5067), .I1(n39_adj_5066), .I2(n37_adj_5065), 
            .I3(n68335), .O(n70310));
    defparam i51040_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49400_4_lut (.I0(n33_adj_5192), .I1(n31_adj_5190), .I2(n29_adj_5187), 
            .I3(n27_adj_5193), .O(n68670));
    defparam i49400_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51549_4_lut (.I0(n69184), .I1(n70607), .I2(n43_adj_5070), 
            .I3(n68323), .O(n70819));   // verilog/uart_rx.v(119[33:55])
    defparam i51549_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2751_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n53098));
    SB_LUT4 i49912_3_lut (.I0(n70456), .I1(baudrate[12]), .I2(n33_adj_5056), 
            .I3(GND_net), .O(n69182));   // verilog/uart_rx.v(119[33:55])
    defparam i49912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5194), .I1(baudrate[9]), 
            .I2(n41_adj_5185), .I3(GND_net), .O(n38_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51611_4_lut (.I0(n69182), .I1(n70819), .I2(n43_adj_5070), 
            .I3(n70310), .O(n70881));   // verilog/uart_rx.v(119[33:55])
    defparam i51611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51612_3_lut (.I0(n70881), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n70882));   // verilog/uart_rx.v(119[33:55])
    defparam i51612_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50905_3_lut (.I0(n26_adj_5196), .I1(baudrate[5]), .I2(n33_adj_5192), 
            .I3(GND_net), .O(n70175));   // verilog/uart_rx.v(119[33:55])
    defparam i50905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n53097), 
            .O(n7986[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2750_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n53096), 
            .O(n7986[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7986[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50906_3_lut (.I0(n70175), .I1(baudrate[6]), .I2(n35_adj_5132), 
            .I3(GND_net), .O(n70176));   // verilog/uart_rx.v(119[33:55])
    defparam i50906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49383_4_lut (.I0(n39_adj_5186), .I1(n37_adj_5131), .I2(n35_adj_5132), 
            .I3(n68670), .O(n68653));
    defparam i49383_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51355_4_lut (.I0(n38_adj_5195), .I1(n28_adj_5197), .I2(n41_adj_5185), 
            .I3(n68650), .O(n70625));   // verilog/uart_rx.v(119[33:55])
    defparam i51355_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49856_3_lut (.I0(n70176), .I1(baudrate[7]), .I2(n37_adj_5131), 
            .I3(GND_net), .O(n69126));   // verilog/uart_rx.v(119[33:55])
    defparam i49856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51555_4_lut (.I0(n69126), .I1(n70625), .I2(n41_adj_5185), 
            .I3(n68653), .O(n70825));   // verilog/uart_rx.v(119[33:55])
    defparam i51555_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51556_3_lut (.I0(n70825), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n70826));   // verilog/uart_rx.v(119[33:55])
    defparam i51556_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8012[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8038[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51497_3_lut (.I0(n70826), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n70767));   // verilog/uart_rx.v(119[33:55])
    defparam i51497_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49862_3_lut (.I0(n70767), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam i49862_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8090[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8064[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8090[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8116[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49291_4_lut (.I0(n27_adj_5204), .I1(n25_adj_5200), .I2(n23_adj_5199), 
            .I3(n21_adj_5205), .O(n68561));
    defparam i49291_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49286_4_lut (.I0(n33_adj_5122), .I1(n31_adj_5119), .I2(n29_adj_5112), 
            .I3(n68561), .O(n68556));
    defparam i49286_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51227_3_lut (.I0(n42_adj_5201), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n70497));   // verilog/uart_rx.v(119[33:55])
    defparam i51227_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49332_4_lut (.I0(n29_adj_5210), .I1(n27_adj_5211), .I2(n25_adj_5212), 
            .I3(n23_adj_5209), .O(n68602));
    defparam i49332_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5214), .I1(baudrate[7]), 
            .I2(n31_adj_5119), .I3(GND_net), .O(n28_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49324_4_lut (.I0(n35_adj_5216), .I1(n33_adj_5203), .I2(n31_adj_5217), 
            .I3(n68602), .O(n68594));
    defparam i49324_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2750_10 (.CI(n53096), .I0(n1553), .I1(n1742), .CO(n53097));
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5218), .I1(baudrate[9]), 
            .I2(n35_adj_5106), .I3(GND_net), .O(n32_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51361_4_lut (.I0(n32_adj_5219), .I1(n22_adj_5220), .I2(n35_adj_5106), 
            .I3(n68552), .O(n70631));   // verilog/uart_rx.v(119[33:55])
    defparam i51361_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51362_3_lut (.I0(n70631), .I1(baudrate[10]), .I2(n37_adj_5102), 
            .I3(GND_net), .O(n70632));   // verilog/uart_rx.v(119[33:55])
    defparam i51362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51202_3_lut (.I0(n70632), .I1(baudrate[11]), .I2(n39_adj_5098), 
            .I3(GND_net), .O(n70472));   // verilog/uart_rx.v(119[33:55])
    defparam i51202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51228_3_lut (.I0(n70497), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n70498));   // verilog/uart_rx.v(119[33:55])
    defparam i51228_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5222), .I1(baudrate[7]), 
            .I2(n33_adj_5203), .I3(GND_net), .O(n30_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51074_4_lut (.I0(n39_adj_5098), .I1(n37_adj_5102), .I2(n35_adj_5106), 
            .I3(n68556), .O(n70344));
    defparam i51074_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51456_4_lut (.I0(n28_adj_5215), .I1(n20_adj_5213), .I2(n31_adj_5119), 
            .I3(n68558), .O(n70726));   // verilog/uart_rx.v(119[33:55])
    defparam i51456_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49882_3_lut (.I0(n70472), .I1(baudrate[12]), .I2(n41_adj_5095), 
            .I3(GND_net), .O(n69152));   // verilog/uart_rx.v(119[33:55])
    defparam i49882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41903_1_lut (.I0(n27742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61126));
    defparam i41903_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51553_4_lut (.I0(n69152), .I1(n70726), .I2(n41_adj_5095), 
            .I3(n70344), .O(n70823));   // verilog/uart_rx.v(119[33:55])
    defparam i51553_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50928_3_lut (.I0(n70498), .I1(baudrate[4]), .I2(n60872), 
            .I3(GND_net), .O(n48_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam i50928_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i49412_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i49412_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7908[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51368_3_lut (.I0(n70637), .I1(baudrate[10]), .I2(n31_adj_5140), 
            .I3(GND_net), .O(n70638));   // verilog/uart_rx.v(119[33:55])
    defparam i51368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51190_3_lut (.I0(n70638), .I1(baudrate[11]), .I2(n33_adj_5030), 
            .I3(GND_net), .O(n70460));   // verilog/uart_rx.v(119[33:55])
    defparam i51190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51554_3_lut (.I0(n70823), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n70824));   // verilog/uart_rx.v(119[33:55])
    defparam i51554_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51499_3_lut (.I0(n70824), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n70769));   // verilog/uart_rx.v(119[33:55])
    defparam i51499_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2750_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n53095), 
            .O(n7986[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_9 (.CI(n53095), .I0(n1554), .I1(n1602), .CO(n53096));
    SB_LUT4 add_2750_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n53094), 
            .O(n7986[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51052_4_lut (.I0(n43_adj_5171), .I1(n41_adj_5172), .I2(n39_adj_5167), 
            .I3(n68399), .O(n70322));
    defparam i51052_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51431_4_lut (.I0(n69178), .I1(n70222), .I2(n45_adj_5169), 
            .I3(n68387), .O(n70701));   // verilog/uart_rx.v(119[33:55])
    defparam i51431_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7934[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7960[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49906_3_lut (.I0(n70460), .I1(baudrate[12]), .I2(n35_adj_5071), 
            .I3(GND_net), .O(n69176));   // verilog/uart_rx.v(119[33:55])
    defparam i49906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51433_4_lut (.I0(n69176), .I1(n70701), .I2(n45_adj_5169), 
            .I3(n70322), .O(n70703));   // verilog/uart_rx.v(119[33:55])
    defparam i51433_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n29821), 
            .D(n479[2]), .R(n31149));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7986[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2750_8 (.CI(n53094), .I0(n1555), .I1(n1459), .CO(n53095));
    SB_LUT4 add_2750_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n53093), 
            .O(n7986[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_7 (.CI(n53093), .I0(n1556), .I1(n1460), .CO(n53094));
    SB_LUT4 add_2750_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n53092), 
            .O(n7986[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_6 (.CI(n53092), .I0(n1557), .I1(n1011), .CO(n53093));
    SB_LUT4 add_2750_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n53091), 
            .O(n7986[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_5 (.CI(n53091), .I0(n1558), .I1(n856), .CO(n53092));
    SB_LUT4 add_2750_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n53090), 
            .O(n7986[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_4 (.CI(n53090), .I0(n1559), .I1(n698), .CO(n53091));
    SB_LUT4 add_2750_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n53089), 
            .O(n7986[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8168[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8012[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8194[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8194[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8220[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8246[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2750_3 (.CI(n53089), .I0(n1560), .I1(n858), .CO(n53090));
    SB_LUT4 i1_3_lut_4_lut_adj_1010 (.I0(n64363), .I1(n64503), .I2(n7986[14]), 
            .I3(n48_adj_5224), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1010.LUT_INIT = 16'h0010;
    SB_LUT4 add_2750_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7986[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .D(n32083));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .D(n55814));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n32231));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2750_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53089));
    SB_LUT4 add_2749_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n53088), 
            .O(n7960[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2749_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n53087), 
            .O(n7960[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_9 (.CI(n53087), .I0(n1409), .I1(n1602), .CO(n53088));
    SB_LUT4 add_2749_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n53086), 
            .O(n7960[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_8 (.CI(n53086), .I0(n1410), .I1(n1459), .CO(n53087));
    SB_LUT4 add_2749_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n53085), 
            .O(n7960[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_7 (.CI(n53085), .I0(n1411), .I1(n1460), .CO(n53086));
    SB_LUT4 add_2749_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n53084), 
            .O(n7960[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_6 (.CI(n53084), .I0(n1412), .I1(n1011), .CO(n53085));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n32087));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2749_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n53083), 
            .O(n7960[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_5 (.CI(n53083), .I0(n1413), .I1(n856), .CO(n53084));
    SB_LUT4 add_2749_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n53082), 
            .O(n7960[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_4 (.CI(n53082), .I0(n1414), .I1(n698), .CO(n53083));
    SB_LUT4 add_2749_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n53081), 
            .O(n7960[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8038[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2749_3 (.CI(n53081), .I0(n1415), .I1(n858), .CO(n53082));
    SB_LUT4 add_2749_2_lut (.I0(n61164), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2749_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53081));
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n32021));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n32020));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2748_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n53080), 
            .O(n7934[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5225), .I1(baudrate[9]), 
            .I2(n37_adj_5208), .I3(GND_net), .O(n34_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n31961));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2748_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n53079), 
            .O(n7934[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_8 (.CI(n53079), .I0(n1262), .I1(n1459), .CO(n53080));
    SB_LUT4 add_2748_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n53078), 
            .O(n7934[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_7 (.CI(n53078), .I0(n1263), .I1(n1460), .CO(n53079));
    SB_LUT4 add_2748_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n53077), 
            .O(n7934[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_6 (.CI(n53077), .I0(n1264), .I1(n1011), .CO(n53078));
    SB_LUT4 add_2748_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n53076), 
            .O(n7934[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_5 (.CI(n53076), .I0(n1265), .I1(n856), .CO(n53077));
    SB_LUT4 add_2748_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n53075), 
            .O(n7934[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_4 (.CI(n53075), .I0(n1266), .I1(n698), .CO(n53076));
    SB_LUT4 add_2748_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n53074), 
            .O(n7934[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_3 (.CI(n53074), .I0(n1267), .I1(n858), .CO(n53075));
    SB_LUT4 add_2748_2_lut (.I0(n61168), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2748_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53074));
    SB_LUT4 add_2747_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n53073), 
            .O(n7908[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1011 (.I0(n63627), .I1(n64447), .I2(n8064[11]), 
            .I3(n48_adj_5198), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1011.LUT_INIT = 16'h0010;
    SB_LUT4 add_2747_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n53072), 
            .O(n7908[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_7 (.CI(n53072), .I0(n1112), .I1(n1460), .CO(n53073));
    SB_LUT4 add_2747_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n53071), 
            .O(n7908[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_6 (.CI(n53071), .I0(n1113), .I1(n1011), .CO(n53072));
    SB_LUT4 add_2747_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n53070), 
            .O(n7908[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_5 (.CI(n53070), .I0(n1114), .I1(n856), .CO(n53071));
    SB_LUT4 i45242_2_lut_3_lut (.I0(n63627), .I1(n64447), .I2(baudrate[12]), 
            .I3(GND_net), .O(n64503));
    defparam i45242_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i51715_2_lut_3_lut (.I0(n63627), .I1(n64447), .I2(n48_adj_5198), 
            .I3(GND_net), .O(n294[11]));
    defparam i51715_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_2747_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n53069), 
            .O(n7908[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_4 (.CI(n53069), .I0(n1115), .I1(n698), .CO(n53070));
    SB_LUT4 add_2747_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n53068), 
            .O(n7908[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_3 (.CI(n53068), .I0(n1116), .I1(n858), .CO(n53069));
    SB_LUT4 add_2747_2_lut (.I0(n61172), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2747_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53068));
    SB_LUT4 i51359_4_lut (.I0(n34_adj_5226), .I1(n24_adj_5227), .I2(n37_adj_5208), 
            .I3(n68592), .O(n70629));   // verilog/uart_rx.v(119[33:55])
    defparam i51359_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2763_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n53314), 
            .O(n8324[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2763_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n53313), 
            .O(n8324[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_24 (.CI(n53313), .I0(n3152), .I1(n3082), .CO(n53314));
    SB_LUT4 add_2763_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n53312), 
            .O(n8324[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_23 (.CI(n53312), .I0(n3153), .I1(n3188), .CO(n53313));
    SB_LUT4 add_2763_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n53311), 
            .O(n8324[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_22 (.CI(n53311), .I0(n3154), .I1(n3084), .CO(n53312));
    SB_LUT4 add_2763_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n53310), 
            .O(n8324[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_21 (.CI(n53310), .I0(n3155), .I1(n2977), .CO(n53311));
    SB_LUT4 add_2763_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n53309), 
            .O(n8324[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_20 (.CI(n53309), .I0(n3156), .I1(n2867), .CO(n53310));
    SB_LUT4 add_2763_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n53308), 
            .O(n8324[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_19 (.CI(n53308), .I0(n3157), .I1(n2754), .CO(n53309));
    SB_LUT4 add_2763_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n53307), 
            .O(n8324[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_18 (.CI(n53307), .I0(n3158), .I1(n2638), .CO(n53308));
    SB_LUT4 add_2763_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n53306), 
            .O(n8324[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_17 (.CI(n53306), .I0(n3159), .I1(n2519), .CO(n53307));
    SB_LUT4 add_2763_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n53305), 
            .O(n8324[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_16 (.CI(n53305), .I0(n3160), .I1(n2397), .CO(n53306));
    SB_LUT4 add_2763_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n53304), 
            .O(n8324[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_15 (.CI(n53304), .I0(n3161), .I1(n2272), .CO(n53305));
    SB_LUT4 add_2763_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n53303), 
            .O(n8324[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_14 (.CI(n53303), .I0(n3162), .I1(n2144), .CO(n53304));
    SB_LUT4 add_2763_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n53302), 
            .O(n8324[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_13 (.CI(n53302), .I0(n3163), .I1(n2013), .CO(n53303));
    SB_LUT4 add_2763_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n53301), 
            .O(n8324[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_12 (.CI(n53301), .I0(n3164), .I1(n1879), .CO(n53302));
    SB_LUT4 add_2763_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n53300), 
            .O(n8324[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_11 (.CI(n53300), .I0(n3165), .I1(n1742), .CO(n53301));
    SB_LUT4 add_2763_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n53299), 
            .O(n8324[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_10 (.CI(n53299), .I0(n3166), .I1(n1602), .CO(n53300));
    SB_LUT4 add_2763_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n53298), 
            .O(n8324[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_9 (.CI(n53298), .I0(n3167), .I1(n1459), .CO(n53299));
    SB_LUT4 add_2763_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n53297), 
            .O(n8324[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_8 (.CI(n53297), .I0(n3168), .I1(n1460), .CO(n53298));
    SB_LUT4 add_2763_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n53296), 
            .O(n8324[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_7 (.CI(n53296), .I0(n3169), .I1(n1011), .CO(n53297));
    SB_LUT4 add_2763_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n53295), 
            .O(n8324[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_6 (.CI(n53295), .I0(n3170), .I1(n856), .CO(n53296));
    SB_LUT4 add_2763_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n53294), 
            .O(n8324[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_5 (.CI(n53294), .I0(n3171), .I1(n698), .CO(n53295));
    SB_LUT4 add_2763_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n53293), 
            .O(n8324[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2763_4 (.CI(n53293), .I0(n3172), .I1(n858), .CO(n53294));
    SB_LUT4 add_2763_3_lut (.I0(n61114), .I1(GND_net), .I2(n538), .I3(n53292), 
            .O(n63077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2763_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2763_3 (.CI(n53292), .I0(GND_net), .I1(n538), .CO(n53293));
    SB_CARRY add_2763_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n53292));
    SB_LUT4 add_2762_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n53291), 
            .O(n8298[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2762_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n53290), 
            .O(n8298[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_22 (.CI(n53290), .I0(n3047), .I1(n3188), .CO(n53291));
    SB_LUT4 add_2762_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n53289), 
            .O(n8298[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_21 (.CI(n53289), .I0(n3048), .I1(n3084), .CO(n53290));
    SB_LUT4 add_2762_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n53288), 
            .O(n8298[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_20 (.CI(n53288), .I0(n3049), .I1(n2977), .CO(n53289));
    SB_LUT4 add_2762_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n53287), 
            .O(n8298[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_19 (.CI(n53287), .I0(n3050), .I1(n2867), .CO(n53288));
    SB_LUT4 add_2762_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n53286), 
            .O(n8298[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_18 (.CI(n53286), .I0(n3051), .I1(n2754), .CO(n53287));
    SB_LUT4 add_2762_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n53285), 
            .O(n8298[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_17 (.CI(n53285), .I0(n3052), .I1(n2638), .CO(n53286));
    SB_LUT4 add_2762_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n53284), 
            .O(n8298[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_16 (.CI(n53284), .I0(n3053), .I1(n2519), .CO(n53285));
    SB_LUT4 add_2762_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n53283), 
            .O(n8298[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_15 (.CI(n53283), .I0(n3054), .I1(n2397), .CO(n53284));
    SB_LUT4 add_2762_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n53282), 
            .O(n8298[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_14 (.CI(n53282), .I0(n3055), .I1(n2272), .CO(n53283));
    SB_LUT4 add_2762_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n53281), 
            .O(n8298[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_13 (.CI(n53281), .I0(n3056), .I1(n2144), .CO(n53282));
    SB_LUT4 add_2762_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n53280), 
            .O(n8298[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_12 (.CI(n53280), .I0(n3057), .I1(n2013), .CO(n53281));
    SB_LUT4 add_2762_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n53279), 
            .O(n8298[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_11 (.CI(n53279), .I0(n3058), .I1(n1879), .CO(n53280));
    SB_LUT4 add_2762_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n53278), 
            .O(n8298[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_10 (.CI(n53278), .I0(n3059), .I1(n1742), .CO(n53279));
    SB_LUT4 add_2762_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n53277), 
            .O(n8298[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_9 (.CI(n53277), .I0(n3060), .I1(n1602), .CO(n53278));
    SB_LUT4 add_2762_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n53276), 
            .O(n8298[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_8 (.CI(n53276), .I0(n3061), .I1(n1459), .CO(n53277));
    SB_LUT4 add_2762_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n53275), 
            .O(n8298[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_7 (.CI(n53275), .I0(n3062), .I1(n1460), .CO(n53276));
    SB_LUT4 add_2762_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n53274), 
            .O(n8298[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_6 (.CI(n53274), .I0(n3063), .I1(n1011), .CO(n53275));
    SB_LUT4 add_2762_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n53273), 
            .O(n8298[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_5 (.CI(n53273), .I0(n3064), .I1(n856), .CO(n53274));
    SB_LUT4 add_2762_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n53272), 
            .O(n8298[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_4 (.CI(n53272), .I0(n3065), .I1(n698), .CO(n53273));
    SB_LUT4 add_2762_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n53271), 
            .O(n8298[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2762_3 (.CI(n53271), .I0(n3066), .I1(n858), .CO(n53272));
    SB_LUT4 i51360_3_lut (.I0(n70629), .I1(baudrate[10]), .I2(n39_adj_5207), 
            .I3(GND_net), .O(n70630));   // verilog/uart_rx.v(119[33:55])
    defparam i51360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2762_2_lut (.I0(n61118), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2762_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2762_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53271));
    SB_LUT4 add_2761_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n53270), 
            .O(n8272[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2761_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n53269), 
            .O(n8272[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_21 (.CI(n53269), .I0(n2939), .I1(n3084), .CO(n53270));
    SB_LUT4 add_2761_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n53268), 
            .O(n8272[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_20 (.CI(n53268), .I0(n2940), .I1(n2977), .CO(n53269));
    SB_LUT4 add_2761_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n53267), 
            .O(n8272[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2761_19 (.CI(n53267), .I0(n2941), .I1(n2867), .CO(n53268));
    SB_LUT4 add_2761_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n53266), 
            .O(n8272[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_18 (.CI(n53266), .I0(n2942), .I1(n2754), .CO(n53267));
    SB_LUT4 add_2761_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n53265), 
            .O(n8272[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_17 (.CI(n53265), .I0(n2943), .I1(n2638), .CO(n53266));
    SB_LUT4 add_2761_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n53264), 
            .O(n8272[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_16 (.CI(n53264), .I0(n2944), .I1(n2519), .CO(n53265));
    SB_LUT4 add_2761_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n53263), 
            .O(n8272[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_15 (.CI(n53263), .I0(n2945), .I1(n2397), .CO(n53264));
    SB_LUT4 add_2761_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n53262), 
            .O(n8272[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_14 (.CI(n53262), .I0(n2946), .I1(n2272), .CO(n53263));
    SB_LUT4 add_2761_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n53261), 
            .O(n8272[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_13 (.CI(n53261), .I0(n2947), .I1(n2144), .CO(n53262));
    SB_LUT4 i1_4_lut_adj_1012 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n63785));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5229));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(r_Clock_Count[3]), .I1(n3_adj_5229), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n63785), .O(n63789));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hffde;
    SB_LUT4 add_2761_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n53260), 
            .O(n8272[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_12 (.CI(n53260), .I0(n2948), .I1(n2013), .CO(n53261));
    SB_LUT4 add_2761_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n53259), 
            .O(n8272[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_11 (.CI(n53259), .I0(n2949), .I1(n1879), .CO(n53260));
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49271_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5232), .I3(\o_Rx_DV_N_3488[8] ), .O(n67700));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49271_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n63789), .O(n63793));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hffde;
    SB_LUT4 i49394_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n59720), 
            .I3(r_SM_Main[0]), .O(n67706));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49394_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5230));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49268_4_lut (.I0(n67700), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67697));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49268_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49276_4_lut (.I0(n67706), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67703));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49276_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 add_2761_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n53258), 
            .O(n8272[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_10 (.CI(n53258), .I0(n2950), .I1(n1742), .CO(n53259));
    SB_LUT4 add_2761_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n53257), 
            .O(n8272[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2761_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2761_9 (.CI(n53257), .I0(n2951), .I1(n1602), .CO(n53258));
    SB_LUT4 i1_4_lut_adj_1015 (.I0(r_Clock_Count[6]), .I1(n8_adj_5230), 
            .I2(n63793), .I3(\o_Rx_DV_N_3488[7] ), .O(n59720));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'hfdfe;
    SB_LUT4 equal_347_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(98[17:39])
    defparam equal_347_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n59686));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i45170_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n59720), .I2(GND_net), 
            .I3(GND_net), .O(n64431));
    defparam i45170_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45292_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n64431), .O(n64553));
    defparam i45292_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n63199), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n64553), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n10015));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n10015), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n67703), .I1(n67697), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_5129));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i51204_3_lut (.I0(n70630), .I1(baudrate[11]), .I2(n41_adj_5206), 
            .I3(GND_net), .O(n70474));   // verilog/uart_rx.v(119[33:55])
    defparam i51204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51080_4_lut (.I0(n41_adj_5206), .I1(n39_adj_5207), .I2(n37_adj_5208), 
            .I3(n68594), .O(n70350));
    defparam i51080_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51116_4_lut (.I0(n30_adj_5223), .I1(n22_adj_5221), .I2(n33_adj_5203), 
            .I3(n68600), .O(n70386));   // verilog/uart_rx.v(119[33:55])
    defparam i51116_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8064[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49876_3_lut (.I0(n70474), .I1(baudrate[12]), .I2(n43_adj_5202), 
            .I3(GND_net), .O(n69146));   // verilog/uart_rx.v(119[33:55])
    defparam i49876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8168[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8194[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8220[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8142[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8168[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8090[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8194[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8220[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n63895));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8142[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8168[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45228_3_lut (.I0(baudrate[19]), .I1(baudrate[4]), .I2(baudrate[20]), 
            .I3(GND_net), .O(n64489));
    defparam i45228_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8194[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8220[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n63623));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n63625));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n63629));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n63631));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'heeee;
    SB_LUT4 i51341_4_lut (.I0(n69146), .I1(n70386), .I2(n43_adj_5202), 
            .I3(n70350), .O(n70611));   // verilog/uart_rx.v(119[33:55])
    defparam i51341_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n63633));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n63637));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 i23780_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n41626));
    defparam i23780_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23778_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n41624));
    defparam i23778_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6222_4_lut (.I0(n804), .I1(n41624), .I2(n23812), .I3(baudrate[2]), 
            .O(n23826));   // verilog/uart_rx.v(119[33:55])
    defparam i6222_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i6262_4_lut (.I0(n960), .I1(n9792), .I2(n23867), .I3(n856), 
            .O(n23869));   // verilog/uart_rx.v(119[33:55])
    defparam i6262_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51342_3_lut (.I0(n70611), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n70612));   // verilog/uart_rx.v(119[33:55])
    defparam i51342_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45009_2_lut (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n63893));
    defparam i45009_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63601));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n63849));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49351_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n68621));
    defparam i49351_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1025 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n63903));
    defparam i1_2_lut_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1026 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n63905));
    defparam i1_2_lut_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1027 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n63769));
    defparam i1_2_lut_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59971));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[8]), .I1(baudrate[9]), .I2(baudrate[10]), 
            .I3(baudrate[11]), .O(n63771));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5240));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5232), 
            .O(n15_adj_5241));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8142[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5241), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5240), 
            .I3(n59971), .O(n71701));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i41911_1_lut (.I0(n27736), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61134));
    defparam i41911_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8168[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45184_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), .I2(n27736), 
            .I3(GND_net), .O(n64445));
    defparam i45184_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8194[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4034_2_lut_4_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam i4034_2_lut_4_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63797));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'heeee;
    SB_LUT4 i41895_1_lut (.I0(n27748), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61118));
    defparam i41895_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n63889));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n63993));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'heeee;
    SB_LUT4 i49475_2_lut (.I0(n59720), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n67642));
    defparam i49475_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i49470_4_lut (.I0(n67642), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n67639));
    defparam i49470_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48595_4_lut (.I0(n67639), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n67636));
    defparam i48595_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i51788_4_lut (.I0(\r_SM_Main[2] ), .I1(n67636), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(\r_SM_Main[1] ), .O(n31162));
    defparam i51788_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(n59720), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n63131));
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n63131), .O(n63137));
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'h0100;
    SB_LUT4 i51680_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n63137), .O(n29942));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51680_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1034 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[4]), .I3(baudrate[5]), .O(n63773));
    defparam i1_2_lut_3_lut_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n63897), .I1(n63893), .I2(n63895), 
            .I3(n63891), .O(n63877));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 i45212_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n64473));
    defparam i45212_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1036 (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n63807));
    defparam i1_2_lut_3_lut_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(n63993), .I1(n63807), .I2(n63889), 
            .I3(n63797), .O(n27748));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'hfffe;
    SB_LUT4 i45271_1_lut (.I0(n64531), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61172));
    defparam i45271_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51893_2_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n29821));
    defparam i51893_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i4039_2_lut_2_lut_4_lut (.I0(baudrate[2]), .I1(n805), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n9628));   // verilog/uart_rx.v(119[33:55])
    defparam i4039_2_lut_2_lut_4_lut.LUT_INIT = 16'h0445;
    SB_LUT4 equal_345_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(98[17:39])
    defparam equal_345_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i23791_rep_5_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n61175));   // verilog/uart_rx.v(119[33:55])
    defparam i23791_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45185_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n27736), .I3(GND_net), .O(n61142));
    defparam i45185_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i45267_1_lut (.I0(n64527), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61164));
    defparam i45267_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n61175), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8220[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1038 (.I0(n63821), .I1(n63897), .I2(n63895), 
            .I3(n63893), .O(n63775));
    defparam i1_2_lut_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 i51221_3_lut (.I0(n42_adj_5244), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n70491));   // verilog/uart_rx.v(119[33:55])
    defparam i51221_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49419_2_lut_3_lut (.I0(n27648), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n67685));   // verilog/uart_rx.v(119[33:55])
    defparam i49419_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut_4_lut_adj_1039 (.I0(n59686), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(\r_SM_Main[1] ), .O(n63175));
    defparam i1_3_lut_4_lut_adj_1039.LUT_INIT = 16'hfdfc;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8116[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23738_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n41584));
    defparam i23738_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51222_3_lut (.I0(n70491), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n70492));   // verilog/uart_rx.v(119[33:55])
    defparam i51222_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45269_1_lut_2_lut (.I0(baudrate[8]), .I1(n64527), .I2(GND_net), 
            .I3(GND_net), .O(n61168));
    defparam i45269_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i50930_3_lut (.I0(n70492), .I1(baudrate[5]), .I2(n60874), 
            .I3(GND_net), .O(n48_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam i50930_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_2_lut_4_lut_adj_1040 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n63833));
    defparam i1_2_lut_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(n63835), .I1(n27748), .I2(n63877), 
            .I3(n63833), .O(n27700));
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8142[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1042 (.I0(n27700), .I1(n48_adj_5245), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1042.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7908[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8168[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4210_2_lut_2_lut (.I0(baudrate[3]), .I1(n42_adj_5094), .I2(GND_net), 
            .I3(GND_net), .O(n9799));   // verilog/uart_rx.v(119[33:55])
    defparam i4210_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8220[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6210_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n23812));   // verilog/uart_rx.v(119[33:55])
    defparam i6210_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i45153_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n64413));
    defparam i45153_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7934[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7960[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49457_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5232), .I3(n59971), .O(n67656));
    defparam i49457_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i49453_4_lut (.I0(n67656), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67653));
    defparam i49453_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n67653), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n29817));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8246[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8194[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n63765));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n63743));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(n63743), .I1(n63903), .I2(n63847), 
            .I3(n63843), .O(n27742));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n67685), .I1(baudrate[2]), 
            .I2(n70911), .I3(n48_adj_5072), .O(n46_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5249), .I1(baudrate[3]), 
            .I2(n60868), .I3(GND_net), .O(n48_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n63773), .I1(n27742), .I2(n63775), 
            .I3(n63771), .O(n27694));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63843));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1048 (.I0(n27694), .I1(n48_adj_5250), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1048.LUT_INIT = 16'hefef;
    SB_LUT4 i45079_1_lut_2_lut (.I0(baudrate[17]), .I1(n27736), .I2(GND_net), 
            .I3(GND_net), .O(n61138));
    defparam i45079_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i51709_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n64503), .I3(n48_adj_5224), .O(n294[14]));
    defparam i51709_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i45266_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n64503), .I3(baudrate[9]), .O(n64527));
    defparam i45266_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45214_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n64475));
    defparam i45214_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i50913_3_lut (.I0(n32_adj_5251), .I1(baudrate[5]), .I2(n39_adj_5248), 
            .I3(GND_net), .O(n70183));   // verilog/uart_rx.v(119[33:55])
    defparam i50913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45280_4_lut (.I0(n64475), .I1(n63889), .I2(n64473), .I3(n63843), 
            .O(n64541));
    defparam i45280_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45281_1_lut (.I0(n64541), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61122));
    defparam i45281_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49322_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n68592));
    defparam i49322_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50914_3_lut (.I0(n70183), .I1(baudrate[6]), .I2(n41_adj_5247), 
            .I3(GND_net), .O(n70184));   // verilog/uart_rx.v(119[33:55])
    defparam i50914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49330_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n68600));
    defparam i49330_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49282_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n68552));
    defparam i49282_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50392_4_lut (.I0(n41_adj_5247), .I1(n39_adj_5248), .I2(n37_adj_5246), 
            .I3(n68753), .O(n69662));
    defparam i50392_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50935_3_lut (.I0(n34_adj_5252), .I1(baudrate[4]), .I2(n37_adj_5246), 
            .I3(GND_net), .O(n70205));   // verilog/uart_rx.v(119[33:55])
    defparam i50935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49288_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n68558));
    defparam i49288_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49848_3_lut (.I0(n70184), .I1(baudrate[7]), .I2(n43_adj_5242), 
            .I3(GND_net), .O(n69118));   // verilog/uart_rx.v(119[33:55])
    defparam i49848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51215_4_lut (.I0(n69118), .I1(n70205), .I2(n43_adj_5242), 
            .I3(n69662), .O(n70485));   // verilog/uart_rx.v(119[33:55])
    defparam i51215_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i4197_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam i4197_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49380_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n68650));
    defparam i49380_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51216_3_lut (.I0(n70485), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n70486));   // verilog/uart_rx.v(119[33:55])
    defparam i51216_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n70486), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2318_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2318_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8012[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49079_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n68349));
    defparam i49079_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8038[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5253), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8064[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41619_2_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n60834));
    defparam i41619_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5232), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n59686), .O(n63167));
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n63167), .O(n63173));
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(n63173), .I1(n6), .I2(\r_SM_Main[1] ), 
            .I3(n27), .O(n31149));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'h0323;
    SB_LUT4 i51706_2_lut_4_lut (.I0(n70203), .I1(baudrate[8]), .I2(n1408), 
            .I3(n64527), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i51706_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1052 (.I0(n70203), .I1(baudrate[8]), .I2(n1408), 
            .I3(n63057), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1052.LUT_INIT = 16'h7100;
    SB_LUT4 i2311_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2311_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8090[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49413_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n68683));
    defparam i49413_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7908[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8116[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45270_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n64527), 
            .I3(GND_net), .O(n64531));
    defparam i45270_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8142[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i41891_1_lut_4_lut (.I0(n63995), .I1(n63997), .I2(n63845), 
            .I3(n63993), .O(n61114));
    defparam i41891_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i49051_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n68321));
    defparam i49051_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49145_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n68415));
    defparam i49145_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49111_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n68381));
    defparam i49111_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8168[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8194[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7934[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7960[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7986[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8012[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7934[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8324[20]), .I3(n294[1]), .O(n41_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8038[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8324[19]), .I3(n294[1]), .O(n39_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8324[16]), .I3(n294[1]), .O(n33_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_4_lut_adj_1053 (.I0(n70490), .I1(baudrate[7]), .I2(n1261), 
            .I3(n63055), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1053.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8324[17]), .I3(n294[1]), .O(n35_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i49022_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n68292));
    defparam i49022_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49206_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n68476));
    defparam i49206_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7960[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8324[18]), .I3(n294[1]), .O(n37_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8324[14]), .I3(n294[1]), .O(n29_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8324[15]), .I3(n294[1]), .O(n31_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8324[11]), .I3(n294[1]), .O(n23_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i48988_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n68258));
    defparam i48988_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8324[12]), .I3(n294[1]), .O(n25_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i45243_1_lut (.I0(n64503), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61155));
    defparam i45243_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8324[22]), .I3(n294[1]), .O(n45_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8324[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8064[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8090[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8324[4]), .I3(n294[1]), .O(n9_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7986[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49219_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n68489));
    defparam i49219_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1054 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n63009));
    defparam i1_3_lut_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8324[8]), .I3(n294[1]), .O(n17_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8116[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8142[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8324[9]), .I3(n294[1]), .O(n19_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8324[10]), .I3(n294[1]), .O(n21_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8324[21]), .I3(n294[1]), .O(n43_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8168[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8194[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51791_2_lut_4_lut (.I0(n70765), .I1(baudrate[13]), .I2(n2098), 
            .I3(n27724), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i51791_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8324[5]), .I3(n294[1]), .O(n11_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1055 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[9]), .I3(baudrate[8]), .O(n63835));
    defparam i1_2_lut_3_lut_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8324[6]), .I3(n294[1]), .O(n13_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8324[7]), .I3(n294[1]), .O(n15_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8324[13]), .I3(n294[1]), .O(n27_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i48701_4_lut (.I0(n27_adj_5272), .I1(n15_adj_5271), .I2(n13_adj_5270), 
            .I3(n11_adj_5269), .O(n67971));
    defparam i48701_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8012[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4205_2_lut_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam i4205_2_lut_4_lut.LUT_INIT = 16'hb2bb;
    SB_LUT4 i51782_2_lut_4_lut (.I0(n70484), .I1(baudrate[10]), .I2(n1693), 
            .I3(n27715), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i51782_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i48709_4_lut (.I0(n21_adj_5267), .I1(n19_adj_5266), .I2(n17_adj_5265), 
            .I3(n9_adj_5264), .O(n67979));
    defparam i48709_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5268), .I3(GND_net), .O(n16_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7908[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48666_2_lut (.I0(n43_adj_5268), .I1(n19_adj_5266), .I2(GND_net), 
            .I3(GND_net), .O(n67936));
    defparam i48666_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5265), .I3(GND_net), .O(n8_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5273), .I1(baudrate[22]), 
            .I2(n45_adj_5263), .I3(GND_net), .O(n24_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8324[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48755_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n68025));
    defparam i48755_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i49749_4_lut (.I0(n13_adj_5270), .I1(n11_adj_5269), .I2(n9_adj_5264), 
            .I3(n68025), .O(n69019));
    defparam i49749_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49737_4_lut (.I0(n19_adj_5266), .I1(n17_adj_5265), .I2(n15_adj_5271), 
            .I3(n69019), .O(n69007));
    defparam i49737_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51161_4_lut (.I0(n25_adj_5262), .I1(n23_adj_5261), .I2(n21_adj_5267), 
            .I3(n69007), .O(n70431));
    defparam i51161_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50502_4_lut (.I0(n31_adj_5260), .I1(n29_adj_5259), .I2(n27_adj_5272), 
            .I3(n70431), .O(n69772));
    defparam i50502_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51403_4_lut (.I0(n37_adj_5258), .I1(n35_adj_5257), .I2(n33_adj_5256), 
            .I3(n69772), .O(n70673));
    defparam i51403_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5256), .I3(GND_net), .O(n12_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63077), .I3(n48), .O(n4_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i51096_3_lut (.I0(n4_adj_5278), .I1(baudrate[13]), .I2(n27_adj_5272), 
            .I3(GND_net), .O(n70366));   // verilog/uart_rx.v(119[33:55])
    defparam i51096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51097_3_lut (.I0(n70366), .I1(baudrate[14]), .I2(n29_adj_5259), 
            .I3(GND_net), .O(n70367));   // verilog/uart_rx.v(119[33:55])
    defparam i51097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48685_2_lut (.I0(n33_adj_5256), .I1(n15_adj_5271), .I2(GND_net), 
            .I3(GND_net), .O(n67955));
    defparam i48685_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8038[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8064[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5270), .I3(GND_net), .O(n10_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5277), .I1(baudrate[17]), 
            .I2(n35_adj_5257), .I3(GND_net), .O(n30_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8090[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48691_4_lut (.I0(n33_adj_5256), .I1(n31_adj_5260), .I2(n29_adj_5259), 
            .I3(n67971), .O(n67961));
    defparam i48691_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_adj_1056 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n63865));
    defparam i1_2_lut_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i51462_4_lut (.I0(n30_adj_5280), .I1(n10_adj_5279), .I2(n35_adj_5257), 
            .I3(n67955), .O(n70732));   // verilog/uart_rx.v(119[33:55])
    defparam i51462_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50973_3_lut (.I0(n70367), .I1(baudrate[15]), .I2(n31_adj_5260), 
            .I3(GND_net), .O(n70243));   // verilog/uart_rx.v(119[33:55])
    defparam i50973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51607_4_lut (.I0(n70243), .I1(n70732), .I2(n35_adj_5257), 
            .I3(n67961), .O(n70877));   // verilog/uart_rx.v(119[33:55])
    defparam i51607_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51608_3_lut (.I0(n70877), .I1(baudrate[18]), .I2(n37_adj_5258), 
            .I3(GND_net), .O(n70878));   // verilog/uart_rx.v(119[33:55])
    defparam i51608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5282), .I1(baudrate[4]), 
            .I2(n41_adj_5274), .I3(GND_net), .O(n40_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51347_4_lut (.I0(n40_adj_5283), .I1(n36_adj_5281), .I2(n41_adj_5274), 
            .I3(n68788), .O(n70617));   // verilog/uart_rx.v(119[33:55])
    defparam i51347_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8116[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51348_3_lut (.I0(n70617), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n70618));   // verilog/uart_rx.v(119[33:55])
    defparam i51348_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51100_3_lut (.I0(n6_adj_5284), .I1(baudrate[10]), .I2(n21_adj_5267), 
            .I3(GND_net), .O(n70370));   // verilog/uart_rx.v(119[33:55])
    defparam i51100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8142[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51101_3_lut (.I0(n70370), .I1(baudrate[11]), .I2(n23_adj_5261), 
            .I3(GND_net), .O(n70371));   // verilog/uart_rx.v(119[33:55])
    defparam i51101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48671_4_lut (.I0(n43_adj_5268), .I1(n25_adj_5262), .I2(n23_adj_5261), 
            .I3(n67979), .O(n67941));
    defparam i48671_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50584_4_lut (.I0(n24_adj_5276), .I1(n8_adj_5275), .I2(n45_adj_5263), 
            .I3(n67936), .O(n69854));   // verilog/uart_rx.v(119[33:55])
    defparam i50584_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50971_3_lut (.I0(n70371), .I1(baudrate[12]), .I2(n25_adj_5262), 
            .I3(GND_net), .O(n70241));   // verilog/uart_rx.v(119[33:55])
    defparam i50971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51544_3_lut (.I0(n70878), .I1(baudrate[19]), .I2(n39_adj_5255), 
            .I3(GND_net), .O(n70814));   // verilog/uart_rx.v(119[33:55])
    defparam i51544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8168[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48673_4_lut (.I0(n43_adj_5268), .I1(n41_adj_5254), .I2(n39_adj_5255), 
            .I3(n70673), .O(n67943));
    defparam i48673_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51251_4_lut (.I0(n70241), .I1(n69854), .I2(n45_adj_5263), 
            .I3(n67941), .O(n70521));   // verilog/uart_rx.v(119[33:55])
    defparam i51251_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51516_3_lut (.I0(n70814), .I1(baudrate[20]), .I2(n41_adj_5254), 
            .I3(GND_net), .O(n40_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam i51516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63029));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8324[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51253_4_lut (.I0(n40_adj_5285), .I1(n70521), .I2(n45_adj_5263), 
            .I3(n67943), .O(n70523));   // verilog/uart_rx.v(119[33:55])
    defparam i51253_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n63991), .I1(n63847), .I2(n63029), 
            .I3(n63845), .O(n63037));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 i48752_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5250), .I2(n27694), 
            .I3(GND_net), .O(n68022));   // verilog/uart_rx.v(119[33:55])
    defparam i48752_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i51799_4_lut (.I0(n63037), .I1(n70523), .I2(baudrate[23]), 
            .I3(n3253), .O(n61968));   // verilog/uart_rx.v(119[33:55])
    defparam i51799_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8194[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1059 (.I0(n70616), .I1(baudrate[6]), .I2(n1111), 
            .I3(n63053), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1059.LUT_INIT = 16'h7100;
    SB_LUT4 i51694_2_lut_4_lut (.I0(n70616), .I1(baudrate[6]), .I2(n1111), 
            .I3(n64531), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i51694_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8194[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1060 (.I0(n69850), .I1(baudrate[21]), .I2(n3046), 
            .I3(n63075), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1060.LUT_INIT = 16'h7100;
    SB_LUT4 i51880_2_lut_4_lut (.I0(n69850), .I1(baudrate[21]), .I2(n3046), 
            .I3(n27748), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i51880_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4203_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9792));   // verilog/uart_rx.v(119[33:55])
    defparam i4203_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45186_2_lut (.I0(baudrate[15]), .I1(n64445), .I2(GND_net), 
            .I3(GND_net), .O(n64447));
    defparam i45186_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45187_1_lut_2_lut (.I0(baudrate[15]), .I1(n64445), .I2(GND_net), 
            .I3(GND_net), .O(n61146));
    defparam i45187_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i51685_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n64531), .I3(n48_adj_5031), .O(n294[19]));
    defparam i51685_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n63627));
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48897_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n68167));
    defparam i48897_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48936_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n68206));
    defparam i48936_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51697_2_lut_4_lut (.I0(n70490), .I1(baudrate[7]), .I2(n1261), 
            .I3(n64529), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i51697_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_1062 (.I0(n27648), .I1(n48_adj_5072), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44));
    defparam i1_3_lut_4_lut_adj_1062.LUT_INIT = 16'hefff;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8298[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8298[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8298[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8298[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8298[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8298[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48744_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5072), .I2(n27648), 
            .I3(GND_net), .O(n68014));   // verilog/uart_rx.v(119[33:55])
    defparam i48744_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_4_lut_adj_1063 (.I0(n70612), .I1(baudrate[14]), .I2(n2227), 
            .I3(n63061), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1063.LUT_INIT = 16'h7100;
    SB_LUT4 i51762_2_lut_4_lut (.I0(n70612), .I1(baudrate[14]), .I2(n2227), 
            .I3(n64447), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i51762_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8298[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8298[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7960[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7986[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8012[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8038[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8298[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8064[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8090[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49244_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n68514));
    defparam i49244_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8116[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8142[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8168[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n63897));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n63821));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'heeee;
    SB_LUT4 i45232_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n64493));
    defparam i45232_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n64363));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51883_2_lut_4_lut (.I0(n70662), .I1(baudrate[22]), .I2(n3151), 
            .I3(n27751), .O(n294[1]));
    defparam i51883_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8298[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8298[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1067 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n63007));
    defparam i1_3_lut_4_lut_adj_1067.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n63891));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'heeee;
    SB_LUT4 i49503_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n68773));   // verilog/uart_rx.v(119[33:55])
    defparam i49503_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i41679_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n60900));
    defparam i41679_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45159_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n64419));
    defparam i45159_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45288_4_lut (.I0(n64419), .I1(n63769), .I2(n64363), .I3(baudrate[9]), 
            .O(n64549));
    defparam i45288_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1069 (.I0(baudrate[17]), .I1(n63637), .I2(baudrate[2]), 
            .I3(n41624), .O(n62985));
    defparam i1_4_lut_adj_1069.LUT_INIT = 16'h0100;
    SB_LUT4 i45264_4_lut (.I0(n63631), .I1(n63627), .I2(n63629), .I3(n63625), 
            .O(n64525));
    defparam i45264_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49536_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n68806));   // verilog/uart_rx.v(119[33:55])
    defparam i49536_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_4_lut_adj_1070 (.I0(n64525), .I1(n62985), .I2(n27736), 
            .I3(n64413), .O(n62075));
    defparam i1_4_lut_adj_1070.LUT_INIT = 16'h0004;
    SB_LUT4 i49518_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n68788));   // verilog/uart_rx.v(119[33:55])
    defparam i49518_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n41626), .O(n63339));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'h0100;
    SB_LUT4 i49483_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n68753));   // verilog/uart_rx.v(119[33:55])
    defparam i49483_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49460_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n68730));   // verilog/uart_rx.v(119[33:55])
    defparam i49460_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(n63339), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n63357));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'h0002;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5286));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49372_4_lut (.I0(n33_adj_5233), .I1(n31_adj_5231), .I2(n29_adj_5232), 
            .I3(n27_adj_5286), .O(n68642));
    defparam i49372_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48795_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n68065));
    defparam i48795_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45302_4_lut (.I0(n64493), .I1(n64413), .I2(n64489), .I3(n63623), 
            .O(n64563));
    defparam i45302_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5239), .I1(baudrate[10]), 
            .I2(n41_adj_5237), .I3(GND_net), .O(n38_adj_5287));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8298[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1073 (.I0(n64549), .I1(n64563), .I2(n60900), 
            .I3(n63357), .O(n61643));
    defparam i1_4_lut_adj_1073.LUT_INIT = 16'h0100;
    SB_LUT4 i23831_rep_3_2_lut (.I0(n8064[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n61149));   // verilog/uart_rx.v(119[33:55])
    defparam i23831_rep_3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8298[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1074 (.I0(n63629), .I1(n63625), .I2(n63627), 
            .I3(n63623), .O(n63647));
    defparam i1_4_lut_adj_1074.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8298[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n61149), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5288));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50901_3_lut (.I0(n26_adj_5288), .I1(baudrate[6]), .I2(n33_adj_5233), 
            .I3(GND_net), .O(n70171));   // verilog/uart_rx.v(119[33:55])
    defparam i50901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50902_3_lut (.I0(n70171), .I1(baudrate[7]), .I2(n35_adj_5234), 
            .I3(GND_net), .O(n70172));   // verilog/uart_rx.v(119[33:55])
    defparam i50902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49360_4_lut (.I0(n39_adj_5235), .I1(n37_adj_5236), .I2(n35_adj_5234), 
            .I3(n68642), .O(n68630));
    defparam i49360_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51357_4_lut (.I0(n38_adj_5287), .I1(n28_adj_5238), .I2(n41_adj_5237), 
            .I3(n68621), .O(n70627));   // verilog/uart_rx.v(119[33:55])
    defparam i51357_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51772_2_lut_4_lut (.I0(n70492), .I1(baudrate[5]), .I2(n60874), 
            .I3(n27700), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i51772_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i49864_3_lut (.I0(n70172), .I1(baudrate[8]), .I2(n37_adj_5236), 
            .I3(GND_net), .O(n69134));   // verilog/uart_rx.v(119[33:55])
    defparam i49864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48843_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n68113));
    defparam i48843_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n63997));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i51557_4_lut (.I0(n69134), .I1(n70627), .I2(n41_adj_5237), 
            .I3(n68630), .O(n70827));   // verilog/uart_rx.v(119[33:55])
    defparam i51557_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51558_3_lut (.I0(n70827), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n70828));   // verilog/uart_rx.v(119[33:55])
    defparam i51558_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n63637), .I1(n63633), .I2(n63635), 
            .I3(n63631), .O(n63649));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1076 (.I0(n63649), .I1(n27739), .I2(n63647), 
            .I3(GND_net), .O(n27648));
    defparam i1_3_lut_adj_1076.LUT_INIT = 16'hfefe;
    SB_LUT4 i51495_3_lut (.I0(n70828), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n70765));   // verilog/uart_rx.v(119[33:55])
    defparam i51495_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n61643), .I1(baudrate[2]), 
            .I2(n62075), .I3(GND_net), .O(n48_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i45078_2_lut (.I0(baudrate[17]), .I1(n27736), .I2(GND_net), 
            .I3(GND_net), .O(n64337));
    defparam i45078_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i49870_3_lut (.I0(n70765), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5289));   // verilog/uart_rx.v(119[33:55])
    defparam i49870_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51703_2_lut (.I0(n48_adj_5072), .I1(n27648), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i51703_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1077 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n63899));
    defparam i1_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8298[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51769_2_lut (.I0(n48_adj_5250), .I1(n27694), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i51769_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1078 (.I0(n63833), .I1(n63897), .I2(baudrate[16]), 
            .I3(n41624), .O(n63691));
    defparam i1_4_lut_adj_1078.LUT_INIT = 16'h0100;
    SB_LUT4 i49541_3_lut (.I0(n61643), .I1(n62075), .I2(baudrate[2]), 
            .I3(GND_net), .O(n67620));   // verilog/uart_rx.v(119[33:55])
    defparam i49541_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8298[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8298[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1079 (.I0(n63849), .I1(n63897), .I2(n63601), 
            .I3(GND_net), .O(n63907));
    defparam i1_3_lut_adj_1079.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(n63907), .I1(n63903), .I2(n63905), 
            .I3(n63899), .O(n27724));
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'hfffe;
    SB_LUT4 i49382_4_lut (.I0(n60900), .I1(n63691), .I2(n63835), .I3(n63765), 
            .O(n67621));   // verilog/uart_rx.v(119[33:55])
    defparam i49382_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n67621), .I1(n67620), .I2(n294[21]), 
            .I3(n64337), .O(n60868));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_4_lut_adj_1081 (.I0(n70219), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63065), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1081.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8012[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51811_2_lut_4_lut (.I0(n70219), .I1(baudrate[16]), .I2(n2476), 
            .I3(n64337), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i51811_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_adj_1082 (.I0(n27724), .I1(n48_adj_5289), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1082.LUT_INIT = 16'hefef;
    SB_LUT4 i49249_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n68519));
    defparam i49249_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (clk16MHz, n29799, \current[15] , n31638, \current[1] , 
            n31637, \current[2] , n31636, \current[3] , n31635, \current[4] , 
            n31634, \current[5] , n31633, \current[6] , n31632, \current[7] , 
            n31631, \current[8] , n31630, \current[9] , n31629, \current[10] , 
            n31628, \current[11] , state_7__N_4319, GND_net, VCC_net, 
            CS_c, n31471, \current[0] , n32396, \data[15] , n32395, 
            \data[12] , n32394, \data[11] , n32393, \data[10] , n32392, 
            \data[9] , n32391, \data[8] , n32390, \data[7] , n32389, 
            \data[6] , n32388, \data[5] , n32387, \data[4] , n32386, 
            \data[3] , n32385, \data[2] , n32384, \data[1] , n32101, 
            \data[0] , CS_CLK_c, n27661, n27667, n11, n27680, n27643, 
            n5, n5_adj_4, n41527, n9) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output n29799;
    output \current[15] ;
    input n31638;
    output \current[1] ;
    input n31637;
    output \current[2] ;
    input n31636;
    output \current[3] ;
    input n31635;
    output \current[4] ;
    input n31634;
    output \current[5] ;
    input n31633;
    output \current[6] ;
    input n31632;
    output \current[7] ;
    input n31631;
    output \current[8] ;
    input n31630;
    output \current[9] ;
    input n31629;
    output \current[10] ;
    input n31628;
    output \current[11] ;
    output state_7__N_4319;
    input GND_net;
    input VCC_net;
    output CS_c;
    input n31471;
    output \current[0] ;
    input n32396;
    output \data[15] ;
    input n32395;
    output \data[12] ;
    input n32394;
    output \data[11] ;
    input n32393;
    output \data[10] ;
    input n32392;
    output \data[9] ;
    input n32391;
    output \data[8] ;
    input n32390;
    output \data[7] ;
    input n32389;
    output \data[6] ;
    input n32388;
    output \data[5] ;
    input n32387;
    output \data[4] ;
    input n32386;
    output \data[3] ;
    input n32385;
    output \data[2] ;
    input n32384;
    output \data[1] ;
    input n32101;
    output \data[0] ;
    output CS_CLK_c;
    output n27661;
    output n27667;
    output n11;
    output n27680;
    output n27643;
    output n5;
    output n5_adj_4;
    output n41527;
    output n9;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire clk_slow_N_4232;
    wire [13:0]n241;
    wire [7:0]n37;
    
    wire n29937;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n31405;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n24764;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4314;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4233, n53460, n53459, n53458, n53457, n53456, 
        n53455, n53454, n53453, n53452, n53451, n53450, n53449, 
        n53448, n41868, n29866, n30889, n53434, n53433, n53432, 
        n53431, n67715, n53430, n2, n67716, n53429, n67717, n53428, 
        n67681, n9_c, clk_out, n31473, n10551, n24768, n24770, 
        n24772, n15, n6, n62736, n12, n10;
    
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n29799), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_2045__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n29937), 
            .D(n37[7]), .R(n31405));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2045__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n29937), 
            .D(n37[6]), .R(n31405));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2045__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n29937), 
            .D(n37[5]), .R(n31405));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2045__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n29937), 
            .D(n37[4]), .R(n31405));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n31638));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n31637));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n31636));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n31635));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n31634));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n31633));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n31632));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n31631));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n31630));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n31629));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n31628));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12070_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29937));
    defparam i12070_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNE bit_counter_2045__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n29937), 
            .D(n24764));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2049_2050__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2051_2052__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 counter_2051_2052_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n53460), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2051_2052_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2051_2052_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n53459), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2051_2052_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2051_2052_add_4_3 (.CI(n53459), .I0(GND_net), .I1(counter[1]), 
            .CO(n53460));
    SB_LUT4 counter_2051_2052_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2051_2052_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2051_2052_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n53459));
    SB_LUT4 delay_counter_2049_2050_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n53458), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2049_2050_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n53457), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_12 (.CI(n53457), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n53458));
    SB_LUT4 delay_counter_2049_2050_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n53456), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_11 (.CI(n53456), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n53457));
    SB_LUT4 delay_counter_2049_2050_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n53455), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_10 (.CI(n53455), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n53456));
    SB_LUT4 delay_counter_2049_2050_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n53454), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_9 (.CI(n53454), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n53455));
    SB_LUT4 delay_counter_2049_2050_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n53453), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_8 (.CI(n53453), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n53454));
    SB_LUT4 delay_counter_2049_2050_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n53452), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_7 (.CI(n53452), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n53453));
    SB_LUT4 delay_counter_2049_2050_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n53451), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_6 (.CI(n53451), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n53452));
    SB_LUT4 delay_counter_2049_2050_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n53450), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_5 (.CI(n53450), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n53451));
    SB_LUT4 delay_counter_2049_2050_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n53449), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_4 (.CI(n53449), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n53450));
    SB_LUT4 delay_counter_2049_2050_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n53448), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_3 (.CI(n53448), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n53449));
    SB_LUT4 delay_counter_2049_2050_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2049_2050_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2049_2050_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n53448));
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n29866), .D(n41868), 
            .S(n30889));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_2045_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n53434), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2045_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n53433), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2045_add_4_8 (.CI(n53433), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n53434));
    SB_LUT4 bit_counter_2045_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n53432), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2045_add_4_7 (.CI(n53432), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n53433));
    SB_LUT4 bit_counter_2045_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n53431), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2045_add_4_6 (.CI(n53431), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n53432));
    SB_LUT4 bit_counter_2045_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n53430), .O(n67715)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2045_add_4_5 (.CI(n53430), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n53431));
    SB_LUT4 bit_counter_2045_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n53429), .O(n67716)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2045_add_4_4 (.CI(n53429), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n53430));
    SB_LUT4 bit_counter_2045_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n53428), .O(n67717)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2045_add_4_3 (.CI(n53428), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n53429));
    SB_LUT4 bit_counter_2045_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n67681)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2045_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2045_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n53428));
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9_c));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n31473));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n31471));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n32396));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n32395));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n32394));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n32393));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n32392));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n32391));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n32390));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n32389));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n32388));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n32387));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n32386));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n32385));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n32384));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n32101));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i51674_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n29799));
    defparam i51674_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2247_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2247_1_lut.LUT_INIT = 16'h5555;
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n29866), .D(n10551), 
            .R(n30889));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2045__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n29937), 
            .D(n24768));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2045__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n29937), 
            .D(n24770));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2045__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n29937), 
            .D(n24772));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2049_2050__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2049_2050__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2051_2052__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2051_2052__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i2183_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2183_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n27661));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_991 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n27667));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_991.LUT_INIT = 16'hffbf;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_992 (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n27680));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_992.LUT_INIT = 16'hfeff;
    SB_LUT4 i7076_3_lut (.I0(state[0]), .I1(n67715), .I2(state[1]), .I3(GND_net), 
            .O(n24772));   // verilog/tli4970.v(55[24:39])
    defparam i7076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7074_3_lut (.I0(state[0]), .I1(n67716), .I2(state[1]), .I3(GND_net), 
            .O(n24770));   // verilog/tli4970.v(55[24:39])
    defparam i7074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7072_3_lut (.I0(state[0]), .I1(n67717), .I2(state[1]), .I3(GND_net), 
            .O(n24768));   // verilog/tli4970.v(55[24:39])
    defparam i7072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2157_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n10551));
    defparam mux_2157_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n27643));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i23681_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n41527));
    defparam i23681_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2525_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2525_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), .I3(delay_counter_15__N_4314), 
            .O(n29866));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i12944_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(delay_counter_15__N_4314), .O(n30889));
    defparam i12944_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_LUT4 i13460_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31405));   // verilog/tli4970.v(55[24:39])
    defparam i13460_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 equal_268_i9_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/tli4970.v(56[12:26])
    defparam equal_268_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51690_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n41868));
    defparam i51690_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i13528_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n31473));
    defparam i13528_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i51886_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9_c));
    defparam i51886_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i2_3_lut (.I0(delay_counter[1]), .I1(delay_counter[4]), .I2(delay_counter[3]), 
            .I3(GND_net), .O(n62736));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2184_4_lut (.I0(delay_counter[0]), .I1(delay_counter[5]), .I2(delay_counter[2]), 
            .I3(n62736), .O(n12));
    defparam i2184_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_993 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_993.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i7069_3_lut (.I0(state[0]), .I1(n67681), .I2(state[1]), .I3(GND_net), 
            .O(n24764));   // verilog/tli4970.v(55[24:39])
    defparam i7069_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2889, pwm_out, clk32MHz, reset, GND_net, \pwm_counter[6] , 
            \pwm_counter[8] , VCC_net, pwm_setpoint, n17, n13) /* synthesis syn_module_defined=1 */ ;
    input n2889;
    output pwm_out;
    input clk32MHz;
    input reset;
    input GND_net;
    output \pwm_counter[6] ;
    output \pwm_counter[8] ;
    input VCC_net;
    input [23:0]pwm_setpoint;
    input n17;
    input n13;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577, n59454;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n58260, n53365, n48, n58300, n53364, n58332, n53363, 
        n58372, n53362, n58412, n53361, n58452, n53360, n58486, 
        n53359, n58530, n53358, n58580, n53357, n58630, n53356, 
        n58666, n53355, n58712, n53354, n58758, n53353, n59460, 
        n59462, n59464, n59326, n59128, n58994, n58948, n58896, 
        n58854, n58802, n53352, n53351, n53350, n53349, n53348, 
        n53347, n53346, n53345, n53344, n53343, n41, n39, n45, 
        n43, n37, n23, n25, n29, n31, n35, n11, n15, n27, 
        n9, n19, n21, n33, n68266, n68186, n12, n30, n68357, 
        n69349, n69337, n70533, n69860, n70695, n6, n69904, n69905, 
        n16, n24, n68124, n8, n68105, n69762, n68930, n4, n69908, 
        n69909, n68156, n10, n68153, n70665, n68928, n70837, n70838, 
        n70747, n68128, n70427, n70112, n70675, n62218, n22, n15_adj_5015, 
        n20, n24_adj_5016, n19_adj_5017;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2889), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_DFFR pwm_counter_2041__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n59454), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2041_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n53365), .O(n58260)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2041_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n53364), .O(n58300)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_24 (.CI(n53364), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n53365));
    SB_LUT4 pwm_counter_2041_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n53363), .O(n58332)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_23 (.CI(n53363), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n53364));
    SB_LUT4 pwm_counter_2041_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n53362), .O(n58372)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_22 (.CI(n53362), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n53363));
    SB_LUT4 pwm_counter_2041_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n53361), .O(n58412)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_21 (.CI(n53361), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n53362));
    SB_LUT4 pwm_counter_2041_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n53360), .O(n58452)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_20 (.CI(n53360), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n53361));
    SB_LUT4 pwm_counter_2041_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n53359), .O(n58486)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_19 (.CI(n53359), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n53360));
    SB_LUT4 pwm_counter_2041_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n53358), .O(n58530)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_18 (.CI(n53358), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n53359));
    SB_LUT4 pwm_counter_2041_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n53357), .O(n58580)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_17 (.CI(n53357), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n53358));
    SB_LUT4 pwm_counter_2041_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n53356), .O(n58630)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_16 (.CI(n53356), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n53357));
    SB_LUT4 pwm_counter_2041_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n53355), .O(n58666)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_15 (.CI(n53355), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n53356));
    SB_LUT4 pwm_counter_2041_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n53354), .O(n58712)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_14 (.CI(n53354), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n53355));
    SB_LUT4 pwm_counter_2041_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n53353), .O(n58758)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_13 (.CI(n53353), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n53354));
    SB_DFFR pwm_counter_2041__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n59460), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n59462), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n59464), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n59326), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n59128), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i6 (.Q(\pwm_counter[6] ), .C(clk32MHz), .D(n58994), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n58948), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i8 (.Q(\pwm_counter[8] ), .C(clk32MHz), .D(n58896), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n58854), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n58802), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n58758), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n58712), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n58666), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n58630), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n58580), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n58530), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n58486), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n58452), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n58412), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n58372), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n58332), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n58300), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2041__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n58260), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2041_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n53352), .O(n58802)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_12 (.CI(n53352), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n53353));
    SB_LUT4 pwm_counter_2041_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n53351), .O(n58854)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_11 (.CI(n53351), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n53352));
    SB_LUT4 pwm_counter_2041_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[8] ), 
            .I3(n53350), .O(n58896)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_10 (.CI(n53350), .I0(GND_net), .I1(\pwm_counter[8] ), 
            .CO(n53351));
    SB_LUT4 pwm_counter_2041_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n53349), .O(n58948)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_9 (.CI(n53349), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n53350));
    SB_LUT4 pwm_counter_2041_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[6] ), 
            .I3(n53348), .O(n58994)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_8 (.CI(n53348), .I0(GND_net), .I1(\pwm_counter[6] ), 
            .CO(n53349));
    SB_LUT4 pwm_counter_2041_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n53347), .O(n59128)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_7 (.CI(n53347), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n53348));
    SB_LUT4 pwm_counter_2041_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n53346), .O(n59326)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_6 (.CI(n53346), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n53347));
    SB_LUT4 pwm_counter_2041_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n53345), .O(n59464)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_5 (.CI(n53345), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n53346));
    SB_LUT4 pwm_counter_2041_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n53344), .O(n59462)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_4 (.CI(n53344), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n53345));
    SB_LUT4 pwm_counter_2041_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n53343), .O(n59460)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_3 (.CI(n53343), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n53344));
    SB_LUT4 pwm_counter_2041_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n59454)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2041_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n53343));
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48996_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n68266));
    defparam i48996_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48916_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n68186));
    defparam i48916_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50079_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n68357), 
            .O(n69349));
    defparam i50079_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50067_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n69349), 
            .O(n69337));
    defparam i50067_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51263_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n69337), 
            .O(n70533));
    defparam i51263_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50590_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n70533), 
            .O(n69860));
    defparam i50590_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51425_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69860), 
            .O(n70695));
    defparam i51425_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50634_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n69904));   // verilog/pwm.v(21[8:24])
    defparam i50634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50635_3_lut (.I0(n69904), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n69905));   // verilog/pwm.v(21[8:24])
    defparam i50635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48854_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n68266), 
            .O(n68124));
    defparam i48854_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50492_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n68105), 
            .O(n69762));   // verilog/pwm.v(21[8:24])
    defparam i50492_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49660_3_lut (.I0(n69905), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n68930));   // verilog/pwm.v(21[8:24])
    defparam i49660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50638_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n69908));   // verilog/pwm.v(21[8:24])
    defparam i50638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50639_3_lut (.I0(n69908), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n69909));   // verilog/pwm.v(21[8:24])
    defparam i50639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48886_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n68186), 
            .O(n68156));
    defparam i48886_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51395_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n68153), 
            .O(n70665));   // verilog/pwm.v(21[8:24])
    defparam i51395_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49658_3_lut (.I0(n69909), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n68928));   // verilog/pwm.v(21[8:24])
    defparam i49658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51567_4_lut (.I0(n68928), .I1(n70665), .I2(n35), .I3(n68156), 
            .O(n70837));   // verilog/pwm.v(21[8:24])
    defparam i51567_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51568_3_lut (.I0(n70837), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n70838));   // verilog/pwm.v(21[8:24])
    defparam i51568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51477_3_lut (.I0(n70838), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n70747));   // verilog/pwm.v(21[8:24])
    defparam i51477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48858_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n70695), 
            .O(n68128));
    defparam i48858_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51157_4_lut (.I0(n68930), .I1(n69762), .I2(n45), .I3(n68124), 
            .O(n70427));   // verilog/pwm.v(21[8:24])
    defparam i51157_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50842_3_lut (.I0(n70747), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n70112));   // verilog/pwm.v(21[8:24])
    defparam i50842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51405_4_lut (.I0(n70112), .I1(n70427), .I2(n45), .I3(n68128), 
            .O(n70675));   // verilog/pwm.v(21[8:24])
    defparam i51405_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51406_3_lut (.I0(n70675), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i51406_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(\pwm_counter[8] ), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48835_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n68105));
    defparam i48835_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(\pwm_counter[6] ), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48883_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n68153));
    defparam i48883_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(\pwm_counter[6] ), .I1(\pwm_counter[8] ), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n62218));   // verilog/pwm.v(17[20:33])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[20]), .I1(pwm_counter[19]), .I2(pwm_counter[16]), 
            .I3(pwm_counter[13]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n62218), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_5015));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[17]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_5015), .I1(n22), .I2(pwm_counter[22]), 
            .I3(pwm_counter[18]), .O(n24_adj_5016));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[15]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5017));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_5017), .I2(n24_adj_5016), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49087_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n68357));   // verilog/pwm.v(21[8:24])
    defparam i49087_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[8] , n335, GND_net, \Ki[9] , \Ki[10] , \Ki[11] , 
            \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , setpoint, IntegralLimit, 
            \Ki[1] , \Ki[0] , \Kp[2] , \Kp[3] , \Kp[4] , \Kp[5] , 
            \Kp[6] , \Ki[2] , control_update, duty, clk16MHz, reset, 
            \Ki[3] , \Kp[7] , \Kp[8] , \Kp[9] , \Kp[10] , \Kp[11] , 
            \Kp[12] , \Ki[4] , \Kp[13] , \Kp[14] , n8, \motor_state[9] , 
            \Kp[1] , \Kp[0] , \Ki[5] , \Kp[15] , \motor_state[8] , 
            \Ki[6] , \motor_state[7] , \Ki[7] , \motor_state[6] , \motor_state[5] , 
            \motor_state[4] , \motor_state[3] , \motor_state[2] , \motor_state[1] , 
            VCC_net, PWMLimit, n32332, \PID_CONTROLLER.integral , n32331, 
            n32330, n32329, n32328, n32327, n32326, n32325, n32324, 
            n32323, n32322, n32321, n32320, n32319, n32318, n32317, 
            n32316, n32315, n32314, n32313, n32312, n32311, n32308, 
            n31436, \motor_state[23] , \motor_state[22] , \motor_state[21] , 
            \motor_state[20] , \motor_state[19] , \motor_state[18] , \motor_state[17] , 
            \motor_state[16] , \motor_state[15] , \motor_state[14] , \motor_state[13] , 
            \motor_state[12] , \motor_state[11] , deadband, n41880, 
            \control_mode[7] , \control_mode[6] , \control_mode[1] , \control_mode[0] , 
            n27629, n29776, n54181, \displacement[0] , n59660, n27538, 
            n28, n31, n45, n30, n70677) /* synthesis syn_module_defined=1 */ ;
    input \Ki[8] ;
    output [23:0]n335;
    input GND_net;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]setpoint;
    input [23:0]IntegralLimit;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Ki[2] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input \Ki[3] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Ki[4] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input n8;
    input \motor_state[9] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[5] ;
    input \Kp[15] ;
    input \motor_state[8] ;
    input \Ki[6] ;
    input \motor_state[7] ;
    input \Ki[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input VCC_net;
    input [23:0]PWMLimit;
    input n32332;
    output [23:0]\PID_CONTROLLER.integral ;
    input n32331;
    input n32330;
    input n32329;
    input n32328;
    input n32327;
    input n32326;
    input n32325;
    input n32324;
    input n32323;
    input n32322;
    input n32321;
    input n32320;
    input n32319;
    input n32318;
    input n32317;
    input n32316;
    input n32315;
    input n32314;
    input n32313;
    input n32312;
    input n32311;
    input n32308;
    input n31436;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input [23:0]deadband;
    output n41880;
    input \control_mode[7] ;
    input \control_mode[6] ;
    input \control_mode[1] ;
    input \control_mode[0] ;
    input n27629;
    output n29776;
    input n54181;
    input \displacement[0] ;
    input n59660;
    input n27538;
    output n28;
    input n31;
    input n45;
    input n30;
    output n70677;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n603;
    wire [18:0]n15513;
    wire [17:0]n16781;
    
    wire n670, n52966, n676, n52967, n749, n597, n52965, n53627;
    wire [17:0]n17167;
    
    wire n743, n53628, n822, n895, n40, n70137, n45_c, n67839, 
        n70453, n524, n52964;
    wire [18:0]n15960;
    
    wire n670_adj_4448, n53626, n968, n451, n52963, n378, n52962, 
        n305, n52961, n1041, n1114, n4;
    wire [23:0]n455;
    wire [23:0]n535;
    
    wire n62410, n7071, n4751, n27540, n9980, n67803, n71680, 
        n71683;
    wire [23:0]n233;
    wire [23:0]n285;
    
    wire n284;
    wire [23:0]n310;
    
    wire n258, n98, n67801, n71674, n89, n71677, n29, n20;
    wire [23:0]n207;
    
    wire n174, n247, n320, n67800, n71668, n71671, n232, n52960, 
        n597_adj_4449, n53625, n524_adj_4450, n53624, n451_adj_4451, 
        n53623, n159, n52959, n378_adj_4452, n53622, n17, n86, 
        n305_adj_4453, n53621, n232_adj_4454, n53620, n67799, n71662, 
        n159_adj_4455, n53619;
    wire [16:0]n17907;
    
    wire n52958, n52957, n71665, n17_adj_4456, n86_adj_4457, n52956, 
        n393, n466, n162, n1111, n52955, n67798, n71656, n1038, 
        n52954, n71659, n965, n52953, n892, n52952, n819, n52951, 
        n746, n52950, n71647, counter_31__N_3714, n673, n52949, 
        n600, n52948, n67797, n71650, n71653, n527, n52947, n67796, 
        n71644, n454, n52946, n381, n52945, n308, n52944, n235, 
        n52943, n171, n244, n539, n612, n685, n52942;
    wire [15:0]n18896;
    
    wire n52941, n52940, n758, n831, n904, n317, n977, n1050, 
        n52939, n52938, n52570, n52571, n52937, n52569, n52936, 
        n52935, n52934, n98_adj_4458, n52933, n29_adj_4459, n171_adj_4460, 
        n52932, n244_adj_4461, n317_adj_4462, n530, n52931, n390, 
        n457, n52930, n463, n536_adj_4463, n609, n682, n755, n828, 
        n901, n384, n52929, n974, n390_adj_4464, n1047, n1120, 
        n52568, n311, n52928, n95, n238, n52927, n26, n165, 
        n52926, n23, n92;
    wire [8:0]n22573;
    wire [7:0]n22752;
    
    wire n700, n52925, n463_adj_4465, n168, n241, n314, n627, 
        n52924, n52567, n387, n536_adj_4466, n460, n533, n606, 
        n554_adj_4467, n52923, n679, n752, n481, n52922, n408, 
        n52921, n609_adj_4468, n335_c, n52920, n262, n52919, n682_adj_4469, 
        n755_adj_4470, n825, n898, n971, n189, n52918, n1044, 
        n828_adj_4471, n47, n116;
    wire [14:0]n19756;
    
    wire n52917, n1117, n52916, n52566, n1117_adj_4472, n92_adj_4473, 
        n1044_adj_4474, n52915, n971_adj_4475, n52914, n898_adj_4476, 
        n52913, n23_adj_4477;
    wire [16:0]n18235;
    
    wire n53598, n825_adj_4478, n52912, n53597, n752_adj_4479, n52911, 
        n165_adj_4480, n679_adj_4481, n52910, n901_adj_4482, n606_adj_4483, 
        n52909, n53596, n533_adj_4484, n52908, n1111_adj_4485, n53595, 
        n238_adj_4486, n1038_adj_4487, n53594, n965_adj_4488, n53593, 
        n892_adj_4489, n53592, n819_adj_4490, n53591, n746_adj_4491, 
        n53590, n673_adj_4492, n53589, n600_adj_4493, n53588, n311_adj_4494, 
        n384_adj_4495, n457_adj_4496, n974_adj_4497, n527_adj_4498, 
        n53587, n454_adj_4499, n53586, n460_adj_4500, n52907, n381_adj_4501, 
        n53585, n308_adj_4502, n53584, n387_adj_4503, n52906, n235_adj_4504, 
        n53583, n162_adj_4505, n53582, n20_adj_4506, n89_adj_4507, 
        n314_adj_4508, n52905;
    wire [15:0]n19169;
    
    wire n53581, n241_adj_4509, n52904, n53580, n1114_adj_4510, n53579, 
        n52565, n1041_adj_4511, n53578, n968_adj_4512, n53577, n895_adj_4513, 
        n53576, n822_adj_4514, n53575, n168_adj_4515, n52903, n1047_adj_4516, 
        n1120_adj_4517, n26_adj_4518, n95_adj_4519, n749_adj_4520, n53574, 
        n52564, n676_adj_4521, n53573, n603_adj_4522, n53572, n530_adj_4523, 
        n53571, n52563;
    wire [13:0]n20475;
    
    wire n52902, n52901, n52900, n53570, n53569, n53568, n53567, 
        n52899, n53566;
    wire [14:0]n19977;
    
    wire n53565, n53564, n52898, n53563, n53562, n53561, n53560, 
        n52897, n52896, n52895, n53559, n53558, n53557, n53556, 
        n53555, n52894, n53554, n53553, n53552, n53551, n52893;
    wire [13:0]n20667;
    
    wire n53550, n53549, n52892, n53548, n53547, n53546, n53545, 
        n53544, n53543, n53542, n53541, n53540, n53539, n53538, 
        n53537;
    wire [12:0]n21245;
    
    wire n53536, n53535, n52891, n53534, n53533, n53532, n53531, 
        n53530, n53529, n52890, n52889, n53528, n53527, n53526, 
        n53525, n53524;
    wire [12:0]n21080;
    
    wire n1050_adj_4524, n52888, n32, n101, n977_adj_4525, n52887;
    wire [11:0]n21718;
    
    wire n980, n53523, n907, n53522, n834, n53521, n761, n53520, 
        n688, n53519, n615, n53518, n904_adj_4526, n52886, n542, 
        n53517, n469, n53516, n396, n53515, n831_adj_4527, n52885, 
        n323, n53514, n758_adj_4528, n52884, n250, n53513, n177, 
        n53512, n685_adj_4529, n52883, n35, n104, n612_adj_4530, 
        n52882, n539_adj_4531, n52881, n466_adj_4532, n52880, n393_adj_4533, 
        n52879, n320_adj_4534, n52878, n52562, n247_adj_4535, n52877, 
        n174_adj_4536, n52876, n52561;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n32_adj_4537, n101_adj_4538;
    wire [6:0]n22878;
    
    wire n630, n52875, n557_adj_4539, n52874, n484, n52873, n411, 
        n52872, n338, n52871;
    wire [10:0]n22091;
    wire [9:0]n22374;
    
    wire n840, n53116, n767, n53115, n694, n53114, n265, n52870, 
        n621, n53113;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n71491, n548, n53112, n192, n52869, n475_adj_4540, n53111, 
        n402, n53110, n50, n119, n329, n53109, n256, n53108;
    wire [11:0]n21578;
    
    wire n980_adj_4541, n52868, n907_adj_4542, n52867, n183, n53107, 
        n41, n110, n834_adj_4543, n52866, n761_adj_4544, n52865, 
        n688_adj_4545, n52864;
    wire [5:0]n22974;
    
    wire n61693, n490, n53906;
    wire [4:0]n23044;
    
    wire n417, n53905, n344, n53904, n53447, n271, n53903, n53446, 
        n198, n53902, n53445, n56, n125, n53444;
    wire [8:0]n22496;
    wire [7:0]n22692;
    
    wire n700_adj_4546, n53901, n627_adj_4547, n53900, n554_adj_4548, 
        n53899, n615_adj_4549, n52863, n53443, n542_adj_4550, n52862, 
        n481_adj_4551, n53898, n469_adj_4552, n52861, n396_adj_4553, 
        n52860, n323_adj_4554, n52859, n250_adj_4555, n52858, n408_adj_4556, 
        n53897, n53442, n335_adj_4557, n53896, n53441, n262_adj_4558, 
        n53895, n53440, n177_adj_4559, n52857, n189_adj_4560, n53894, 
        n47_adj_4561, n116_adj_4562, n35_adj_4563, n104_adj_4564, n53439;
    wire [10:0]n21974;
    
    wire n910, n52856;
    wire [6:0]n22833;
    
    wire n630_adj_4565, n53893, n53438, n837, n52855, n557_adj_4566, 
        n53892, n484_adj_4567, n53891, n764, n52854, n53437, n411_adj_4568, 
        n53890, n53436, n338_adj_4569, n53889, n53435, n265_adj_4570, 
        n53888, n192_adj_4571, n53887, n691, n52853, n50_adj_4572, 
        n119_adj_4573, n71311, n618, n52852, n545, n52851, n71293, 
        n71287, n71281, n71275, n71269, n71263, n71257, n71251, 
        n71245, n71239, n71233, n71227, n71221, n71215, n71209, 
        n472, n52850, n399, n52849, n326_adj_4574, n52848, n67744, 
        n71488, n253, n52847, n180, n52846, n38, n107, n560, 
        n52845, n487, n52844, n414, n52843, n341, n52842, n268, 
        n52841, n195, n52840, n53, n122;
    wire [9:0]n22278;
    
    wire n840_adj_4575, n52839, n767_adj_4576, n52838, n694_adj_4577, 
        n52837, n621_adj_4578, n52836, n548_adj_4579, n52835, n70449, 
        n27506, n27508, n475_adj_4581, n52834, n402_adj_4582, n52833, 
        n329_adj_4583, n52832, n256_adj_4584, n52831, n183_adj_4585, 
        n52830, n41_adj_4586, n110_adj_4587, n770, n52829, n697, 
        n52828, n624, n52827, n68118, n551, n52826, n6, n478_adj_4588, 
        n52825;
    wire [0:0]n10812;
    wire [0:0]n10020;
    
    wire n52629, n405, n52824, n332, n52823, n259, n52822;
    wire [43:0]n360;
    wire [47:0]n36;
    
    wire n52628, n186, n52821, n44, n113, n52627, n52626, n52625;
    wire [5:0]n22942;
    
    wire n560_adj_4592, n53773, n487_adj_4593, n53772, n52624, n414_adj_4594, 
        n53771, n52623, n341_adj_4596, n53770, n268_adj_4597, n53769, 
        n195_adj_4598, n53768, n53_adj_4599, n122_adj_4600, n52622, 
        n52621, n52620, n52619, n52618, n52617, n52616, n910_adj_4606, 
        n53325, n837_adj_4607, n53324, n764_adj_4608, n53323, n52615, 
        n691_adj_4609, n53322, n618_adj_4610, n53321, n545_adj_4611, 
        n53320, n52614, n472_adj_4613, n53319, n770_adj_4614, n53067, 
        n697_adj_4615, n53066, n399_adj_4616, n53318, n326_adj_4617, 
        n53317, n62793, n490_adj_4618, n53744;
    wire [4:0]n23023;
    
    wire n417_adj_4619, n53743, n253_adj_4620, n53316, n344_adj_4621, 
        n53742, n180_adj_4622, n53315, n271_adj_4623, n53741, n38_adj_4624, 
        n107_adj_4625, n52613, n198_adj_4627, n53740, n56_adj_4628, 
        n125_adj_4629;
    wire [21:0]n11271;
    
    wire n53739, n53738, n624_adj_4630, n53065, n53737, n52612, 
        n551_adj_4631, n53064, n53736, n53735, n53734, n53733, n53732, 
        n1096, n53731, n1023, n53730, n950, n53729, n478_adj_4632, 
        n53063, n877, n53728, n804, n53727, n52611, n405_adj_4634, 
        n53062, n731, n53726, n52610, n658, n53725, n585, n53724, 
        n52609, n512, n53723, n332_adj_4635, n53061, n259_adj_4636, 
        n53060, n439_adj_4637, n53722, n366, n53721, n293, n53720, 
        n220_adj_4638, n53719, n186_adj_4639, n53059, n147, n53718, 
        n5, n74_adj_4641;
    wire [20:0]n13100;
    
    wire n53696, n44_adj_4642, n113_adj_4643;
    wire [21:0]n10527;
    
    wire n53058, n53695, n53057, n53056, n53055, n53694, n53054, 
        n53053, n53693, n53052, n52608, n53051, n52607, n1096_adj_4645, 
        n53050, n53692;
    wire [23:0]n1_adj_5012;
    
    wire n52775, n1023_adj_4646, n53049, n52774, n53691, n53690, 
        n950_adj_4647, n53048, n52773, n877_adj_4649, n53047, n52772, 
        n1099, n53689, n804_adj_4652, n53046, n52771, n52606, n52605, 
        n52770, n731_adj_4655, n53045, n52769, n52604, n658_adj_4658, 
        n53044, n52768, n585_adj_4659, n53043, n1026, n53688, n512_adj_4660, 
        n53042, n439_adj_4661, n53041, n52767, n953, n53687, n366_adj_4662, 
        n53040, n293_adj_4663, n53039, n52766, n52765, n220_adj_4665, 
        n53038, n52603, n880, n53686, n52764, n52602, n147_adj_4667, 
        n53037, n52763, n52762, n52601, n52600, n807, n53685, 
        n5_adj_4669, n74_adj_4670, n52761, n734, n53684;
    wire [20:0]n12521;
    
    wire n53036, n52760, n53035, n52759, n661, n53683, n53034, 
        n52758, n53033, n588, n53682, n52757, n52756, n52599, 
        n52598, n515, n53681, n53032, n52755, n53031, n52754, 
        n442_adj_4676, n53680, n52753, n53030, n52597, n369, n53679, 
        n1099_adj_4677, n53029, n47_adj_4678;
    wire [23:0]n1_adj_5013;
    
    wire n52752;
    wire [23:0]n46;
    
    wire n52751, n1026_adj_4681, n53028, n52750, n296, n53678, n953_adj_4684, 
        n53027, n52749, n223_adj_4686, n53677, n880_adj_4687, n53026, 
        n52748, n150, n53676, n807_adj_4689, n53025, n52747, n52596, 
        n734_adj_4693, n53024, n52746, n52595, n52594, n661_adj_4695, 
        n53023, n52745, n588_adj_4697, n53022, n52744, n52743, n8_adj_4701, 
        n77, n515_adj_4702, n53021, n52742, n442_adj_4704, n53020, 
        n52741;
    wire [19:0]n14607;
    
    wire n53675, n369_adj_4706, n53019, n52740, n53674, n296_adj_4708, 
        n53018, n52739, n52593, n53673, n223_adj_4710, n53017, n52738, 
        n52592, n150_adj_4712, n53016, n52737, n52591, n8_adj_4714, 
        n77_adj_4715, n52736, n53672, n52735;
    wire [19:0]n14096;
    
    wire n53015, n53671, n53014, n52734, n53013, n52733, n53670, 
        n53012, n52732, n1102, n53669, n53011, n52590, n67600, 
        n71308, n52589, n53010, n52731, n1029, n53668, n1102_adj_4723, 
        n53009, n52730, n67612, n41898, n1029_adj_4726, n53008;
    wire [23:0]n1_adj_5014;
    
    wire n52729, n52728, n956, n53667, n883, n53666, n956_adj_4729, 
        n53007, n52727, n52588, n883_adj_4731, n53006, n52726, n52725, 
        n52587, n810, n53005, n52724, n52723, n810_adj_4737, n53665, 
        n737, n53004, n52722, n52586, n52721, n52585, n664, n53003, 
        n52720, n52719, n52584, n737_adj_4745, n53664, n591, n53002, 
        n52718, n52717, n518, n53001, n664_adj_4748, n53663, n445_adj_4749, 
        n53000, n372, n52999, n591_adj_4750, n53662, n299_adj_4751, 
        n52998, n518_adj_4752, n53661, n226_adj_4753, n52997, n52716, 
        n52715, n153, n52996, n52714, n52583, n52582, n11_adj_4757, 
        n80, n52713, n445_adj_4759, n53660, n52995, n52994, n52712, 
        n52581, n372_adj_4761, n53659, n52580, n52711, n52579, n52993, 
        n52710, n52992, n299_adj_4765, n53658, n52991, n1105, n52990, 
        n52578, n52709, n52577, n1032, n52989, n226_adj_4767, n53657, 
        n52708, n52576, n153_adj_4769, n53656, n959, n52988, n886, 
        n52987, n11_adj_4770, n80_adj_4771, n52707, n52575, n813, 
        n52986, n53655, n740, n52985, n53654, n667, n52984, n52574, 
        n53653, n594, n52983, n52573, n521, n52982, n448_adj_4775, 
        n52981, n53652, n375, n52980, n52572, n53651, n302_adj_4776, 
        n52979, n229, n52978, n156, n52977, n1105_adj_4777, n53650, 
        n14_adj_4778, n83, n1032_adj_4779, n53649, n52976, n959_adj_4780, 
        n53648, n886_adj_4781, n53647, n52975, n52974, n52973, n813_adj_4782, 
        n53646, n1108, n52972, n740_adj_4783, n53645, n1035, n52971, 
        n962, n52970, n667_adj_4784, n53644, n889, n52969, n594_adj_4785, 
        n53643, n521_adj_4786, n53642, n448_adj_4787, n53641, n375_adj_4788, 
        n53640, n302_adj_4789, n53639, n229_adj_4790, n53638, n816, 
        n52968, n156_adj_4791, n53637, n743_adj_4792, n14_adj_4793, 
        n83_adj_4794, n53636, n53635, n53634, n53633, n1108_adj_4795, 
        n53632, n1035_adj_4796, n53631, n962_adj_4797, n53630, n889_adj_4798, 
        n53629, n816_adj_4799, n9_adj_4800, n11_adj_4801, n13_adj_4802, 
        n15_adj_4803, n21_adj_4804, n19_adj_4805, n17_adj_4806, n23_adj_4807, 
        n25_adj_4808, n9_adj_4809, n11_adj_4810, n13_adj_4811, n15_adj_4812, 
        n64295, n67833, n23_adj_4813, n21_adj_4814, n19_adj_4815, 
        n17_adj_4816, n23_adj_4817, n22_adj_4818, n25_adj_4819, n27, 
        n26_adj_4820, n67845, n67934, n68007, n45_adj_4821, n41_adj_4822, 
        n43, n37, n39, n33, n31_c, n27_adj_4823, n35_adj_4824, 
        n29_adj_4825, n68460, n68447, n68231, n12_adj_4826, n68264, 
        n68309, n27602;
    wire [3:0]n23080;
    
    wire n6_adj_4828, n32_adj_4829, n204, n68604, n34;
    wire [1:0]n23138;
    
    wire n52254;
    wire [2:0]n23117;
    
    wire n131, n62_adj_4830, n68761, n10_adj_4831, n6_adj_4832, n68697, 
        n8_adj_4833, n10_adj_4834, n68343, n30_c, n53911, n52279, 
        n63933, n63937, n63935, n52224, n63943, n4_adj_4836, n8_adj_4837, 
        n6_adj_4838, n68482, n68521, n68478, n69469, n69461, n70577, 
        n69984, n70716, n16_adj_4839, n6_adj_4840, n70274, n70275, 
        n8_adj_4841, n24_adj_4842, n68417, n68411, n69782, n68964, 
        n68435, n4_adj_4843, n70270, n70271, n68441, n70593, n68966, 
        n70805, n70806, n70792, n68421, n70437, n68972, n39_adj_4849, 
        n41_adj_4850, n45_adj_4851, n43_adj_4852, n29_adj_4853, n31_adj_4854, 
        n37_adj_4855, n23_adj_4856, n25_adj_4857, n35_adj_4858, n41540, 
        n41850, n11_adj_4859, n13_adj_4860, n68307, n6_adj_4861, n7073, 
        n67557, n27_adj_4862, n67558, n67559, n67563, n9_adj_4863, 
        n67564, n67565, n67566, n67567, n17_adj_4864, n67568, n19_adj_4865, 
        n21_adj_4866, n15_adj_4867, n33_adj_4868, n70681, n68573, 
        n68548, n12_adj_4869, n10_adj_4870, n30_adj_4871, n67593, 
        n67587, n67584, n67569, n67570, n67575, n67926, n68596, 
        n69569, n6_adj_4872, n69555, n70619, n70024, n68_adj_4874, 
        n63987, n70734, n16_adj_4875, n6_adj_4876, n70284, n70285, 
        n70679, n8_adj_4877, n24_adj_4878, n68484, n69780, n68954, 
        n4_adj_4879, n70280, n70281, n68527, n70591, n45_adj_4880, 
        n71290, n68956, n70803, n39_adj_4882, n70804, n70794, n68487, 
        n70435, n68962, n41_adj_4883, n43_adj_4884, n41_adj_4885, 
        n37_adj_4886, n39_adj_4887, n43_adj_4888, n31_adj_4889, n29_adj_4891, 
        n31_adj_4892, n33_adj_4893, n37_adj_4894, n17_adj_4895, n19_adj_4896, 
        n21_adj_4897, n23_adj_4898, n25_adj_4899, n52284, n9_adj_4900, 
        n29_adj_4901, n35_adj_4902, n71284, n33_adj_4903;
    wire [3:0]n23092;
    
    wire n4_adj_4904, n35_adj_4905, n347_adj_4906, n6_adj_4907, n60085, 
        n11_adj_4908, n13_adj_4909, n63983, n68375, n63973, n72161, 
        n63977, n8_adj_4910, n6_adj_4911, n15_adj_4912, n27_adj_4913, 
        n41_adj_4914, n68359, n39_adj_4915, n15_adj_4916, n13_adj_4917, 
        n19_adj_4918, n12_adj_4919, n17_adj_4920, n7_adj_4921, n9_adj_4922, 
        n11_adj_4923, n5_adj_4924, n68763, n71278, n16_adj_4925, n4_adj_4926, 
        n12_adj_4927, n68755, n70589, n69778, n70844, n70845, n70739, 
        n70125, n10_adj_4928, n33_adj_4929, n30_adj_4930, n35_adj_4931, 
        n37_adj_4932, n43_adj_4933, n68623, n42, n70286, n70287, 
        n68608, n70127, n68952, n105, n41_adj_4937, n39_adj_4938, 
        n45_adj_4939, n29_adj_4940, n31_adj_4941, n43_adj_4942, n37_adj_4943, 
        n17_adj_4944, n19_adj_4945, n21_adj_4946, n71272, n23_adj_4947, 
        n25_adj_4948, n9_adj_4949, n35_adj_4950, n68409, n69403, n33_adj_4951, 
        n11_adj_4952, n13_adj_4953, n15_adj_4954, n27_adj_4955, n69387, 
        n68220, n69243, n71827, n69209, n71822, n68209, n69235, 
        n71842, n69229, n71837, n70563, n16_adj_4956, n68120, n8_adj_4957, 
        n24_adj_4958, n69948, n68229, n71835, n68222, n71863, n69888, 
        n71860, n70712, n16_adj_4959, n69239, n6_adj_4960, n70266, 
        n70254, n70267, n68194, n8_adj_4961, n24_adj_4962, n71825, 
        n68315, n69862, n71854, n70509, n71816, n69784, n68974, 
        n70770, n4_adj_4963, n71813, n68278, n12_adj_4964, n10_adj_4965, 
        n70264, n30_adj_4966, n70265, n69311, n69303, n70553, n69912, 
        n70708, n16_adj_4967, n71266, n8_adj_4968, n24_adj_4969, n68351, 
        n70260, n70261, n68286, n68236, n69786, n70595, n68976, 
        n68984, n4_adj_4970, n69874, n70809, n69875, n12_adj_4971, 
        n68151, n71848, n10_adj_4972, n30_adj_4973, n68165, n70810, 
        n70790, n70362, n68996, n68319, n70718, n70439, n70719, 
        n70705, n6_adj_4974, n68982, n69878, n69879, n68122, n70683, 
        n71810, n69788, n68994, n68133, n70443, n69002, n70687, 
        n4_adj_4975, n70258, n70259, n68270, n70599, n68986, n70811, 
        n71260, n70812, n70788, n68251, n70441, n68992, n70688, 
        n70685, n4_adj_4976, n52388, n4_adj_4977, n39_adj_4978, n41_adj_4979, 
        n45_adj_4980, n43_adj_4981, n37_adj_4982, n29_adj_4983, n31_adj_4984, 
        n23_adj_4985, n25_adj_4986, n35_adj_4987, n33_adj_4988, n11_adj_4989, 
        n71254, n71248, n13_adj_4990, n71242, n15_adj_4991, n27_adj_4992, 
        n9_adj_4993, n17_adj_4994, n19_adj_4995, n21_adj_4996, n68072, 
        n71236, n71230, n68036, n12_adj_4997, n10_adj_4998, n30_adj_4999, 
        n69066, n69062, n70469, n71224, n69804, n70689, n16_adj_5000, 
        n69866, n71218, n69867, n8_adj_5001, n24_adj_5002, n71212, 
        n67946, n71206, n69790, n69004, n4_adj_5003, n69864, n69865, 
        n68009, n70720, n69006, n70869, n70870, n70832, n67948, 
        n70447, n40_adj_5004, n67859, n12_adj_5005, n10_adj_5006, 
        n30_adj_5007, n68889, n68883, n70415, n69720, n70671, n70360, 
        n70361, n16_adj_5008, n8_adj_5009, n24_adj_5010, n67886, n67835, 
        n69792, n70132, n4_adj_5011, n70356, n70357, n67847, n70722, 
        n70134, n70871, n70872, n70830;
    
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5097_10_lut (.I0(GND_net), .I1(n16781[7]), .I2(n670), 
            .I3(n52966), .O(n15513[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5097_10 (.CI(n52966), .I0(n16781[7]), .I1(n670), .CO(n52967));
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5097_9_lut (.I0(GND_net), .I1(n16781[6]), .I2(n597), .I3(n52965), 
            .O(n15513[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_11 (.CI(n53627), .I0(n17167[8]), .I1(n743), .CO(n53628));
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51183_4_lut (.I0(n40), .I1(n70137), .I2(n45_c), .I3(n67839), 
            .O(n70453));   // verilog/motorControl.v(65[25:41])
    defparam i51183_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5097_9 (.CI(n52965), .I0(n16781[6]), .I1(n597), .CO(n52966));
    SB_LUT4 add_5097_8_lut (.I0(GND_net), .I1(n16781[5]), .I2(n524), .I3(n52964), 
            .O(n15513[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_10_lut (.I0(GND_net), .I1(n17167[7]), .I2(n670_adj_4448), 
            .I3(n53626), .O(n15960[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_8 (.CI(n52964), .I0(n16781[5]), .I1(n524), .CO(n52965));
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5097_7_lut (.I0(GND_net), .I1(n16781[4]), .I2(n451), .I3(n52963), 
            .O(n15513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_7 (.CI(n52963), .I0(n16781[4]), .I1(n451), .CO(n52964));
    SB_LUT4 add_5097_6_lut (.I0(GND_net), .I1(n16781[3]), .I2(n378), .I3(n52962), 
            .O(n15513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_6 (.CI(n52962), .I0(n16781[3]), .I1(n378), .CO(n52963));
    SB_LUT4 add_5097_5_lut (.I0(GND_net), .I1(n16781[2]), .I2(n305), .I3(n52961), 
            .O(n15513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_5 (.CI(n52961), .I0(n16781[2]), .I1(n305), .CO(n52962));
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n70453), .I1(n4), .I2(n455[23]), .I3(n535[23]), 
            .O(n62410));
    defparam i2_4_lut.LUT_INIT = 16'hdfcd;
    SB_LUT4 i4431_4_lut (.I0(n7071), .I1(n4751), .I2(n62410), .I3(n27540), 
            .O(n9980));
    defparam i4431_4_lut.LUT_INIT = 16'hbbab;
    SB_LUT4 n9980_bdd_4_lut (.I0(n9980), .I1(n67803), .I2(setpoint[6]), 
            .I3(n4751), .O(n71680));
    defparam n9980_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71680_bdd_4_lut (.I0(n71680), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4751), .O(n71683));
    defparam n71680_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n335[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n335[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9980_bdd_4_lut_52320 (.I0(n9980), .I1(n67801), .I2(setpoint[5]), 
            .I3(n4751), .O(n71674));
    defparam n9980_bdd_4_lut_52320.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71674_bdd_4_lut (.I0(n71674), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4751), .O(n71677));
    defparam n71674_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9980_bdd_4_lut_52315 (.I0(n9980), .I1(n67800), .I2(setpoint[4]), 
            .I3(n4751), .O(n71668));
    defparam n9980_bdd_4_lut_52315.LUT_INIT = 16'he4aa;
    SB_LUT4 n71668_bdd_4_lut (.I0(n71668), .I1(n535[4]), .I2(n455[4]), 
            .I3(n4751), .O(n71671));
    defparam n71668_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5097_4_lut (.I0(GND_net), .I1(n16781[1]), .I2(n232), .I3(n52960), 
            .O(n15513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_10 (.CI(n53626), .I0(n17167[7]), .I1(n670_adj_4448), 
            .CO(n53627));
    SB_LUT4 add_5118_9_lut (.I0(GND_net), .I1(n17167[6]), .I2(n597_adj_4449), 
            .I3(n53625), .O(n15960[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_9 (.CI(n53625), .I0(n17167[6]), .I1(n597_adj_4449), 
            .CO(n53626));
    SB_LUT4 add_5118_8_lut (.I0(GND_net), .I1(n17167[5]), .I2(n524_adj_4450), 
            .I3(n53624), .O(n15960[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_8 (.CI(n53624), .I0(n17167[5]), .I1(n524_adj_4450), 
            .CO(n53625));
    SB_LUT4 add_5118_7_lut (.I0(GND_net), .I1(n17167[4]), .I2(n451_adj_4451), 
            .I3(n53623), .O(n15960[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_4 (.CI(n52960), .I0(n16781[1]), .I1(n232), .CO(n52961));
    SB_LUT4 add_5097_3_lut (.I0(GND_net), .I1(n16781[0]), .I2(n159), .I3(n52959), 
            .O(n15513[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_7 (.CI(n53623), .I0(n17167[4]), .I1(n451_adj_4451), 
            .CO(n53624));
    SB_CARRY add_5097_3 (.CI(n52959), .I0(n16781[0]), .I1(n159), .CO(n52960));
    SB_LUT4 add_5118_6_lut (.I0(GND_net), .I1(n17167[3]), .I2(n378_adj_4452), 
            .I3(n53622), .O(n15960[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_6 (.CI(n53622), .I0(n17167[3]), .I1(n378_adj_4452), 
            .CO(n53623));
    SB_LUT4 add_5097_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n15513[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_5_lut (.I0(GND_net), .I1(n17167[2]), .I2(n305_adj_4453), 
            .I3(n53621), .O(n15960[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_5 (.CI(n53621), .I0(n17167[2]), .I1(n305_adj_4453), 
            .CO(n53622));
    SB_LUT4 add_5118_4_lut (.I0(GND_net), .I1(n17167[1]), .I2(n232_adj_4454), 
            .I3(n53620), .O(n15960[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_4 (.CI(n53620), .I0(n17167[1]), .I1(n232_adj_4454), 
            .CO(n53621));
    SB_LUT4 n9980_bdd_4_lut_52310 (.I0(n9980), .I1(n67799), .I2(setpoint[3]), 
            .I3(n4751), .O(n71662));
    defparam n9980_bdd_4_lut_52310.LUT_INIT = 16'he4aa;
    SB_CARRY add_5097_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n52959));
    SB_LUT4 add_5118_3_lut (.I0(GND_net), .I1(n17167[0]), .I2(n159_adj_4455), 
            .I3(n53619), .O(n15960[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_19_lut (.I0(GND_net), .I1(n17907[16]), .I2(GND_net), 
            .I3(n52958), .O(n16781[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_18_lut (.I0(GND_net), .I1(n17907[15]), .I2(GND_net), 
            .I3(n52957), .O(n16781[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_3 (.CI(n53619), .I0(n17167[0]), .I1(n159_adj_4455), 
            .CO(n53620));
    SB_LUT4 n71662_bdd_4_lut (.I0(n71662), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4751), .O(n71665));
    defparam n71662_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5118_2_lut (.I0(GND_net), .I1(n17_adj_4456), .I2(n86_adj_4457), 
            .I3(GND_net), .O(n15960[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_2 (.CI(GND_net), .I0(n17_adj_4456), .I1(n86_adj_4457), 
            .CO(n53619));
    SB_CARRY add_5153_18 (.CI(n52957), .I0(n17907[15]), .I1(GND_net), 
            .CO(n52958));
    SB_LUT4 add_5153_17_lut (.I0(GND_net), .I1(n17907[14]), .I2(GND_net), 
            .I3(n52956), .O(n16781[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5153_17 (.CI(n52956), .I0(n17907[14]), .I1(GND_net), 
            .CO(n52957));
    SB_LUT4 add_5153_16_lut (.I0(GND_net), .I1(n17907[13]), .I2(n1111), 
            .I3(n52955), .O(n16781[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_16 (.CI(n52955), .I0(n17907[13]), .I1(n1111), .CO(n52956));
    SB_LUT4 n9980_bdd_4_lut_52305 (.I0(n9980), .I1(n67798), .I2(setpoint[2]), 
            .I3(n4751), .O(n71656));
    defparam n9980_bdd_4_lut_52305.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5153_15_lut (.I0(GND_net), .I1(n17907[12]), .I2(n1038), 
            .I3(n52954), .O(n16781[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_15 (.CI(n52954), .I0(n17907[12]), .I1(n1038), .CO(n52955));
    SB_LUT4 n71656_bdd_4_lut (.I0(n71656), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4751), .O(n71659));
    defparam n71656_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5153_14_lut (.I0(GND_net), .I1(n17907[11]), .I2(n965), 
            .I3(n52953), .O(n16781[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_14 (.CI(n52953), .I0(n17907[11]), .I1(n965), .CO(n52954));
    SB_LUT4 add_5153_13_lut (.I0(GND_net), .I1(n17907[10]), .I2(n892), 
            .I3(n52952), .O(n16781[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_13 (.CI(n52952), .I0(n17907[10]), .I1(n892), .CO(n52953));
    SB_LUT4 add_5153_12_lut (.I0(GND_net), .I1(n17907[9]), .I2(n819), 
            .I3(n52951), .O(n16781[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_12 (.CI(n52951), .I0(n17907[9]), .I1(n819), .CO(n52952));
    SB_LUT4 add_5153_11_lut (.I0(GND_net), .I1(n17907[8]), .I2(n746), 
            .I3(n52950), .O(n16781[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_11 (.CI(n52950), .I0(n17907[8]), .I1(n746), .CO(n52951));
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n71647), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_LUT4 add_5153_10_lut (.I0(GND_net), .I1(n17907[7]), .I2(n673), 
            .I3(n52949), .O(n16781[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_10 (.CI(n52949), .I0(n17907[7]), .I1(n673), .CO(n52950));
    SB_LUT4 add_5153_9_lut (.I0(GND_net), .I1(n17907[6]), .I2(n600), .I3(n52948), 
            .O(n16781[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9980_bdd_4_lut_52300 (.I0(n9980), .I1(n67797), .I2(setpoint[1]), 
            .I3(n4751), .O(n71650));
    defparam n9980_bdd_4_lut_52300.LUT_INIT = 16'he4aa;
    SB_CARRY add_5153_9 (.CI(n52948), .I0(n17907[6]), .I1(n600), .CO(n52949));
    SB_LUT4 n71650_bdd_4_lut (.I0(n71650), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4751), .O(n71653));
    defparam n71650_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5153_8_lut (.I0(GND_net), .I1(n17907[5]), .I2(n527), .I3(n52947), 
            .O(n16781[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9980_bdd_4_lut_52295 (.I0(n9980), .I1(n67796), .I2(setpoint[0]), 
            .I3(n4751), .O(n71644));
    defparam n9980_bdd_4_lut_52295.LUT_INIT = 16'he4aa;
    SB_CARRY add_5153_8 (.CI(n52947), .I0(n17907[5]), .I1(n527), .CO(n52948));
    SB_LUT4 add_5153_7_lut (.I0(GND_net), .I1(n17907[4]), .I2(n454), .I3(n52946), 
            .O(n16781[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_7 (.CI(n52946), .I0(n17907[4]), .I1(n454), .CO(n52947));
    SB_LUT4 add_5153_6_lut (.I0(GND_net), .I1(n17907[3]), .I2(n381), .I3(n52945), 
            .O(n16781[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71644_bdd_4_lut (.I0(n71644), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4751), .O(n71647));
    defparam n71644_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_5153_6 (.CI(n52945), .I0(n17907[3]), .I1(n381), .CO(n52946));
    SB_LUT4 add_5153_5_lut (.I0(GND_net), .I1(n17907[2]), .I2(n308), .I3(n52944), 
            .O(n16781[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_5 (.CI(n52944), .I0(n17907[2]), .I1(n308), .CO(n52945));
    SB_LUT4 add_5153_4_lut (.I0(GND_net), .I1(n17907[1]), .I2(n235), .I3(n52943), 
            .O(n16781[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5153_4 (.CI(n52943), .I0(n17907[1]), .I1(n235), .CO(n52944));
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5153_3_lut (.I0(GND_net), .I1(n17907[0]), .I2(n162), .I3(n52942), 
            .O(n16781[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_3 (.CI(n52942), .I0(n17907[0]), .I1(n162), .CO(n52943));
    SB_LUT4 add_5153_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n16781[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n52942));
    SB_LUT4 add_5206_18_lut (.I0(GND_net), .I1(n18896[15]), .I2(GND_net), 
            .I3(n52941), .O(n17907[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5206_17_lut (.I0(GND_net), .I1(n18896[14]), .I2(GND_net), 
            .I3(n52940), .O(n17907[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5206_17 (.CI(n52940), .I0(n18896[14]), .I1(GND_net), 
            .CO(n52941));
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5206_16_lut (.I0(GND_net), .I1(n18896[13]), .I2(n1114), 
            .I3(n52939), .O(n17907[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_16 (.CI(n52939), .I0(n18896[13]), .I1(n1114), .CO(n52940));
    SB_LUT4 add_5206_15_lut (.I0(GND_net), .I1(n18896[12]), .I2(n1041), 
            .I3(n52938), .O(n17907[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_15 (.CI(n52938), .I0(n18896[12]), .I1(n1041), .CO(n52939));
    SB_CARRY sub_15_add_2_12 (.CI(n52570), .I0(setpoint[10]), .I1(n8), 
            .CO(n52571));
    SB_LUT4 add_5206_14_lut (.I0(GND_net), .I1(n18896[11]), .I2(n968), 
            .I3(n52937), .O(n17907[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n52569), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_14 (.CI(n52937), .I0(n18896[11]), .I1(n968), .CO(n52938));
    SB_LUT4 add_5206_13_lut (.I0(GND_net), .I1(n18896[10]), .I2(n895), 
            .I3(n52936), .O(n17907[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_13 (.CI(n52936), .I0(n18896[10]), .I1(n895), .CO(n52937));
    SB_LUT4 add_5206_12_lut (.I0(GND_net), .I1(n18896[9]), .I2(n822), 
            .I3(n52935), .O(n17907[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_12 (.CI(n52935), .I0(n18896[9]), .I1(n822), .CO(n52936));
    SB_LUT4 add_5206_11_lut (.I0(GND_net), .I1(n18896[8]), .I2(n749), 
            .I3(n52934), .O(n17907[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_11 (.CI(n52934), .I0(n18896[8]), .I1(n749), .CO(n52935));
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4458));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5206_10_lut (.I0(GND_net), .I1(n18896[7]), .I2(n676), 
            .I3(n52933), .O(n17907[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_10 (.CI(n52933), .I0(n18896[7]), .I1(n676), .CO(n52934));
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4459));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4460));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5206_9_lut (.I0(GND_net), .I1(n18896[6]), .I2(n603), .I3(n52932), 
            .O(n17907[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4461));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4462));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5206_9 (.CI(n52932), .I0(n18896[6]), .I1(n603), .CO(n52933));
    SB_LUT4 add_5206_8_lut (.I0(GND_net), .I1(n18896[5]), .I2(n530), .I3(n52931), 
            .O(n17907[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5206_8 (.CI(n52931), .I0(n18896[5]), .I1(n530), .CO(n52932));
    SB_LUT4 add_5206_7_lut (.I0(GND_net), .I1(n18896[4]), .I2(n457), .I3(n52930), 
            .O(n17907[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_11 (.CI(n52569), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n52570));
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5206_7 (.CI(n52930), .I0(n18896[4]), .I1(n457), .CO(n52931));
    SB_LUT4 add_5206_6_lut (.I0(GND_net), .I1(n18896[3]), .I2(n384), .I3(n52929), 
            .O(n17907[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4464));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n52568), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_6 (.CI(n52929), .I0(n18896[3]), .I1(n384), .CO(n52930));
    SB_LUT4 add_5206_5_lut (.I0(GND_net), .I1(n18896[2]), .I2(n311), .I3(n52928), 
            .O(n17907[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_5 (.CI(n52928), .I0(n18896[2]), .I1(n311), .CO(n52929));
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5206_4_lut (.I0(GND_net), .I1(n18896[1]), .I2(n238), .I3(n52927), 
            .O(n17907[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_4 (.CI(n52927), .I0(n18896[1]), .I1(n238), .CO(n52928));
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_10 (.CI(n52568), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n52569));
    SB_LUT4 add_5206_3_lut (.I0(GND_net), .I1(n18896[0]), .I2(n165), .I3(n52926), 
            .O(n17907[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_3 (.CI(n52926), .I0(n18896[0]), .I1(n165), .CO(n52927));
    SB_LUT4 add_5206_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n17907[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n52926));
    SB_LUT4 add_5483_10_lut (.I0(GND_net), .I1(n22752[7]), .I2(n700), 
            .I3(n52925), .O(n22573[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4465));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_9_lut (.I0(GND_net), .I1(n22752[6]), .I2(n627), .I3(n52924), 
            .O(n22573[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5483_9 (.CI(n52924), .I0(n22752[6]), .I1(n627), .CO(n52925));
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n52567), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4466));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_8_lut (.I0(GND_net), .I1(n22752[5]), .I2(n554_adj_4467), 
            .I3(n52923), .O(n22573[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n52567), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n52568));
    SB_CARRY add_5483_8 (.CI(n52923), .I0(n22752[5]), .I1(n554_adj_4467), 
            .CO(n52924));
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_7_lut (.I0(GND_net), .I1(n22752[4]), .I2(n481), .I3(n52922), 
            .O(n22573[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5483_7 (.CI(n52922), .I0(n22752[4]), .I1(n481), .CO(n52923));
    SB_LUT4 add_5483_6_lut (.I0(GND_net), .I1(n22752[3]), .I2(n408), .I3(n52921), 
            .O(n22573[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5483_6 (.CI(n52921), .I0(n22752[3]), .I1(n408), .CO(n52922));
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4468));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_5_lut (.I0(GND_net), .I1(n22752[2]), .I2(n335_c), 
            .I3(n52920), .O(n22573[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5483_5 (.CI(n52920), .I0(n22752[2]), .I1(n335_c), .CO(n52921));
    SB_LUT4 add_5483_4_lut (.I0(GND_net), .I1(n22752[1]), .I2(n262), .I3(n52919), 
            .O(n22573[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4469));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4470));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5483_4 (.CI(n52919), .I0(n22752[1]), .I1(n262), .CO(n52920));
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_3_lut (.I0(GND_net), .I1(n22752[0]), .I2(n189), .I3(n52918), 
            .O(n22573[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5483_3 (.CI(n52918), .I0(n22752[0]), .I1(n189), .CO(n52919));
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4471));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5483_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n22573[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5483_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5483_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n52918));
    SB_LUT4 add_5254_17_lut (.I0(GND_net), .I1(n19756[14]), .I2(GND_net), 
            .I3(n52917), .O(n18896[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_16_lut (.I0(GND_net), .I1(n19756[13]), .I2(n1117), 
            .I3(n52916), .O(n18896[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_16 (.CI(n52916), .I0(n19756[13]), .I1(n1117), .CO(n52917));
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n52566), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_8 (.CI(n52566), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n52567));
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4472));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4473));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5254_15_lut (.I0(GND_net), .I1(n19756[12]), .I2(n1044_adj_4474), 
            .I3(n52915), .O(n18896[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_15 (.CI(n52915), .I0(n19756[12]), .I1(n1044_adj_4474), 
            .CO(n52916));
    SB_LUT4 add_5254_14_lut (.I0(GND_net), .I1(n19756[11]), .I2(n971_adj_4475), 
            .I3(n52914), .O(n18896[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_14 (.CI(n52914), .I0(n19756[11]), .I1(n971_adj_4475), 
            .CO(n52915));
    SB_LUT4 add_5254_13_lut (.I0(GND_net), .I1(n19756[10]), .I2(n898_adj_4476), 
            .I3(n52913), .O(n18896[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_13 (.CI(n52913), .I0(n19756[10]), .I1(n898_adj_4476), 
            .CO(n52914));
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4477));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5172_19_lut (.I0(GND_net), .I1(n18235[16]), .I2(GND_net), 
            .I3(n53598), .O(n17167[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_12_lut (.I0(GND_net), .I1(n19756[9]), .I2(n825_adj_4478), 
            .I3(n52912), .O(n18896[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_12 (.CI(n52912), .I0(n19756[9]), .I1(n825_adj_4478), 
            .CO(n52913));
    SB_LUT4 add_5172_18_lut (.I0(GND_net), .I1(n18235[15]), .I2(GND_net), 
            .I3(n53597), .O(n17167[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_11_lut (.I0(GND_net), .I1(n19756[8]), .I2(n752_adj_4479), 
            .I3(n52911), .O(n18896[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_18 (.CI(n53597), .I0(n18235[15]), .I1(GND_net), 
            .CO(n53598));
    SB_CARRY add_5254_11 (.CI(n52911), .I0(n19756[8]), .I1(n752_adj_4479), 
            .CO(n52912));
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4480));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5254_10_lut (.I0(GND_net), .I1(n19756[7]), .I2(n679_adj_4481), 
            .I3(n52910), .O(n18896[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4448));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5254_10 (.CI(n52910), .I0(n19756[7]), .I1(n679_adj_4481), 
            .CO(n52911));
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4482));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5254_9_lut (.I0(GND_net), .I1(n19756[6]), .I2(n606_adj_4483), 
            .I3(n52909), .O(n18896[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_9 (.CI(n52909), .I0(n19756[6]), .I1(n606_adj_4483), 
            .CO(n52910));
    SB_LUT4 add_5172_17_lut (.I0(GND_net), .I1(n18235[14]), .I2(GND_net), 
            .I3(n53596), .O(n17167[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_8_lut (.I0(GND_net), .I1(n19756[5]), .I2(n533_adj_4484), 
            .I3(n52908), .O(n18896[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_17 (.CI(n53596), .I0(n18235[14]), .I1(GND_net), 
            .CO(n53597));
    SB_LUT4 add_5172_16_lut (.I0(GND_net), .I1(n18235[13]), .I2(n1111_adj_4485), 
            .I3(n53595), .O(n17167[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_16 (.CI(n53595), .I0(n18235[13]), .I1(n1111_adj_4485), 
            .CO(n53596));
    SB_CARRY add_5254_8 (.CI(n52908), .I0(n19756[5]), .I1(n533_adj_4484), 
            .CO(n52909));
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4486));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5172_15_lut (.I0(GND_net), .I1(n18235[12]), .I2(n1038_adj_4487), 
            .I3(n53594), .O(n17167[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_15 (.CI(n53594), .I0(n18235[12]), .I1(n1038_adj_4487), 
            .CO(n53595));
    SB_LUT4 add_5172_14_lut (.I0(GND_net), .I1(n18235[11]), .I2(n965_adj_4488), 
            .I3(n53593), .O(n17167[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_14 (.CI(n53593), .I0(n18235[11]), .I1(n965_adj_4488), 
            .CO(n53594));
    SB_LUT4 add_5172_13_lut (.I0(GND_net), .I1(n18235[10]), .I2(n892_adj_4489), 
            .I3(n53592), .O(n17167[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_13 (.CI(n53592), .I0(n18235[10]), .I1(n892_adj_4489), 
            .CO(n53593));
    SB_LUT4 add_5172_12_lut (.I0(GND_net), .I1(n18235[9]), .I2(n819_adj_4490), 
            .I3(n53591), .O(n17167[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_12 (.CI(n53591), .I0(n18235[9]), .I1(n819_adj_4490), 
            .CO(n53592));
    SB_LUT4 add_5172_11_lut (.I0(GND_net), .I1(n18235[8]), .I2(n746_adj_4491), 
            .I3(n53590), .O(n17167[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_11 (.CI(n53590), .I0(n18235[8]), .I1(n746_adj_4491), 
            .CO(n53591));
    SB_LUT4 add_5172_10_lut (.I0(GND_net), .I1(n18235[7]), .I2(n673_adj_4492), 
            .I3(n53589), .O(n17167[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_10 (.CI(n53589), .I0(n18235[7]), .I1(n673_adj_4492), 
            .CO(n53590));
    SB_LUT4 add_5172_9_lut (.I0(GND_net), .I1(n18235[6]), .I2(n600_adj_4493), 
            .I3(n53588), .O(n17167[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_9 (.CI(n53588), .I0(n18235[6]), .I1(n600_adj_4493), 
            .CO(n53589));
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4494));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4495));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4496));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5172_8_lut (.I0(GND_net), .I1(n18235[5]), .I2(n527_adj_4498), 
            .I3(n53587), .O(n17167[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_8 (.CI(n53587), .I0(n18235[5]), .I1(n527_adj_4498), 
            .CO(n53588));
    SB_LUT4 add_5172_7_lut (.I0(GND_net), .I1(n18235[4]), .I2(n454_adj_4499), 
            .I3(n53586), .O(n17167[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_7 (.CI(n53586), .I0(n18235[4]), .I1(n454_adj_4499), 
            .CO(n53587));
    SB_LUT4 add_5254_7_lut (.I0(GND_net), .I1(n19756[4]), .I2(n460_adj_4500), 
            .I3(n52907), .O(n18896[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_7 (.CI(n52907), .I0(n19756[4]), .I1(n460_adj_4500), 
            .CO(n52908));
    SB_LUT4 add_5172_6_lut (.I0(GND_net), .I1(n18235[3]), .I2(n381_adj_4501), 
            .I3(n53585), .O(n17167[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_6 (.CI(n53585), .I0(n18235[3]), .I1(n381_adj_4501), 
            .CO(n53586));
    SB_LUT4 add_5172_5_lut (.I0(GND_net), .I1(n18235[2]), .I2(n308_adj_4502), 
            .I3(n53584), .O(n17167[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_6_lut (.I0(GND_net), .I1(n19756[3]), .I2(n387_adj_4503), 
            .I3(n52906), .O(n18896[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_5 (.CI(n53584), .I0(n18235[2]), .I1(n308_adj_4502), 
            .CO(n53585));
    SB_LUT4 add_5172_4_lut (.I0(GND_net), .I1(n18235[1]), .I2(n235_adj_4504), 
            .I3(n53583), .O(n17167[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_4 (.CI(n53583), .I0(n18235[1]), .I1(n235_adj_4504), 
            .CO(n53584));
    SB_CARRY add_5254_6 (.CI(n52906), .I0(n19756[3]), .I1(n387_adj_4503), 
            .CO(n52907));
    SB_LUT4 add_5172_3_lut (.I0(GND_net), .I1(n18235[0]), .I2(n162_adj_4505), 
            .I3(n53582), .O(n17167[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_3 (.CI(n53582), .I0(n18235[0]), .I1(n162_adj_4505), 
            .CO(n53583));
    SB_LUT4 add_5172_2_lut (.I0(GND_net), .I1(n20_adj_4506), .I2(n89_adj_4507), 
            .I3(GND_net), .O(n17167[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_5_lut (.I0(GND_net), .I1(n19756[2]), .I2(n314_adj_4508), 
            .I3(n52905), .O(n18896[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_5 (.CI(n52905), .I0(n19756[2]), .I1(n314_adj_4508), 
            .CO(n52906));
    SB_CARRY add_5172_2 (.CI(GND_net), .I0(n20_adj_4506), .I1(n89_adj_4507), 
            .CO(n53582));
    SB_LUT4 add_5223_18_lut (.I0(GND_net), .I1(n19169[15]), .I2(GND_net), 
            .I3(n53581), .O(n18235[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_4_lut (.I0(GND_net), .I1(n19756[1]), .I2(n241_adj_4509), 
            .I3(n52904), .O(n18896[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5223_17_lut (.I0(GND_net), .I1(n19169[14]), .I2(GND_net), 
            .I3(n53580), .O(n18235[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_17 (.CI(n53580), .I0(n19169[14]), .I1(GND_net), 
            .CO(n53581));
    SB_LUT4 add_5223_16_lut (.I0(GND_net), .I1(n19169[13]), .I2(n1114_adj_4510), 
            .I3(n53579), .O(n18235[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n52565), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_4 (.CI(n52904), .I0(n19756[1]), .I1(n241_adj_4509), 
            .CO(n52905));
    SB_CARRY add_5223_16 (.CI(n53579), .I0(n19169[13]), .I1(n1114_adj_4510), 
            .CO(n53580));
    SB_LUT4 add_5223_15_lut (.I0(GND_net), .I1(n19169[12]), .I2(n1041_adj_4511), 
            .I3(n53578), .O(n18235[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_7 (.CI(n52565), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n52566));
    SB_CARRY add_5223_15 (.CI(n53578), .I0(n19169[12]), .I1(n1041_adj_4511), 
            .CO(n53579));
    SB_LUT4 add_5223_14_lut (.I0(GND_net), .I1(n19169[11]), .I2(n968_adj_4512), 
            .I3(n53577), .O(n18235[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_14 (.CI(n53577), .I0(n19169[11]), .I1(n968_adj_4512), 
            .CO(n53578));
    SB_LUT4 add_5223_13_lut (.I0(GND_net), .I1(n19169[10]), .I2(n895_adj_4513), 
            .I3(n53576), .O(n18235[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_13 (.CI(n53576), .I0(n19169[10]), .I1(n895_adj_4513), 
            .CO(n53577));
    SB_LUT4 add_5223_12_lut (.I0(GND_net), .I1(n19169[9]), .I2(n822_adj_4514), 
            .I3(n53575), .O(n18235[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_12 (.CI(n53575), .I0(n19169[9]), .I1(n822_adj_4514), 
            .CO(n53576));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(n8), 
            .I3(n52570), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_3_lut (.I0(GND_net), .I1(n19756[0]), .I2(n168_adj_4515), 
            .I3(n52903), .O(n18896[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4516));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4517));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5254_3 (.CI(n52903), .I0(n19756[0]), .I1(n168_adj_4515), 
            .CO(n52904));
    SB_LUT4 add_5254_2_lut (.I0(GND_net), .I1(n26_adj_4518), .I2(n95_adj_4519), 
            .I3(GND_net), .O(n18896[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5223_11_lut (.I0(GND_net), .I1(n19169[8]), .I2(n749_adj_4520), 
            .I3(n53574), .O(n18235[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_2 (.CI(GND_net), .I0(n26_adj_4518), .I1(n95_adj_4519), 
            .CO(n52903));
    SB_CARRY add_5223_11 (.CI(n53574), .I0(n19169[8]), .I1(n749_adj_4520), 
            .CO(n53575));
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n52564), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5223_10_lut (.I0(GND_net), .I1(n19169[7]), .I2(n676_adj_4521), 
            .I3(n53573), .O(n18235[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_10 (.CI(n53573), .I0(n19169[7]), .I1(n676_adj_4521), 
            .CO(n53574));
    SB_CARRY sub_15_add_2_6 (.CI(n52564), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n52565));
    SB_LUT4 add_5223_9_lut (.I0(GND_net), .I1(n19169[6]), .I2(n603_adj_4522), 
            .I3(n53572), .O(n18235[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_9 (.CI(n53572), .I0(n19169[6]), .I1(n603_adj_4522), 
            .CO(n53573));
    SB_LUT4 add_5223_8_lut (.I0(GND_net), .I1(n19169[5]), .I2(n530_adj_4523), 
            .I3(n53571), .O(n18235[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_8 (.CI(n53571), .I0(n19169[5]), .I1(n530_adj_4523), 
            .CO(n53572));
    SB_CARRY sub_15_add_2_5 (.CI(n52563), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n52564));
    SB_LUT4 add_5299_16_lut (.I0(GND_net), .I1(n20475[13]), .I2(n1120_adj_4517), 
            .I3(n52902), .O(n19756[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_15_lut (.I0(GND_net), .I1(n20475[12]), .I2(n1047_adj_4516), 
            .I3(n52901), .O(n19756[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_15 (.CI(n52901), .I0(n20475[12]), .I1(n1047_adj_4516), 
            .CO(n52902));
    SB_LUT4 add_5299_14_lut (.I0(GND_net), .I1(n20475[11]), .I2(n974_adj_4497), 
            .I3(n52900), .O(n19756[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5223_7_lut (.I0(GND_net), .I1(n19169[4]), .I2(n457_adj_4496), 
            .I3(n53570), .O(n18235[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_7 (.CI(n53570), .I0(n19169[4]), .I1(n457_adj_4496), 
            .CO(n53571));
    SB_LUT4 add_5223_6_lut (.I0(GND_net), .I1(n19169[3]), .I2(n384_adj_4495), 
            .I3(n53569), .O(n18235[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_6 (.CI(n53569), .I0(n19169[3]), .I1(n384_adj_4495), 
            .CO(n53570));
    SB_LUT4 add_5223_5_lut (.I0(GND_net), .I1(n19169[2]), .I2(n311_adj_4494), 
            .I3(n53568), .O(n18235[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_5 (.CI(n53568), .I0(n19169[2]), .I1(n311_adj_4494), 
            .CO(n53569));
    SB_CARRY add_5299_14 (.CI(n52900), .I0(n20475[11]), .I1(n974_adj_4497), 
            .CO(n52901));
    SB_LUT4 add_5223_4_lut (.I0(GND_net), .I1(n19169[1]), .I2(n238_adj_4486), 
            .I3(n53567), .O(n18235[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_4 (.CI(n53567), .I0(n19169[1]), .I1(n238_adj_4486), 
            .CO(n53568));
    SB_LUT4 add_5299_13_lut (.I0(GND_net), .I1(n20475[10]), .I2(n901_adj_4482), 
            .I3(n52899), .O(n19756[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5223_3_lut (.I0(GND_net), .I1(n19169[0]), .I2(n165_adj_4480), 
            .I3(n53566), .O(n18235[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_3 (.CI(n53566), .I0(n19169[0]), .I1(n165_adj_4480), 
            .CO(n53567));
    SB_CARRY add_5299_13 (.CI(n52899), .I0(n20475[10]), .I1(n901_adj_4482), 
            .CO(n52900));
    SB_LUT4 add_5223_2_lut (.I0(GND_net), .I1(n23_adj_4477), .I2(n92_adj_4473), 
            .I3(GND_net), .O(n18235[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5223_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5223_2 (.CI(GND_net), .I0(n23_adj_4477), .I1(n92_adj_4473), 
            .CO(n53566));
    SB_LUT4 add_5269_17_lut (.I0(GND_net), .I1(n19977[14]), .I2(GND_net), 
            .I3(n53565), .O(n19169[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5269_16_lut (.I0(GND_net), .I1(n19977[13]), .I2(n1117_adj_4472), 
            .I3(n53564), .O(n19169[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_12_lut (.I0(GND_net), .I1(n20475[9]), .I2(n828_adj_4471), 
            .I3(n52898), .O(n19756[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_16 (.CI(n53564), .I0(n19977[13]), .I1(n1117_adj_4472), 
            .CO(n53565));
    SB_LUT4 add_5269_15_lut (.I0(GND_net), .I1(n19977[12]), .I2(n1044), 
            .I3(n53563), .O(n19169[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_12 (.CI(n52898), .I0(n20475[9]), .I1(n828_adj_4471), 
            .CO(n52899));
    SB_CARRY add_5269_15 (.CI(n53563), .I0(n19977[12]), .I1(n1044), .CO(n53564));
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4523));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5269_14_lut (.I0(GND_net), .I1(n19977[11]), .I2(n971), 
            .I3(n53562), .O(n19169[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_14 (.CI(n53562), .I0(n19977[11]), .I1(n971), .CO(n53563));
    SB_LUT4 add_5269_13_lut (.I0(GND_net), .I1(n19977[10]), .I2(n898), 
            .I3(n53561), .O(n19169[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_13 (.CI(n53561), .I0(n19977[10]), .I1(n898), .CO(n53562));
    SB_LUT4 add_5269_12_lut (.I0(GND_net), .I1(n19977[9]), .I2(n825), 
            .I3(n53560), .O(n19169[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_11_lut (.I0(GND_net), .I1(n20475[8]), .I2(n755_adj_4470), 
            .I3(n52897), .O(n19756[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_11 (.CI(n52897), .I0(n20475[8]), .I1(n755_adj_4470), 
            .CO(n52898));
    SB_LUT4 add_5299_10_lut (.I0(GND_net), .I1(n20475[7]), .I2(n682_adj_4469), 
            .I3(n52896), .O(n19756[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_10 (.CI(n52896), .I0(n20475[7]), .I1(n682_adj_4469), 
            .CO(n52897));
    SB_LUT4 add_5299_9_lut (.I0(GND_net), .I1(n20475[6]), .I2(n609_adj_4468), 
            .I3(n52895), .O(n19756[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_12 (.CI(n53560), .I0(n19977[9]), .I1(n825), .CO(n53561));
    SB_CARRY add_5299_9 (.CI(n52895), .I0(n20475[6]), .I1(n609_adj_4468), 
            .CO(n52896));
    SB_LUT4 add_5269_11_lut (.I0(GND_net), .I1(n19977[8]), .I2(n752), 
            .I3(n53559), .O(n19169[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_11 (.CI(n53559), .I0(n19977[8]), .I1(n752), .CO(n53560));
    SB_LUT4 add_5269_10_lut (.I0(GND_net), .I1(n19977[7]), .I2(n679), 
            .I3(n53558), .O(n19169[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4522));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5269_10 (.CI(n53558), .I0(n19977[7]), .I1(n679), .CO(n53559));
    SB_LUT4 add_5269_9_lut (.I0(GND_net), .I1(n19977[6]), .I2(n606), .I3(n53557), 
            .O(n19169[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_9 (.CI(n53557), .I0(n19977[6]), .I1(n606), .CO(n53558));
    SB_LUT4 add_5269_8_lut (.I0(GND_net), .I1(n19977[5]), .I2(n533), .I3(n53556), 
            .O(n19169[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4521));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5269_8 (.CI(n53556), .I0(n19977[5]), .I1(n533), .CO(n53557));
    SB_LUT4 add_5269_7_lut (.I0(GND_net), .I1(n19977[4]), .I2(n460), .I3(n53555), 
            .O(n19169[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_8_lut (.I0(GND_net), .I1(n20475[5]), .I2(n536_adj_4466), 
            .I3(n52894), .O(n19756[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_7 (.CI(n53555), .I0(n19977[4]), .I1(n460), .CO(n53556));
    SB_LUT4 add_5269_6_lut (.I0(GND_net), .I1(n19977[3]), .I2(n387), .I3(n53554), 
            .O(n19169[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_6 (.CI(n53554), .I0(n19977[3]), .I1(n387), .CO(n53555));
    SB_LUT4 add_5269_5_lut (.I0(GND_net), .I1(n19977[2]), .I2(n314), .I3(n53553), 
            .O(n19169[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_8 (.CI(n52894), .I0(n20475[5]), .I1(n536_adj_4466), 
            .CO(n52895));
    SB_CARRY add_5269_5 (.CI(n53553), .I0(n19977[2]), .I1(n314), .CO(n53554));
    SB_LUT4 add_5269_4_lut (.I0(GND_net), .I1(n19977[1]), .I2(n241), .I3(n53552), 
            .O(n19169[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_4 (.CI(n53552), .I0(n19977[1]), .I1(n241), .CO(n53553));
    SB_LUT4 add_5269_3_lut (.I0(GND_net), .I1(n19977[0]), .I2(n168), .I3(n53551), 
            .O(n19169[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_7_lut (.I0(GND_net), .I1(n20475[4]), .I2(n463_adj_4465), 
            .I3(n52893), .O(n19756[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_3 (.CI(n53551), .I0(n19977[0]), .I1(n168), .CO(n53552));
    SB_LUT4 add_5269_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n19169[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n53551));
    SB_CARRY add_5299_7 (.CI(n52893), .I0(n20475[4]), .I1(n463_adj_4465), 
            .CO(n52894));
    SB_LUT4 add_5312_16_lut (.I0(GND_net), .I1(n20667[13]), .I2(n1120), 
            .I3(n53550), .O(n19977[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5312_15_lut (.I0(GND_net), .I1(n20667[12]), .I2(n1047), 
            .I3(n53549), .O(n19977[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_6_lut (.I0(GND_net), .I1(n20475[3]), .I2(n390_adj_4464), 
            .I3(n52892), .O(n19756[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_15 (.CI(n53549), .I0(n20667[12]), .I1(n1047), .CO(n53550));
    SB_LUT4 add_5312_14_lut (.I0(GND_net), .I1(n20667[11]), .I2(n974), 
            .I3(n53548), .O(n19977[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_14 (.CI(n53548), .I0(n20667[11]), .I1(n974), .CO(n53549));
    SB_LUT4 add_5312_13_lut (.I0(GND_net), .I1(n20667[10]), .I2(n901), 
            .I3(n53547), .O(n19977[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_13 (.CI(n53547), .I0(n20667[10]), .I1(n901), .CO(n53548));
    SB_LUT4 add_5312_12_lut (.I0(GND_net), .I1(n20667[9]), .I2(n828), 
            .I3(n53546), .O(n19977[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_12 (.CI(n53546), .I0(n20667[9]), .I1(n828), .CO(n53547));
    SB_LUT4 add_5312_11_lut (.I0(GND_net), .I1(n20667[8]), .I2(n755), 
            .I3(n53545), .O(n19977[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_11 (.CI(n53545), .I0(n20667[8]), .I1(n755), .CO(n53546));
    SB_LUT4 add_5312_10_lut (.I0(GND_net), .I1(n20667[7]), .I2(n682), 
            .I3(n53544), .O(n19977[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_10 (.CI(n53544), .I0(n20667[7]), .I1(n682), .CO(n53545));
    SB_LUT4 add_5312_9_lut (.I0(GND_net), .I1(n20667[6]), .I2(n609), .I3(n53543), 
            .O(n19977[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_9 (.CI(n53543), .I0(n20667[6]), .I1(n609), .CO(n53544));
    SB_LUT4 add_5312_8_lut (.I0(GND_net), .I1(n20667[5]), .I2(n536_adj_4463), 
            .I3(n53542), .O(n19977[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_8 (.CI(n53542), .I0(n20667[5]), .I1(n536_adj_4463), 
            .CO(n53543));
    SB_LUT4 add_5312_7_lut (.I0(GND_net), .I1(n20667[4]), .I2(n463), .I3(n53541), 
            .O(n19977[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_7 (.CI(n53541), .I0(n20667[4]), .I1(n463), .CO(n53542));
    SB_LUT4 add_5312_6_lut (.I0(GND_net), .I1(n20667[3]), .I2(n390), .I3(n53540), 
            .O(n19977[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_6 (.CI(n53540), .I0(n20667[3]), .I1(n390), .CO(n53541));
    SB_LUT4 add_5312_5_lut (.I0(GND_net), .I1(n20667[2]), .I2(n317_adj_4462), 
            .I3(n53539), .O(n19977[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_5 (.CI(n53539), .I0(n20667[2]), .I1(n317_adj_4462), 
            .CO(n53540));
    SB_LUT4 add_5312_4_lut (.I0(GND_net), .I1(n20667[1]), .I2(n244_adj_4461), 
            .I3(n53538), .O(n19977[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_4 (.CI(n53538), .I0(n20667[1]), .I1(n244_adj_4461), 
            .CO(n53539));
    SB_LUT4 add_5312_3_lut (.I0(GND_net), .I1(n20667[0]), .I2(n171_adj_4460), 
            .I3(n53537), .O(n19977[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5312_3 (.CI(n53537), .I0(n20667[0]), .I1(n171_adj_4460), 
            .CO(n53538));
    SB_LUT4 add_5312_2_lut (.I0(GND_net), .I1(n29_adj_4459), .I2(n98_adj_4458), 
            .I3(GND_net), .O(n19977[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5312_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_6 (.CI(n52892), .I0(n20475[3]), .I1(n390_adj_4464), 
            .CO(n52893));
    SB_CARRY add_5312_2 (.CI(GND_net), .I0(n29_adj_4459), .I1(n98_adj_4458), 
            .CO(n53537));
    SB_LUT4 add_5350_15_lut (.I0(GND_net), .I1(n21245[12]), .I2(n1050), 
            .I3(n53536), .O(n20667[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5350_14_lut (.I0(GND_net), .I1(n21245[11]), .I2(n977), 
            .I3(n53535), .O(n20667[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_14 (.CI(n53535), .I0(n21245[11]), .I1(n977), .CO(n53536));
    SB_LUT4 add_5299_5_lut (.I0(GND_net), .I1(n20475[2]), .I2(n317), .I3(n52891), 
            .O(n19756[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5350_13_lut (.I0(GND_net), .I1(n21245[10]), .I2(n904), 
            .I3(n53534), .O(n20667[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_13 (.CI(n53534), .I0(n21245[10]), .I1(n904), .CO(n53535));
    SB_LUT4 add_5350_12_lut (.I0(GND_net), .I1(n21245[9]), .I2(n831), 
            .I3(n53533), .O(n20667[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_12 (.CI(n53533), .I0(n21245[9]), .I1(n831), .CO(n53534));
    SB_LUT4 add_5350_11_lut (.I0(GND_net), .I1(n21245[8]), .I2(n758), 
            .I3(n53532), .O(n20667[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_11 (.CI(n53532), .I0(n21245[8]), .I1(n758), .CO(n53533));
    SB_LUT4 add_5350_10_lut (.I0(GND_net), .I1(n21245[7]), .I2(n685), 
            .I3(n53531), .O(n20667[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_10 (.CI(n53531), .I0(n21245[7]), .I1(n685), .CO(n53532));
    SB_LUT4 add_5350_9_lut (.I0(GND_net), .I1(n21245[6]), .I2(n612), .I3(n53530), 
            .O(n20667[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_9 (.CI(n53530), .I0(n21245[6]), .I1(n612), .CO(n53531));
    SB_CARRY add_5299_5 (.CI(n52891), .I0(n20475[2]), .I1(n317), .CO(n52892));
    SB_LUT4 add_5350_8_lut (.I0(GND_net), .I1(n21245[5]), .I2(n539), .I3(n53529), 
            .O(n20667[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_4_lut (.I0(GND_net), .I1(n20475[1]), .I2(n244), .I3(n52890), 
            .O(n19756[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_4 (.CI(n52890), .I0(n20475[1]), .I1(n244), .CO(n52891));
    SB_LUT4 add_5299_3_lut (.I0(GND_net), .I1(n20475[0]), .I2(n171), .I3(n52889), 
            .O(n19756[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_8 (.CI(n53529), .I0(n21245[5]), .I1(n539), .CO(n53530));
    SB_LUT4 add_5350_7_lut (.I0(GND_net), .I1(n21245[4]), .I2(n466), .I3(n53528), 
            .O(n20667[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_7 (.CI(n53528), .I0(n21245[4]), .I1(n466), .CO(n53529));
    SB_LUT4 add_5350_6_lut (.I0(GND_net), .I1(n21245[3]), .I2(n393), .I3(n53527), 
            .O(n20667[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_6 (.CI(n53527), .I0(n21245[3]), .I1(n393), .CO(n53528));
    SB_CARRY add_5299_3 (.CI(n52889), .I0(n20475[0]), .I1(n171), .CO(n52890));
    SB_LUT4 add_5350_5_lut (.I0(GND_net), .I1(n21245[2]), .I2(n320), .I3(n53526), 
            .O(n20667[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_5 (.CI(n53526), .I0(n21245[2]), .I1(n320), .CO(n53527));
    SB_LUT4 add_5350_4_lut (.I0(GND_net), .I1(n21245[1]), .I2(n247), .I3(n53525), 
            .O(n20667[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_4 (.CI(n53525), .I0(n21245[1]), .I1(n247), .CO(n53526));
    SB_LUT4 add_5350_3_lut (.I0(GND_net), .I1(n21245[0]), .I2(n174), .I3(n53524), 
            .O(n20667[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n19756[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_3 (.CI(n53524), .I0(n21245[0]), .I1(n174), .CO(n53525));
    SB_CARRY add_5299_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n52889));
    SB_LUT4 add_5338_15_lut (.I0(GND_net), .I1(n21080[12]), .I2(n1050_adj_4524), 
            .I3(n52888), .O(n20475[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5350_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n20667[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5350_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5350_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n53524));
    SB_LUT4 add_5338_14_lut (.I0(GND_net), .I1(n21080[11]), .I2(n977_adj_4525), 
            .I3(n52887), .O(n20475[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_14_lut (.I0(GND_net), .I1(n21718[11]), .I2(n980), 
            .I3(n53523), .O(n21245[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_13_lut (.I0(GND_net), .I1(n21718[10]), .I2(n907), 
            .I3(n53522), .O(n21245[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_13 (.CI(n53522), .I0(n21718[10]), .I1(n907), .CO(n53523));
    SB_LUT4 add_5385_12_lut (.I0(GND_net), .I1(n21718[9]), .I2(n834), 
            .I3(n53521), .O(n21245[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_12 (.CI(n53521), .I0(n21718[9]), .I1(n834), .CO(n53522));
    SB_LUT4 add_5385_11_lut (.I0(GND_net), .I1(n21718[8]), .I2(n761), 
            .I3(n53520), .O(n21245[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_14 (.CI(n52887), .I0(n21080[11]), .I1(n977_adj_4525), 
            .CO(n52888));
    SB_CARRY add_5385_11 (.CI(n53520), .I0(n21718[8]), .I1(n761), .CO(n53521));
    SB_LUT4 add_5385_10_lut (.I0(GND_net), .I1(n21718[7]), .I2(n688), 
            .I3(n53519), .O(n21245[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_10 (.CI(n53519), .I0(n21718[7]), .I1(n688), .CO(n53520));
    SB_LUT4 add_5385_9_lut (.I0(GND_net), .I1(n21718[6]), .I2(n615), .I3(n53518), 
            .O(n21245[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_13_lut (.I0(GND_net), .I1(n21080[10]), .I2(n904_adj_4526), 
            .I3(n52886), .O(n20475[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_9 (.CI(n53518), .I0(n21718[6]), .I1(n615), .CO(n53519));
    SB_LUT4 add_5385_8_lut (.I0(GND_net), .I1(n21718[5]), .I2(n542), .I3(n53517), 
            .O(n21245[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_8 (.CI(n53517), .I0(n21718[5]), .I1(n542), .CO(n53518));
    SB_CARRY add_5338_13 (.CI(n52886), .I0(n21080[10]), .I1(n904_adj_4526), 
            .CO(n52887));
    SB_LUT4 add_5385_7_lut (.I0(GND_net), .I1(n21718[4]), .I2(n469), .I3(n53516), 
            .O(n21245[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_7 (.CI(n53516), .I0(n21718[4]), .I1(n469), .CO(n53517));
    SB_LUT4 add_5385_6_lut (.I0(GND_net), .I1(n21718[3]), .I2(n396), .I3(n53515), 
            .O(n21245[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_6 (.CI(n53515), .I0(n21718[3]), .I1(n396), .CO(n53516));
    SB_LUT4 add_5338_12_lut (.I0(GND_net), .I1(n21080[9]), .I2(n831_adj_4527), 
            .I3(n52885), .O(n20475[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_5_lut (.I0(GND_net), .I1(n21718[2]), .I2(n323), .I3(n53514), 
            .O(n21245[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_12 (.CI(n52885), .I0(n21080[9]), .I1(n831_adj_4527), 
            .CO(n52886));
    SB_LUT4 add_5338_11_lut (.I0(GND_net), .I1(n21080[8]), .I2(n758_adj_4528), 
            .I3(n52884), .O(n20475[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_5 (.CI(n53514), .I0(n21718[2]), .I1(n323), .CO(n53515));
    SB_CARRY add_5338_11 (.CI(n52884), .I0(n21080[8]), .I1(n758_adj_4528), 
            .CO(n52885));
    SB_LUT4 add_5385_4_lut (.I0(GND_net), .I1(n21718[1]), .I2(n250), .I3(n53513), 
            .O(n21245[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_4 (.CI(n53513), .I0(n21718[1]), .I1(n250), .CO(n53514));
    SB_LUT4 add_5385_3_lut (.I0(GND_net), .I1(n21718[0]), .I2(n177), .I3(n53512), 
            .O(n21245[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_10_lut (.I0(GND_net), .I1(n21080[7]), .I2(n685_adj_4529), 
            .I3(n52883), .O(n20475[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_3 (.CI(n53512), .I0(n21718[0]), .I1(n177), .CO(n53513));
    SB_LUT4 add_5385_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n21245[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n53512));
    SB_CARRY add_5338_10 (.CI(n52883), .I0(n21080[7]), .I1(n685_adj_4529), 
            .CO(n52884));
    SB_LUT4 add_5338_9_lut (.I0(GND_net), .I1(n21080[6]), .I2(n612_adj_4530), 
            .I3(n52882), .O(n20475[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_9 (.CI(n52882), .I0(n21080[6]), .I1(n612_adj_4530), 
            .CO(n52883));
    SB_LUT4 add_5338_8_lut (.I0(GND_net), .I1(n21080[5]), .I2(n539_adj_4531), 
            .I3(n52881), .O(n20475[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_8 (.CI(n52881), .I0(n21080[5]), .I1(n539_adj_4531), 
            .CO(n52882));
    SB_LUT4 add_5338_7_lut (.I0(GND_net), .I1(n21080[4]), .I2(n466_adj_4532), 
            .I3(n52880), .O(n20475[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_7 (.CI(n52880), .I0(n21080[4]), .I1(n466_adj_4532), 
            .CO(n52881));
    SB_LUT4 add_5338_6_lut (.I0(GND_net), .I1(n21080[3]), .I2(n393_adj_4533), 
            .I3(n52879), .O(n20475[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_6 (.CI(n52879), .I0(n21080[3]), .I1(n393_adj_4533), 
            .CO(n52880));
    SB_LUT4 add_5338_5_lut (.I0(GND_net), .I1(n21080[2]), .I2(n320_adj_4534), 
            .I3(n52878), .O(n20475[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_4 (.CI(n52562), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n52563));
    SB_CARRY add_5338_5 (.CI(n52878), .I0(n21080[2]), .I1(n320_adj_4534), 
            .CO(n52879));
    SB_LUT4 add_5338_4_lut (.I0(GND_net), .I1(n21080[1]), .I2(n247_adj_4535), 
            .I3(n52877), .O(n20475[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_4 (.CI(n52877), .I0(n21080[1]), .I1(n247_adj_4535), 
            .CO(n52878));
    SB_LUT4 add_5338_3_lut (.I0(GND_net), .I1(n21080[0]), .I2(n174_adj_4536), 
            .I3(n52876), .O(n20475[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_3 (.CI(n52561), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n52562));
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n52561));
    SB_CARRY add_5338_3 (.CI(n52876), .I0(n21080[0]), .I1(n174_adj_4536), 
            .CO(n52877));
    SB_LUT4 add_5338_2_lut (.I0(GND_net), .I1(n32_adj_4537), .I2(n101_adj_4538), 
            .I3(GND_net), .O(n20475[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_2 (.CI(GND_net), .I0(n32_adj_4537), .I1(n101_adj_4538), 
            .CO(n52876));
    SB_LUT4 add_5499_9_lut (.I0(GND_net), .I1(n22878[6]), .I2(n630), .I3(n52875), 
            .O(n22752[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5499_8_lut (.I0(GND_net), .I1(n22878[5]), .I2(n557_adj_4539), 
            .I3(n52874), .O(n22752[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_8 (.CI(n52874), .I0(n22878[5]), .I1(n557_adj_4539), 
            .CO(n52875));
    SB_LUT4 add_5499_7_lut (.I0(GND_net), .I1(n22878[4]), .I2(n484), .I3(n52873), 
            .O(n22752[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_7 (.CI(n52873), .I0(n22878[4]), .I1(n484), .CO(n52874));
    SB_LUT4 add_5499_6_lut (.I0(GND_net), .I1(n22878[3]), .I2(n411), .I3(n52872), 
            .O(n22752[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_6 (.CI(n52872), .I0(n22878[3]), .I1(n411), .CO(n52873));
    SB_LUT4 add_5499_5_lut (.I0(GND_net), .I1(n22878[2]), .I2(n338), .I3(n52871), 
            .O(n22752[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5442_12_lut (.I0(GND_net), .I1(n22374[9]), .I2(n840), 
            .I3(n53116), .O(n22091[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5442_11_lut (.I0(GND_net), .I1(n22374[8]), .I2(n767), 
            .I3(n53115), .O(n22091[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_5 (.CI(n52871), .I0(n22878[2]), .I1(n338), .CO(n52872));
    SB_CARRY add_5442_11 (.CI(n53115), .I0(n22374[8]), .I1(n767), .CO(n53116));
    SB_LUT4 add_5442_10_lut (.I0(GND_net), .I1(n22374[7]), .I2(n694), 
            .I3(n53114), .O(n22091[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5499_4_lut (.I0(GND_net), .I1(n22878[1]), .I2(n265), .I3(n52870), 
            .O(n22752[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4520));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5442_10 (.CI(n53114), .I0(n22374[7]), .I1(n694), .CO(n53115));
    SB_LUT4 add_5442_9_lut (.I0(GND_net), .I1(n22374[6]), .I2(n621), .I3(n53113), 
            .O(n22091[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_4 (.CI(n52870), .I0(n22878[1]), .I1(n265), .CO(n52871));
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n335[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR counter_2046_2047__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n71491), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_5442_9 (.CI(n53113), .I0(n22374[6]), .I1(n621), .CO(n53114));
    SB_LUT4 add_5442_8_lut (.I0(GND_net), .I1(n22374[5]), .I2(n548), .I3(n53112), 
            .O(n22091[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5442_8 (.CI(n53112), .I0(n22374[5]), .I1(n548), .CO(n53113));
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4519));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5499_3_lut (.I0(GND_net), .I1(n22878[0]), .I2(n192), .I3(n52869), 
            .O(n22752[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_3 (.CI(n52869), .I0(n22878[0]), .I1(n192), .CO(n52870));
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5442_7_lut (.I0(GND_net), .I1(n22374[4]), .I2(n475_adj_4540), 
            .I3(n53111), .O(n22091[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5442_7 (.CI(n53111), .I0(n22374[4]), .I1(n475_adj_4540), 
            .CO(n53112));
    SB_LUT4 add_5442_6_lut (.I0(GND_net), .I1(n22374[3]), .I2(n402), .I3(n53110), 
            .O(n22091[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5442_6 (.CI(n53110), .I0(n22374[3]), .I1(n402), .CO(n53111));
    SB_LUT4 add_5499_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n22752[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5499_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5442_5_lut (.I0(GND_net), .I1(n22374[2]), .I2(n329), .I3(n53109), 
            .O(n22091[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5499_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n52869));
    SB_CARRY add_5442_5 (.CI(n53109), .I0(n22374[2]), .I1(n329), .CO(n53110));
    SB_LUT4 add_5442_4_lut (.I0(GND_net), .I1(n22374[1]), .I2(n256), .I3(n53108), 
            .O(n22091[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_14_lut (.I0(GND_net), .I1(n21578[11]), .I2(n980_adj_4541), 
            .I3(n52868), .O(n21080[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5442_4 (.CI(n53108), .I0(n22374[1]), .I1(n256), .CO(n53109));
    SB_LUT4 add_5374_13_lut (.I0(GND_net), .I1(n21578[10]), .I2(n907_adj_4542), 
            .I3(n52867), .O(n21080[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5442_3_lut (.I0(GND_net), .I1(n22374[0]), .I2(n183), .I3(n53107), 
            .O(n22091[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_13 (.CI(n52867), .I0(n21578[10]), .I1(n907_adj_4542), 
            .CO(n52868));
    SB_CARRY add_5442_3 (.CI(n53107), .I0(n22374[0]), .I1(n183), .CO(n53108));
    SB_LUT4 add_5442_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n22091[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5442_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_12_lut (.I0(GND_net), .I1(n21578[9]), .I2(n834_adj_4543), 
            .I3(n52866), .O(n21080[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_12 (.CI(n52866), .I0(n21578[9]), .I1(n834_adj_4543), 
            .CO(n52867));
    SB_LUT4 add_5374_11_lut (.I0(GND_net), .I1(n21578[8]), .I2(n761_adj_4544), 
            .I3(n52865), .O(n21080[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5442_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n53107));
    SB_CARRY add_5374_11 (.CI(n52865), .I0(n21578[8]), .I1(n761_adj_4544), 
            .CO(n52866));
    SB_LUT4 add_5374_10_lut (.I0(GND_net), .I1(n21578[7]), .I2(n688_adj_4545), 
            .I3(n52864), .O(n21080[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5525_7_lut (.I0(GND_net), .I1(n61693), .I2(n490), .I3(n53906), 
            .O(n22974[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5525_6_lut (.I0(GND_net), .I1(n23044[3]), .I2(n417), .I3(n53905), 
            .O(n22974[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5525_6 (.CI(n53905), .I0(n23044[3]), .I1(n417), .CO(n53906));
    SB_LUT4 add_5525_5_lut (.I0(GND_net), .I1(n23044[2]), .I2(n344), .I3(n53904), 
            .O(n22974[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5525_5 (.CI(n53904), .I0(n23044[2]), .I1(n344), .CO(n53905));
    SB_LUT4 counter_2046_2047_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n53447), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5525_4_lut (.I0(GND_net), .I1(n23044[1]), .I2(n271), .I3(n53903), 
            .O(n22974[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5525_4 (.CI(n53903), .I0(n23044[1]), .I1(n271), .CO(n53904));
    SB_LUT4 counter_2046_2047_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n53446), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_14 (.CI(n53446), .I0(GND_net), .I1(counter[12]), 
            .CO(n53447));
    SB_LUT4 add_5525_3_lut (.I0(GND_net), .I1(n23044[0]), .I2(n198), .I3(n53902), 
            .O(n22974[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5525_3 (.CI(n53902), .I0(n23044[0]), .I1(n198), .CO(n53903));
    SB_LUT4 counter_2046_2047_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n53445), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_13 (.CI(n53445), .I0(GND_net), .I1(counter[11]), 
            .CO(n53446));
    SB_LUT4 add_5525_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n22974[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5525_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5525_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n53902));
    SB_LUT4 counter_2046_2047_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n53444), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_12 (.CI(n53444), .I0(GND_net), .I1(counter[10]), 
            .CO(n53445));
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5476_10_lut (.I0(GND_net), .I1(n22692[7]), .I2(n700_adj_4546), 
            .I3(n53901), .O(n22496[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_10 (.CI(n52864), .I0(n21578[7]), .I1(n688_adj_4545), 
            .CO(n52865));
    SB_LUT4 add_5476_9_lut (.I0(GND_net), .I1(n22692[6]), .I2(n627_adj_4547), 
            .I3(n53900), .O(n22496[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5476_9 (.CI(n53900), .I0(n22692[6]), .I1(n627_adj_4547), 
            .CO(n53901));
    SB_LUT4 add_5476_8_lut (.I0(GND_net), .I1(n22692[5]), .I2(n554_adj_4548), 
            .I3(n53899), .O(n22496[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_9_lut (.I0(GND_net), .I1(n21578[6]), .I2(n615_adj_4549), 
            .I3(n52863), .O(n21080[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5476_8 (.CI(n53899), .I0(n22692[5]), .I1(n554_adj_4548), 
            .CO(n53900));
    SB_LUT4 counter_2046_2047_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n53443), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_11 (.CI(n53443), .I0(GND_net), .I1(counter[9]), 
            .CO(n53444));
    SB_CARRY add_5374_9 (.CI(n52863), .I0(n21578[6]), .I1(n615_adj_4549), 
            .CO(n52864));
    SB_LUT4 add_5374_8_lut (.I0(GND_net), .I1(n21578[5]), .I2(n542_adj_4550), 
            .I3(n52862), .O(n21080[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5476_7_lut (.I0(GND_net), .I1(n22692[4]), .I2(n481_adj_4551), 
            .I3(n53898), .O(n22496[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_8 (.CI(n52862), .I0(n21578[5]), .I1(n542_adj_4550), 
            .CO(n52863));
    SB_LUT4 add_5374_7_lut (.I0(GND_net), .I1(n21578[4]), .I2(n469_adj_4552), 
            .I3(n52861), .O(n21080[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_7 (.CI(n52861), .I0(n21578[4]), .I1(n469_adj_4552), 
            .CO(n52862));
    SB_LUT4 add_5374_6_lut (.I0(GND_net), .I1(n21578[3]), .I2(n396_adj_4553), 
            .I3(n52860), .O(n21080[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_6 (.CI(n52860), .I0(n21578[3]), .I1(n396_adj_4553), 
            .CO(n52861));
    SB_LUT4 add_5374_5_lut (.I0(GND_net), .I1(n21578[2]), .I2(n323_adj_4554), 
            .I3(n52859), .O(n21080[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_5 (.CI(n52859), .I0(n21578[2]), .I1(n323_adj_4554), 
            .CO(n52860));
    SB_LUT4 add_5374_4_lut (.I0(GND_net), .I1(n21578[1]), .I2(n250_adj_4555), 
            .I3(n52858), .O(n21080[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5476_7 (.CI(n53898), .I0(n22692[4]), .I1(n481_adj_4551), 
            .CO(n53899));
    SB_LUT4 add_5476_6_lut (.I0(GND_net), .I1(n22692[3]), .I2(n408_adj_4556), 
            .I3(n53897), .O(n22496[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2046_2047_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n53442), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_10 (.CI(n53442), .I0(GND_net), .I1(counter[8]), 
            .CO(n53443));
    SB_CARRY add_5476_6 (.CI(n53897), .I0(n22692[3]), .I1(n408_adj_4556), 
            .CO(n53898));
    SB_CARRY add_5374_4 (.CI(n52858), .I0(n21578[1]), .I1(n250_adj_4555), 
            .CO(n52859));
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4514));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5476_5_lut (.I0(GND_net), .I1(n22692[2]), .I2(n335_adj_4557), 
            .I3(n53896), .O(n22496[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2046_2047_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n53441), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4513));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5476_5 (.CI(n53896), .I0(n22692[2]), .I1(n335_adj_4557), 
            .CO(n53897));
    SB_LUT4 add_5476_4_lut (.I0(GND_net), .I1(n22692[1]), .I2(n262_adj_4558), 
            .I3(n53895), .O(n22496[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5476_4 (.CI(n53895), .I0(n22692[1]), .I1(n262_adj_4558), 
            .CO(n53896));
    SB_CARRY counter_2046_2047_add_4_9 (.CI(n53441), .I0(GND_net), .I1(counter[7]), 
            .CO(n53442));
    SB_LUT4 counter_2046_2047_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n53440), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5374_3_lut (.I0(GND_net), .I1(n21578[0]), .I2(n177_adj_4559), 
            .I3(n52857), .O(n21080[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5476_3_lut (.I0(GND_net), .I1(n22692[0]), .I2(n189_adj_4560), 
            .I3(n53894), .O(n22496[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5476_3 (.CI(n53894), .I0(n22692[0]), .I1(n189_adj_4560), 
            .CO(n53895));
    SB_CARRY add_5374_3 (.CI(n52857), .I0(n21578[0]), .I1(n177_adj_4559), 
            .CO(n52858));
    SB_LUT4 add_5476_2_lut (.I0(GND_net), .I1(n47_adj_4561), .I2(n116_adj_4562), 
            .I3(GND_net), .O(n22496[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5476_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_8 (.CI(n53440), .I0(GND_net), .I1(counter[6]), 
            .CO(n53441));
    SB_CARRY add_5476_2 (.CI(GND_net), .I0(n47_adj_4561), .I1(n116_adj_4562), 
            .CO(n53894));
    SB_LUT4 add_5374_2_lut (.I0(GND_net), .I1(n35_adj_4563), .I2(n104_adj_4564), 
            .I3(GND_net), .O(n21080[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5374_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5374_2 (.CI(GND_net), .I0(n35_adj_4563), .I1(n104_adj_4564), 
            .CO(n52857));
    SB_LUT4 counter_2046_2047_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n53439), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5406_13_lut (.I0(GND_net), .I1(n21974[10]), .I2(n910), 
            .I3(n52856), .O(n21578[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5493_9_lut (.I0(GND_net), .I1(n22833[6]), .I2(n630_adj_4565), 
            .I3(n53893), .O(n22692[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_7 (.CI(n53439), .I0(GND_net), .I1(counter[5]), 
            .CO(n53440));
    SB_LUT4 counter_2046_2047_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n53438), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5406_12_lut (.I0(GND_net), .I1(n21974[9]), .I2(n837), 
            .I3(n52855), .O(n21578[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5493_8_lut (.I0(GND_net), .I1(n22833[5]), .I2(n557_adj_4566), 
            .I3(n53892), .O(n22692[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5493_8 (.CI(n53892), .I0(n22833[5]), .I1(n557_adj_4566), 
            .CO(n53893));
    SB_LUT4 add_5493_7_lut (.I0(GND_net), .I1(n22833[4]), .I2(n484_adj_4567), 
            .I3(n53891), .O(n22692[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_6 (.CI(n53438), .I0(GND_net), .I1(counter[4]), 
            .CO(n53439));
    SB_CARRY add_5406_12 (.CI(n52855), .I0(n21974[9]), .I1(n837), .CO(n52856));
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5406_11_lut (.I0(GND_net), .I1(n21974[8]), .I2(n764), 
            .I3(n52854), .O(n21578[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2046_2047_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n53437), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5493_7 (.CI(n53891), .I0(n22833[4]), .I1(n484_adj_4567), 
            .CO(n53892));
    SB_LUT4 add_5493_6_lut (.I0(GND_net), .I1(n22833[3]), .I2(n411_adj_4568), 
            .I3(n53890), .O(n22692[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_5 (.CI(n53437), .I0(GND_net), .I1(counter[3]), 
            .CO(n53438));
    SB_LUT4 counter_2046_2047_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n53436), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4511));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5493_6 (.CI(n53890), .I0(n22833[3]), .I1(n411_adj_4568), 
            .CO(n53891));
    SB_LUT4 add_5493_5_lut (.I0(GND_net), .I1(n22833[2]), .I2(n338_adj_4569), 
            .I3(n53889), .O(n22692[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_4 (.CI(n53436), .I0(GND_net), .I1(counter[2]), 
            .CO(n53437));
    SB_LUT4 counter_2046_2047_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n53435), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5406_11 (.CI(n52854), .I0(n21974[8]), .I1(n764), .CO(n52855));
    SB_CARRY add_5493_5 (.CI(n53889), .I0(n22833[2]), .I1(n338_adj_4569), 
            .CO(n53890));
    SB_CARRY counter_2046_2047_add_4_3 (.CI(n53435), .I0(GND_net), .I1(counter[1]), 
            .CO(n53436));
    SB_LUT4 add_5493_4_lut (.I0(GND_net), .I1(n22833[1]), .I2(n265_adj_4570), 
            .I3(n53888), .O(n22692[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2046_2047_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2046_2047_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2046_2047_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n53435));
    SB_CARRY add_5493_4 (.CI(n53888), .I0(n22833[1]), .I1(n265_adj_4570), 
            .CO(n53889));
    SB_LUT4 add_5493_3_lut (.I0(GND_net), .I1(n22833[0]), .I2(n192_adj_4571), 
            .I3(n53887), .O(n22692[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5406_10_lut (.I0(GND_net), .I1(n21974[7]), .I2(n691), 
            .I3(n52853), .O(n21578[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5493_3 (.CI(n53887), .I0(n22833[0]), .I1(n192_adj_4571), 
            .CO(n53888));
    SB_LUT4 add_5493_2_lut (.I0(GND_net), .I1(n50_adj_4572), .I2(n119_adj_4573), 
            .I3(GND_net), .O(n22692[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5493_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n71311), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_5493_2 (.CI(GND_net), .I0(n50_adj_4572), .I1(n119_adj_4573), 
            .CO(n53887));
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5406_10 (.CI(n52853), .I0(n21974[7]), .I1(n691), .CO(n52854));
    SB_LUT4 add_5406_9_lut (.I0(GND_net), .I1(n21974[6]), .I2(n618), .I3(n52852), 
            .O(n21578[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5406_9 (.CI(n52852), .I0(n21974[6]), .I1(n618), .CO(n52853));
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4510));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5406_8_lut (.I0(GND_net), .I1(n21974[5]), .I2(n545), .I3(n52851), 
            .O(n21578[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4509));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n71293), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n71287), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n71281), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n71275), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n71269), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n71263), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n71257), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n71251), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n71245), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n71239), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_5406_8 (.CI(n52851), .I0(n21974[5]), .I1(n545), .CO(n52852));
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n71233), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n71227), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n71221), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n71215), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n71209), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n71683), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n71677), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_5406_7_lut (.I0(GND_net), .I1(n21974[4]), .I2(n472), .I3(n52850), 
            .O(n21578[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n71671), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_5406_7 (.CI(n52850), .I0(n21974[4]), .I1(n472), .CO(n52851));
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n71665), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n71659), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n71653), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_5406_6_lut (.I0(GND_net), .I1(n21974[3]), .I2(n399), .I3(n52849), 
            .O(n21578[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4508));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4507));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5406_6 (.CI(n52849), .I0(n21974[3]), .I1(n399), .CO(n52850));
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4506));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4505));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4504));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5406_5_lut (.I0(GND_net), .I1(n21974[2]), .I2(n326_adj_4574), 
            .I3(n52848), .O(n21578[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4503));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5406_5 (.CI(n52848), .I0(n21974[2]), .I1(n326_adj_4574), 
            .CO(n52849));
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4502));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4501));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4500));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4499));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4498));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4493));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4492));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4491));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4489));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9980_bdd_4_lut_52290 (.I0(n9980), .I1(n67744), .I2(setpoint[23]), 
            .I3(n4751), .O(n71488));
    defparam n9980_bdd_4_lut_52290.LUT_INIT = 16'he4aa;
    SB_LUT4 n71488_bdd_4_lut (.I0(n71488), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4751), .O(n71491));
    defparam n71488_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5406_4_lut (.I0(GND_net), .I1(n21974[1]), .I2(n253), .I3(n52847), 
            .O(n21578[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5406_4 (.CI(n52847), .I0(n21974[1]), .I1(n253), .CO(n52848));
    SB_LUT4 add_5406_3_lut (.I0(GND_net), .I1(n21974[0]), .I2(n180), .I3(n52846), 
            .O(n21578[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5406_3 (.CI(n52846), .I0(n21974[0]), .I1(n180), .CO(n52847));
    SB_LUT4 add_5406_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n21578[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5406_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n52846));
    SB_LUT4 add_5513_8_lut (.I0(GND_net), .I1(n22974[5]), .I2(n560), .I3(n52845), 
            .O(n22878[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5513_7_lut (.I0(GND_net), .I1(n22974[4]), .I2(n487), .I3(n52844), 
            .O(n22878[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_7 (.CI(n52844), .I0(n22974[4]), .I1(n487), .CO(n52845));
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4488));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4485));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4484));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4483));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5513_6_lut (.I0(GND_net), .I1(n22974[3]), .I2(n414), .I3(n52843), 
            .O(n22878[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_6 (.CI(n52843), .I0(n22974[3]), .I1(n414), .CO(n52844));
    SB_LUT4 add_5513_5_lut (.I0(GND_net), .I1(n22974[2]), .I2(n341), .I3(n52842), 
            .O(n22878[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_5 (.CI(n52842), .I0(n22974[2]), .I1(n341), .CO(n52843));
    SB_LUT4 add_5513_4_lut (.I0(GND_net), .I1(n22974[1]), .I2(n268), .I3(n52841), 
            .O(n22878[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_4 (.CI(n52841), .I0(n22974[1]), .I1(n268), .CO(n52842));
    SB_LUT4 add_5513_3_lut (.I0(GND_net), .I1(n22974[0]), .I2(n195), .I3(n52840), 
            .O(n22878[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_3 (.CI(n52840), .I0(n22974[0]), .I1(n195), .CO(n52841));
    SB_LUT4 add_5513_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n22878[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5513_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5513_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n52840));
    SB_LUT4 add_5433_12_lut (.I0(GND_net), .I1(n22278[9]), .I2(n840_adj_4575), 
            .I3(n52839), .O(n21974[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5433_11_lut (.I0(GND_net), .I1(n22278[8]), .I2(n767_adj_4576), 
            .I3(n52838), .O(n21974[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_11 (.CI(n52838), .I0(n22278[8]), .I1(n767_adj_4576), 
            .CO(n52839));
    SB_LUT4 add_5433_10_lut (.I0(GND_net), .I1(n22278[7]), .I2(n694_adj_4577), 
            .I3(n52837), .O(n21974[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_10 (.CI(n52837), .I0(n22278[7]), .I1(n694_adj_4577), 
            .CO(n52838));
    SB_LUT4 add_5433_9_lut (.I0(GND_net), .I1(n22278[6]), .I2(n621_adj_4578), 
            .I3(n52836), .O(n21974[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_9 (.CI(n52836), .I0(n22278[6]), .I1(n621_adj_4578), 
            .CO(n52837));
    SB_LUT4 add_5433_8_lut (.I0(GND_net), .I1(n22278[5]), .I2(n548_adj_4579), 
            .I3(n52835), .O(n21974[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5433_8 (.CI(n52835), .I0(n22278[5]), .I1(n548_adj_4579), 
            .CO(n52836));
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4479));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i11_3_lut (.I0(n233[10]), .I1(n285[10]), .I2(n284), 
            .I3(GND_net), .O(n310[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4478));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i11_3_lut (.I0(n310[10]), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n335[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4538));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4537));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4536));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(n70449), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n27506), .O(n27508));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff71;
    SB_LUT4 i1_2_lut_4_lut_adj_969 (.I0(n70449), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n27506), .O(n4));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_969.LUT_INIT = 16'hff8e;
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4476));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4535));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5433_7_lut (.I0(GND_net), .I1(n22278[4]), .I2(n475_adj_4581), 
            .I3(n52834), .O(n21974[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_7 (.CI(n52834), .I0(n22278[4]), .I1(n475_adj_4581), 
            .CO(n52835));
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4475));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n32332), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n32331), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n32330), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n32329), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n32328), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n32327), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n32326), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n32325), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n32324), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n32323), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n32322), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n32321), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n32320), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n32319), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n32318), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n32317), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n32316), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n32315), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n32314), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n32313), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n32312), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n32311), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n32308), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_5433_6_lut (.I0(GND_net), .I1(n22278[3]), .I2(n402_adj_4582), 
            .I3(n52833), .O(n21974[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4474));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5433_6 (.CI(n52833), .I0(n22278[3]), .I1(n402_adj_4582), 
            .CO(n52834));
    SB_LUT4 add_5433_5_lut (.I0(GND_net), .I1(n22278[2]), .I2(n329_adj_4583), 
            .I3(n52832), .O(n21974[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_5 (.CI(n52832), .I0(n22278[2]), .I1(n329_adj_4583), 
            .CO(n52833));
    SB_LUT4 add_5433_4_lut (.I0(GND_net), .I1(n22278[1]), .I2(n256_adj_4584), 
            .I3(n52831), .O(n21974[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_4 (.CI(n52831), .I0(n22278[1]), .I1(n256_adj_4584), 
            .CO(n52832));
    SB_LUT4 add_5433_3_lut (.I0(GND_net), .I1(n22278[0]), .I2(n183_adj_4585), 
            .I3(n52830), .O(n21974[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_3 (.CI(n52830), .I0(n22278[0]), .I1(n183_adj_4585), 
            .CO(n52831));
    SB_LUT4 add_5433_2_lut (.I0(GND_net), .I1(n41_adj_4586), .I2(n110_adj_4587), 
            .I3(GND_net), .O(n21974[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5433_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5433_2 (.CI(GND_net), .I0(n41_adj_4586), .I1(n110_adj_4587), 
            .CO(n52830));
    SB_LUT4 add_5456_11_lut (.I0(GND_net), .I1(n22496[8]), .I2(n770), 
            .I3(n52829), .O(n22278[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5456_10_lut (.I0(GND_net), .I1(n22496[7]), .I2(n697), 
            .I3(n52828), .O(n22278[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_10 (.CI(n52828), .I0(n22496[7]), .I1(n697), .CO(n52829));
    SB_LUT4 add_5456_9_lut (.I0(GND_net), .I1(n22496[6]), .I2(n624), .I3(n52827), 
            .O(n22278[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_9 (.CI(n52827), .I0(n22496[6]), .I1(n624), .CO(n52828));
    SB_LUT4 i48848_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(PWMLimit[2]), .O(n68118));   // verilog/motorControl.v(63[16:31])
    defparam i48848_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5456_8_lut (.I0(GND_net), .I1(n22496[5]), .I2(n551), .I3(n52826), 
            .O(n22278[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_8 (.CI(n52826), .I0(n22496[5]), .I1(n551), .CO(n52827));
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_5456_7_lut (.I0(GND_net), .I1(n22496[4]), .I2(n478_adj_4588), 
            .I3(n52825), .O(n22278[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n10812[0]), .I2(n10020[0]), 
            .I3(n52629), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_7 (.CI(n52825), .I0(n22496[4]), .I1(n478_adj_4588), 
            .CO(n52826));
    SB_LUT4 add_5456_6_lut (.I0(GND_net), .I1(n22496[3]), .I2(n405), .I3(n52824), 
            .O(n22278[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5456_6 (.CI(n52824), .I0(n22496[3]), .I1(n405), .CO(n52825));
    SB_LUT4 add_5456_5_lut (.I0(GND_net), .I1(n22496[2]), .I2(n332), .I3(n52823), 
            .O(n22278[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5456_5 (.CI(n52823), .I0(n22496[2]), .I1(n332), .CO(n52824));
    SB_LUT4 add_5456_4_lut (.I0(GND_net), .I1(n22496[1]), .I2(n259), .I3(n52822), 
            .O(n22278[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n36[22]), 
            .I3(n52628), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_24 (.CI(n52628), .I0(n360[22]), .I1(n36[22]), .CO(n52629));
    SB_DFFSR counter_2046_2047__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY add_5456_4 (.CI(n52822), .I0(n22496[1]), .I1(n259), .CO(n52823));
    SB_LUT4 add_5456_3_lut (.I0(GND_net), .I1(n22496[0]), .I2(n186), .I3(n52821), 
            .O(n22278[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_2046_2047__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2046_2047__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY add_5456_3 (.CI(n52821), .I0(n22496[0]), .I1(n186), .CO(n52822));
    SB_LUT4 add_5456_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n22278[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5456_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n31436), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5456_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n52821));
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n36[21]), 
            .I3(n52627), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n52627), .I0(n360[21]), .I1(n36[21]), .CO(n52628));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n36[20]), 
            .I3(n52626), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n52626), .I0(n360[20]), .I1(n36[20]), .CO(n52627));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n36[19]), 
            .I3(n52625), .O(n455[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5508_8_lut (.I0(GND_net), .I1(n22942[5]), .I2(n560_adj_4592), 
            .I3(n53773), .O(n22833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5508_7_lut (.I0(GND_net), .I1(n22942[4]), .I2(n487_adj_4593), 
            .I3(n53772), .O(n22833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n52625), .I0(n360[19]), .I1(n36[19]), .CO(n52626));
    SB_CARRY add_5508_7 (.CI(n53772), .I0(n22942[4]), .I1(n487_adj_4593), 
            .CO(n53773));
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n36[18]), 
            .I3(n52624), .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n52624), .I0(n360[18]), .I1(n36[18]), .CO(n52625));
    SB_LUT4 add_5508_6_lut (.I0(GND_net), .I1(n22942[3]), .I2(n414_adj_4594), 
            .I3(n53771), .O(n22833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5508_6 (.CI(n53771), .I0(n22942[3]), .I1(n414_adj_4594), 
            .CO(n53772));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n36[17]), 
            .I3(n52623), .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5508_5_lut (.I0(GND_net), .I1(n22942[2]), .I2(n341_adj_4596), 
            .I3(n53770), .O(n22833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5508_5 (.CI(n53770), .I0(n22942[2]), .I1(n341_adj_4596), 
            .CO(n53771));
    SB_LUT4 add_5508_4_lut (.I0(GND_net), .I1(n22942[1]), .I2(n268_adj_4597), 
            .I3(n53769), .O(n22833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5508_4 (.CI(n53769), .I0(n22942[1]), .I1(n268_adj_4597), 
            .CO(n53770));
    SB_LUT4 add_5508_3_lut (.I0(GND_net), .I1(n22942[0]), .I2(n195_adj_4598), 
            .I3(n53768), .O(n22833[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5508_3 (.CI(n53768), .I0(n22942[0]), .I1(n195_adj_4598), 
            .CO(n53769));
    SB_LUT4 add_5508_2_lut (.I0(GND_net), .I1(n53_adj_4599), .I2(n122_adj_4600), 
            .I3(GND_net), .O(n22833[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5508_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5508_2 (.CI(GND_net), .I0(n53_adj_4599), .I1(n122_adj_4600), 
            .CO(n53768));
    SB_CARRY add_25_19 (.CI(n52623), .I0(n360[17]), .I1(n36[17]), .CO(n52624));
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n36[16]), 
            .I3(n52622), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n52622), .I0(n360[16]), .I1(n36[16]), .CO(n52623));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n36[15]), 
            .I3(n52621), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_17 (.CI(n52621), .I0(n360[15]), .I1(n36[15]), .CO(n52622));
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n36[14]), 
            .I3(n52620), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_16 (.CI(n52620), .I0(n360[14]), .I1(n36[14]), .CO(n52621));
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n36[13]), 
            .I3(n52619), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n52619), .I0(n360[13]), .I1(n36[13]), .CO(n52620));
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n36[12]), 
            .I3(n52618), .O(n455[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n52618), .I0(n360[12]), .I1(n36[12]), .CO(n52619));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n36[11]), 
            .I3(n52617), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n52617), .I0(n360[11]), .I1(n36[11]), .CO(n52618));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n36[10]), 
            .I3(n52616), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5416_13_lut (.I0(GND_net), .I1(n22091[10]), .I2(n910_adj_4606), 
            .I3(n53325), .O(n21718[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5416_12_lut (.I0(GND_net), .I1(n22091[9]), .I2(n837_adj_4607), 
            .I3(n53324), .O(n21718[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_12 (.CI(n53324), .I0(n22091[9]), .I1(n837_adj_4607), 
            .CO(n53325));
    SB_LUT4 add_5416_11_lut (.I0(GND_net), .I1(n22091[8]), .I2(n764_adj_4608), 
            .I3(n53323), .O(n21718[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_12 (.CI(n52616), .I0(n360[10]), .I1(n36[10]), .CO(n52617));
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n36[9]), .I3(n52615), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_11 (.CI(n52615), .I0(n360[9]), .I1(n36[9]), .CO(n52616));
    SB_CARRY add_5416_11 (.CI(n53323), .I0(n22091[8]), .I1(n764_adj_4608), 
            .CO(n53324));
    SB_LUT4 add_5416_10_lut (.I0(GND_net), .I1(n22091[7]), .I2(n691_adj_4609), 
            .I3(n53322), .O(n21718[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_10 (.CI(n53322), .I0(n22091[7]), .I1(n691_adj_4609), 
            .CO(n53323));
    SB_LUT4 add_5416_9_lut (.I0(GND_net), .I1(n22091[6]), .I2(n618_adj_4610), 
            .I3(n53321), .O(n21718[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_9 (.CI(n53321), .I0(n22091[6]), .I1(n618_adj_4610), 
            .CO(n53322));
    SB_LUT4 add_5416_8_lut (.I0(GND_net), .I1(n22091[5]), .I2(n545_adj_4611), 
            .I3(n53320), .O(n21718[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_8 (.CI(n53320), .I0(n22091[5]), .I1(n545_adj_4611), 
            .CO(n53321));
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n36[8]), .I3(n52614), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_10 (.CI(n52614), .I0(n360[8]), .I1(n36[8]), .CO(n52615));
    SB_LUT4 add_5416_7_lut (.I0(GND_net), .I1(n22091[4]), .I2(n472_adj_4613), 
            .I3(n53319), .O(n21718[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5464_11_lut (.I0(GND_net), .I1(n22573[8]), .I2(n770_adj_4614), 
            .I3(n53067), .O(n22374[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5464_10_lut (.I0(GND_net), .I1(n22573[7]), .I2(n697_adj_4615), 
            .I3(n53066), .O(n22374[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_7 (.CI(n53319), .I0(n22091[4]), .I1(n472_adj_4613), 
            .CO(n53320));
    SB_LUT4 add_5416_6_lut (.I0(GND_net), .I1(n22091[3]), .I2(n399_adj_4616), 
            .I3(n53318), .O(n21718[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_6 (.CI(n53318), .I0(n22091[3]), .I1(n399_adj_4616), 
            .CO(n53319));
    SB_LUT4 add_5416_5_lut (.I0(GND_net), .I1(n22091[2]), .I2(n326_adj_4617), 
            .I3(n53317), .O(n21718[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_5 (.CI(n53317), .I0(n22091[2]), .I1(n326_adj_4617), 
            .CO(n53318));
    SB_LUT4 add_5521_7_lut (.I0(GND_net), .I1(n62793), .I2(n490_adj_4618), 
            .I3(n53744), .O(n22942[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5521_6_lut (.I0(GND_net), .I1(n23023[3]), .I2(n417_adj_4619), 
            .I3(n53743), .O(n22942[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5416_4_lut (.I0(GND_net), .I1(n22091[1]), .I2(n253_adj_4620), 
            .I3(n53316), .O(n21718[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_6 (.CI(n53743), .I0(n23023[3]), .I1(n417_adj_4619), 
            .CO(n53744));
    SB_LUT4 add_5521_5_lut (.I0(GND_net), .I1(n23023[2]), .I2(n344_adj_4621), 
            .I3(n53742), .O(n22942[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_4 (.CI(n53316), .I0(n22091[1]), .I1(n253_adj_4620), 
            .CO(n53317));
    SB_LUT4 add_5416_3_lut (.I0(GND_net), .I1(n22091[0]), .I2(n180_adj_4622), 
            .I3(n53315), .O(n21718[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_5 (.CI(n53742), .I0(n23023[2]), .I1(n344_adj_4621), 
            .CO(n53743));
    SB_LUT4 add_5521_4_lut (.I0(GND_net), .I1(n23023[1]), .I2(n271_adj_4623), 
            .I3(n53741), .O(n22942[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_3 (.CI(n53315), .I0(n22091[0]), .I1(n180_adj_4622), 
            .CO(n53316));
    SB_LUT4 add_5416_2_lut (.I0(GND_net), .I1(n38_adj_4624), .I2(n107_adj_4625), 
            .I3(GND_net), .O(n21718[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5416_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n36[7]), .I3(n52613), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_4 (.CI(n53741), .I0(n23023[1]), .I1(n271_adj_4623), 
            .CO(n53742));
    SB_LUT4 add_5521_3_lut (.I0(GND_net), .I1(n23023[0]), .I2(n198_adj_4627), 
            .I3(n53740), .O(n22942[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_3 (.CI(n53740), .I0(n23023[0]), .I1(n198_adj_4627), 
            .CO(n53741));
    SB_LUT4 add_5521_2_lut (.I0(GND_net), .I1(n56_adj_4628), .I2(n125_adj_4629), 
            .I3(GND_net), .O(n22942[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5416_2 (.CI(GND_net), .I0(n38_adj_4624), .I1(n107_adj_4625), 
            .CO(n53315));
    SB_CARRY add_5521_2 (.CI(GND_net), .I0(n56_adj_4628), .I1(n125_adj_4629), 
            .CO(n53740));
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n11271[21]), .I2(GND_net), 
            .I3(n53739), .O(n10812[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n11271[20]), .I2(GND_net), 
            .I3(n53738), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n53738), .I0(n11271[20]), .I1(GND_net), 
            .CO(n53739));
    SB_CARRY add_5464_10 (.CI(n53066), .I0(n22573[7]), .I1(n697_adj_4615), 
            .CO(n53067));
    SB_LUT4 add_5464_9_lut (.I0(GND_net), .I1(n22573[6]), .I2(n624_adj_4630), 
            .I3(n53065), .O(n22374[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n11271[19]), .I2(GND_net), 
            .I3(n53737), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_9 (.CI(n53065), .I0(n22573[6]), .I1(n624_adj_4630), 
            .CO(n53066));
    SB_CARRY add_25_9 (.CI(n52613), .I0(n360[7]), .I1(n36[7]), .CO(n52614));
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n36[6]), .I3(n52612), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5464_8_lut (.I0(GND_net), .I1(n22573[5]), .I2(n551_adj_4631), 
            .I3(n53064), .O(n22374[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_8 (.CI(n52612), .I0(n360[6]), .I1(n36[6]), .CO(n52613));
    SB_CARRY mult_23_add_1221_22 (.CI(n53737), .I0(n11271[19]), .I1(GND_net), 
            .CO(n53738));
    SB_CARRY add_5464_8 (.CI(n53064), .I0(n22573[5]), .I1(n551_adj_4631), 
            .CO(n53065));
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n11271[18]), .I2(GND_net), 
            .I3(n53736), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n53736), .I0(n11271[18]), .I1(GND_net), 
            .CO(n53737));
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n11271[17]), .I2(GND_net), 
            .I3(n53735), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_20 (.CI(n53735), .I0(n11271[17]), .I1(GND_net), 
            .CO(n53736));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n11271[16]), .I2(GND_net), 
            .I3(n53734), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n53734), .I0(n11271[16]), .I1(GND_net), 
            .CO(n53735));
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n11271[15]), .I2(GND_net), 
            .I3(n53733), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_18 (.CI(n53733), .I0(n11271[15]), .I1(GND_net), 
            .CO(n53734));
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n11271[14]), .I2(GND_net), 
            .I3(n53732), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_17 (.CI(n53732), .I0(n11271[14]), .I1(GND_net), 
            .CO(n53733));
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n11271[13]), .I2(n1096), 
            .I3(n53731), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n53731), .I0(n11271[13]), .I1(n1096), 
            .CO(n53732));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n11271[12]), .I2(n1023), 
            .I3(n53730), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_15 (.CI(n53730), .I0(n11271[12]), .I1(n1023), 
            .CO(n53731));
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n11271[11]), .I2(n950), 
            .I3(n53729), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5464_7_lut (.I0(GND_net), .I1(n22573[4]), .I2(n478_adj_4632), 
            .I3(n53063), .O(n22374[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_14 (.CI(n53729), .I0(n11271[11]), .I1(n950), 
            .CO(n53730));
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n11271[10]), .I2(n877), 
            .I3(n53728), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_13 (.CI(n53728), .I0(n11271[10]), .I1(n877), 
            .CO(n53729));
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n11271[9]), .I2(n804), 
            .I3(n53727), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n36[5]), .I3(n52611), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_7 (.CI(n53063), .I0(n22573[4]), .I1(n478_adj_4632), 
            .CO(n53064));
    SB_CARRY add_25_7 (.CI(n52611), .I0(n360[5]), .I1(n36[5]), .CO(n52612));
    SB_LUT4 add_5464_6_lut (.I0(GND_net), .I1(n22573[3]), .I2(n405_adj_4634), 
            .I3(n53062), .O(n22374[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_12 (.CI(n53727), .I0(n11271[9]), .I1(n804), 
            .CO(n53728));
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n11271[8]), .I2(n731), 
            .I3(n53726), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_6 (.CI(n53062), .I0(n22573[3]), .I1(n405_adj_4634), 
            .CO(n53063));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n36[4]), .I3(n52610), 
            .O(n455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_11 (.CI(n53726), .I0(n11271[8]), .I1(n731), 
            .CO(n53727));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n11271[7]), .I2(n658), 
            .I3(n53725), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_10 (.CI(n53725), .I0(n11271[7]), .I1(n658), 
            .CO(n53726));
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n11271[6]), .I2(n585), 
            .I3(n53724), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n52610), .I0(n360[4]), .I1(n36[4]), .CO(n52611));
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n36[3]), .I3(n52609), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n53724), .I0(n11271[6]), .I1(n585), 
            .CO(n53725));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n11271[5]), .I2(n512), 
            .I3(n53723), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_8 (.CI(n53723), .I0(n11271[5]), .I1(n512), 
            .CO(n53724));
    SB_LUT4 add_5464_5_lut (.I0(GND_net), .I1(n22573[2]), .I2(n332_adj_4635), 
            .I3(n53061), .O(n22374[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_5 (.CI(n53061), .I0(n22573[2]), .I1(n332_adj_4635), 
            .CO(n53062));
    SB_LUT4 add_5464_4_lut (.I0(GND_net), .I1(n22573[1]), .I2(n259_adj_4636), 
            .I3(n53060), .O(n22374[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n11271[4]), .I2(n439_adj_4637), 
            .I3(n53722), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_7 (.CI(n53722), .I0(n11271[4]), .I1(n439_adj_4637), 
            .CO(n53723));
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n11271[3]), .I2(n366), 
            .I3(n53721), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n53721), .I0(n11271[3]), .I1(n366), 
            .CO(n53722));
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n11271[2]), .I2(n293), 
            .I3(n53720), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_5 (.CI(n53720), .I0(n11271[2]), .I1(n293), 
            .CO(n53721));
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n11271[1]), .I2(n220_adj_4638), 
            .I3(n53719), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_4 (.CI(n53060), .I0(n22573[1]), .I1(n259_adj_4636), 
            .CO(n53061));
    SB_LUT4 add_5464_3_lut (.I0(GND_net), .I1(n22573[0]), .I2(n186_adj_4639), 
            .I3(n53059), .O(n22374[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_4 (.CI(n53719), .I0(n11271[1]), .I1(n220_adj_4638), 
            .CO(n53720));
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n11271[0]), .I2(n147), 
            .I3(n53718), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_3 (.CI(n53718), .I0(n11271[0]), .I1(n147), 
            .CO(n53719));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5), .I2(n74_adj_4641), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5), .I1(n74_adj_4641), 
            .CO(n53718));
    SB_CARRY add_5464_3 (.CI(n53059), .I0(n22573[0]), .I1(n186_adj_4639), 
            .CO(n53060));
    SB_LUT4 add_4795_23_lut (.I0(GND_net), .I1(n13100[20]), .I2(GND_net), 
            .I3(n53696), .O(n11271[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5464_2_lut (.I0(GND_net), .I1(n44_adj_4642), .I2(n113_adj_4643), 
            .I3(GND_net), .O(n22374[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5464_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5464_2 (.CI(GND_net), .I0(n44_adj_4642), .I1(n113_adj_4643), 
            .CO(n53059));
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n335[23]), .I1(n10527[21]), .I2(GND_net), 
            .I3(n53058), .O(n10020[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4795_22_lut (.I0(GND_net), .I1(n13100[19]), .I2(GND_net), 
            .I3(n53695), .O(n11271[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n10527[20]), .I2(GND_net), 
            .I3(n53057), .O(n36[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4467));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_23 (.CI(n53057), .I0(n10527[20]), .I1(GND_net), 
            .CO(n53058));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n10527[19]), .I2(GND_net), 
            .I3(n53056), .O(n36[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_22 (.CI(n53056), .I0(n10527[19]), .I1(GND_net), 
            .CO(n53057));
    SB_CARRY add_4795_22 (.CI(n53695), .I0(n13100[19]), .I1(GND_net), 
            .CO(n53696));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n10527[18]), .I2(GND_net), 
            .I3(n53055), .O(n36[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_21 (.CI(n53055), .I0(n10527[18]), .I1(GND_net), 
            .CO(n53056));
    SB_LUT4 add_4795_21_lut (.I0(GND_net), .I1(n13100[18]), .I2(GND_net), 
            .I3(n53694), .O(n11271[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n10527[17]), .I2(GND_net), 
            .I3(n53054), .O(n36[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n53054), .I0(n10527[17]), .I1(GND_net), 
            .CO(n53055));
    SB_CARRY add_4795_21 (.CI(n53694), .I0(n13100[18]), .I1(GND_net), 
            .CO(n53695));
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n10527[16]), .I2(GND_net), 
            .I3(n53053), .O(n36[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_19 (.CI(n53053), .I0(n10527[16]), .I1(GND_net), 
            .CO(n53054));
    SB_CARRY add_25_5 (.CI(n52609), .I0(n360[3]), .I1(n36[3]), .CO(n52610));
    SB_LUT4 add_4795_20_lut (.I0(GND_net), .I1(n13100[17]), .I2(GND_net), 
            .I3(n53693), .O(n11271[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n10527[15]), .I2(GND_net), 
            .I3(n53052), .O(n36[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n36[2]), .I3(n52608), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_4 (.CI(n52608), .I0(n360[2]), .I1(n36[2]), .CO(n52609));
    SB_CARRY mult_24_add_1225_18 (.CI(n53052), .I0(n10527[15]), .I1(GND_net), 
            .CO(n53053));
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n10527[14]), .I2(GND_net), 
            .I3(n53051), .O(n36[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n36[1]), .I3(n52607), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_3 (.CI(n52607), .I0(n360[1]), .I1(n36[1]), .CO(n52608));
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n36[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_20 (.CI(n53693), .I0(n13100[17]), .I1(GND_net), 
            .CO(n53694));
    SB_CARRY mult_24_add_1225_17 (.CI(n53051), .I0(n10527[14]), .I1(GND_net), 
            .CO(n53052));
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n10527[13]), .I2(n1096_adj_4645), 
            .I3(n53050), .O(n36[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_19_lut (.I0(GND_net), .I1(n13100[16]), .I2(GND_net), 
            .I3(n53692), .O(n11271[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_16 (.CI(n53050), .I0(n10527[13]), .I1(n1096_adj_4645), 
            .CO(n53051));
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[23]), 
            .I3(n52775), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n10527[12]), .I2(n1023_adj_4646), 
            .I3(n53049), .O(n36[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[22]), 
            .I3(n52774), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_19 (.CI(n53692), .I0(n13100[16]), .I1(GND_net), 
            .CO(n53693));
    SB_LUT4 add_4795_18_lut (.I0(GND_net), .I1(n13100[15]), .I2(GND_net), 
            .I3(n53691), .O(n11271[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_18 (.CI(n53691), .I0(n13100[15]), .I1(GND_net), 
            .CO(n53692));
    SB_CARRY mult_24_add_1225_15 (.CI(n53049), .I0(n10527[12]), .I1(n1023_adj_4646), 
            .CO(n53050));
    SB_LUT4 add_4795_17_lut (.I0(GND_net), .I1(n13100[14]), .I2(GND_net), 
            .I3(n53690), .O(n11271[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n52774), .I0(GND_net), .I1(n1_adj_5012[22]), 
            .CO(n52775));
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n10527[11]), .I2(n950_adj_4647), 
            .I3(n53048), .O(n36[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[21]), 
            .I3(n52773), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_14 (.CI(n53048), .I0(n10527[11]), .I1(n950_adj_4647), 
            .CO(n53049));
    SB_CARRY unary_minus_33_add_3_23 (.CI(n52773), .I0(GND_net), .I1(n1_adj_5012[21]), 
            .CO(n52774));
    SB_CARRY add_4795_17 (.CI(n53690), .I0(n13100[14]), .I1(GND_net), 
            .CO(n53691));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n10527[10]), .I2(n877_adj_4649), 
            .I3(n53047), .O(n36[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n36[0]), .CO(n52607));
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[20]), 
            .I3(n52772), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_13 (.CI(n53047), .I0(n10527[10]), .I1(n877_adj_4649), 
            .CO(n53048));
    SB_CARRY unary_minus_33_add_3_22 (.CI(n52772), .I0(GND_net), .I1(n1_adj_5012[20]), 
            .CO(n52773));
    SB_LUT4 add_4795_16_lut (.I0(GND_net), .I1(n13100[13]), .I2(n1099), 
            .I3(n53689), .O(n11271[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n10527[9]), .I2(n804_adj_4652), 
            .I3(n53046), .O(n36[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[19]), 
            .I3(n52771), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n52771), .I0(GND_net), .I1(n1_adj_5012[19]), 
            .CO(n52772));
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n52606), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_12 (.CI(n53046), .I0(n10527[9]), .I1(n804_adj_4652), 
            .CO(n53047));
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n52605), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[18]), 
            .I3(n52770), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n10527[8]), .I2(n731_adj_4655), 
            .I3(n53045), .O(n36[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_24 (.CI(n52605), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n52606));
    SB_CARRY unary_minus_33_add_3_20 (.CI(n52770), .I0(GND_net), .I1(n1_adj_5012[18]), 
            .CO(n52771));
    SB_CARRY mult_24_add_1225_11 (.CI(n53045), .I0(n10527[8]), .I1(n731_adj_4655), 
            .CO(n53046));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[17]), 
            .I3(n52769), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n52769), .I0(GND_net), .I1(n1_adj_5012[17]), 
            .CO(n52770));
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n52604), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n10527[7]), .I2(n658_adj_4658), 
            .I3(n53044), .O(n36[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_16 (.CI(n53689), .I0(n13100[13]), .I1(n1099), .CO(n53690));
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[16]), 
            .I3(n52768), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n53044), .I0(n10527[7]), .I1(n658_adj_4658), 
            .CO(n53045));
    SB_CARRY add_16_23 (.CI(n52604), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n52605));
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n10527[6]), .I2(n585_adj_4659), 
            .I3(n53043), .O(n36[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_15_lut (.I0(GND_net), .I1(n13100[12]), .I2(n1026), 
            .I3(n53688), .O(n11271[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_9 (.CI(n53043), .I0(n10527[6]), .I1(n585_adj_4659), 
            .CO(n53044));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n10527[5]), .I2(n512_adj_4660), 
            .I3(n53042), .O(n36[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n53042), .I0(n10527[5]), .I1(n512_adj_4660), 
            .CO(n53043));
    SB_CARRY add_4795_15 (.CI(n53688), .I0(n13100[12]), .I1(n1026), .CO(n53689));
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n10527[4]), .I2(n439_adj_4661), 
            .I3(n53041), .O(n36[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n52768), .I0(GND_net), .I1(n1_adj_5012[16]), 
            .CO(n52769));
    SB_CARRY mult_24_add_1225_7 (.CI(n53041), .I0(n10527[4]), .I1(n439_adj_4661), 
            .CO(n53042));
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[15]), 
            .I3(n52767), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_14_lut (.I0(GND_net), .I1(n13100[11]), .I2(n953), 
            .I3(n53687), .O(n11271[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n10527[3]), .I2(n366_adj_4662), 
            .I3(n53040), .O(n36[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_6 (.CI(n53040), .I0(n10527[3]), .I1(n366_adj_4662), 
            .CO(n53041));
    SB_CARRY unary_minus_33_add_3_17 (.CI(n52767), .I0(GND_net), .I1(n1_adj_5012[15]), 
            .CO(n52768));
    SB_CARRY add_4795_14 (.CI(n53687), .I0(n13100[11]), .I1(n953), .CO(n53688));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n10527[2]), .I2(n293_adj_4663), 
            .I3(n53039), .O(n36[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[14]), 
            .I3(n52766), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_5 (.CI(n53039), .I0(n10527[2]), .I1(n293_adj_4663), 
            .CO(n53040));
    SB_CARRY unary_minus_33_add_3_16 (.CI(n52766), .I0(GND_net), .I1(n1_adj_5012[14]), 
            .CO(n52767));
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[13]), 
            .I3(n52765), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n10527[1]), .I2(n220_adj_4665), 
            .I3(n53038), .O(n36[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n52603), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_22 (.CI(n52603), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n52604));
    SB_LUT4 add_4795_13_lut (.I0(GND_net), .I1(n13100[10]), .I2(n880), 
            .I3(n53686), .O(n11271[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_4 (.CI(n53038), .I0(n10527[1]), .I1(n220_adj_4665), 
            .CO(n53039));
    SB_CARRY unary_minus_33_add_3_15 (.CI(n52765), .I0(GND_net), .I1(n1_adj_5012[13]), 
            .CO(n52766));
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[12]), 
            .I3(n52764), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_14 (.CI(n52764), .I0(GND_net), .I1(n1_adj_5012[12]), 
            .CO(n52765));
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n52602), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n52602), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n52603));
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n10527[0]), .I2(n147_adj_4667), 
            .I3(n53037), .O(n36[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[11]), 
            .I3(n52763), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n52763), .I0(GND_net), .I1(n1_adj_5012[11]), 
            .CO(n52764));
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[10]), 
            .I3(n52762), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n52601), .O(n233[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_20 (.CI(n52601), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n52602));
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n52600), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_13 (.CI(n53686), .I0(n13100[10]), .I1(n880), .CO(n53687));
    SB_LUT4 add_4795_12_lut (.I0(GND_net), .I1(n13100[9]), .I2(n807), 
            .I3(n53685), .O(n11271[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_12 (.CI(n53685), .I0(n13100[9]), .I1(n807), .CO(n53686));
    SB_CARRY mult_24_add_1225_3 (.CI(n53037), .I0(n10527[0]), .I1(n147_adj_4667), 
            .CO(n53038));
    SB_CARRY unary_minus_33_add_3_12 (.CI(n52762), .I0(GND_net), .I1(n1_adj_5012[10]), 
            .CO(n52763));
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4669), .I2(n74_adj_4670), 
            .I3(GND_net), .O(n36[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[9]), 
            .I3(n52761), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_11_lut (.I0(GND_net), .I1(n13100[8]), .I2(n734), 
            .I3(n53684), .O(n11271[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5_adj_4669), .I1(n74_adj_4670), 
            .CO(n53037));
    SB_CARRY unary_minus_33_add_3_11 (.CI(n52761), .I0(GND_net), .I1(n1_adj_5012[9]), 
            .CO(n52762));
    SB_LUT4 add_4514_23_lut (.I0(GND_net), .I1(n12521[20]), .I2(GND_net), 
            .I3(n53036), .O(n10527[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[8]), 
            .I3(n52760), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_11 (.CI(n53684), .I0(n13100[8]), .I1(n734), .CO(n53685));
    SB_LUT4 add_4514_22_lut (.I0(GND_net), .I1(n12521[19]), .I2(GND_net), 
            .I3(n53035), .O(n10527[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_10 (.CI(n52760), .I0(GND_net), .I1(n1_adj_5012[8]), 
            .CO(n52761));
    SB_CARRY add_4514_22 (.CI(n53035), .I0(n12521[19]), .I1(GND_net), 
            .CO(n53036));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[7]), 
            .I3(n52759), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n52759), .I0(GND_net), .I1(n1_adj_5012[7]), 
            .CO(n52760));
    SB_LUT4 add_4795_10_lut (.I0(GND_net), .I1(n13100[7]), .I2(n661), 
            .I3(n53683), .O(n11271[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_21_lut (.I0(GND_net), .I1(n12521[18]), .I2(GND_net), 
            .I3(n53034), .O(n10527[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[6]), 
            .I3(n52758), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_21 (.CI(n53034), .I0(n12521[18]), .I1(GND_net), 
            .CO(n53035));
    SB_CARRY unary_minus_33_add_3_8 (.CI(n52758), .I0(GND_net), .I1(n1_adj_5012[6]), 
            .CO(n52759));
    SB_LUT4 add_4514_20_lut (.I0(GND_net), .I1(n12521[17]), .I2(GND_net), 
            .I3(n53033), .O(n10527[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_10 (.CI(n53683), .I0(n13100[7]), .I1(n661), .CO(n53684));
    SB_LUT4 add_4795_9_lut (.I0(GND_net), .I1(n13100[6]), .I2(n588), .I3(n53682), 
            .O(n11271[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_20 (.CI(n53033), .I0(n12521[17]), .I1(GND_net), 
            .CO(n53034));
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[5]), 
            .I3(n52757), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n52757), .I0(GND_net), .I1(n1_adj_5012[5]), 
            .CO(n52758));
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[4]), 
            .I3(n52756), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_19 (.CI(n52600), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n52601));
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n52599), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_6 (.CI(n52756), .I0(GND_net), .I1(n1_adj_5012[4]), 
            .CO(n52757));
    SB_CARRY add_4795_9 (.CI(n53682), .I0(n13100[6]), .I1(n588), .CO(n53683));
    SB_CARRY add_16_18 (.CI(n52599), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n52600));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n52598), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_8_lut (.I0(GND_net), .I1(n13100[5]), .I2(n515), .I3(n53681), 
            .O(n11271[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_19_lut (.I0(GND_net), .I1(n12521[16]), .I2(GND_net), 
            .I3(n53032), .O(n10527[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[3]), 
            .I3(n52755), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_8 (.CI(n53681), .I0(n13100[5]), .I1(n515), .CO(n53682));
    SB_CARRY add_4514_19 (.CI(n53032), .I0(n12521[16]), .I1(GND_net), 
            .CO(n53033));
    SB_CARRY unary_minus_33_add_3_5 (.CI(n52755), .I0(GND_net), .I1(n1_adj_5012[3]), 
            .CO(n52756));
    SB_LUT4 add_4514_18_lut (.I0(GND_net), .I1(n12521[15]), .I2(GND_net), 
            .I3(n53031), .O(n10527[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[2]), 
            .I3(n52754), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_7_lut (.I0(GND_net), .I1(n13100[4]), .I2(n442_adj_4676), 
            .I3(n53680), .O(n11271[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_18 (.CI(n53031), .I0(n12521[15]), .I1(GND_net), 
            .CO(n53032));
    SB_CARRY unary_minus_33_add_3_4 (.CI(n52754), .I0(GND_net), .I1(n1_adj_5012[2]), 
            .CO(n52755));
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[1]), 
            .I3(n52753), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_3 (.CI(n52753), .I0(GND_net), .I1(n1_adj_5012[1]), 
            .CO(n52754));
    SB_LUT4 add_4514_17_lut (.I0(GND_net), .I1(n12521[14]), .I2(GND_net), 
            .I3(n53030), .O(n10527[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5012[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_7 (.CI(n53680), .I0(n13100[4]), .I1(n442_adj_4676), 
            .CO(n53681));
    SB_CARRY add_4514_17 (.CI(n53030), .I0(n12521[14]), .I1(GND_net), 
            .CO(n53031));
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5012[0]), 
            .CO(n52753));
    SB_CARRY add_16_17 (.CI(n52598), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n52599));
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n52597), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_6_lut (.I0(GND_net), .I1(n13100[3]), .I2(n369), .I3(n53679), 
            .O(n11271[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_16_lut (.I0(GND_net), .I1(n12521[13]), .I2(n1099_adj_4677), 
            .I3(n53029), .O(n10527[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_5013[23]), 
            .I3(n52752), .O(n47_adj_4678)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4514_16 (.CI(n53029), .I0(n12521[13]), .I1(n1099_adj_4677), 
            .CO(n53030));
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[22]), 
            .I3(n52751), .O(n46[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_6 (.CI(n53679), .I0(n13100[3]), .I1(n369), .CO(n53680));
    SB_LUT4 add_4514_15_lut (.I0(GND_net), .I1(n12521[12]), .I2(n1026_adj_4681), 
            .I3(n53028), .O(n10527[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n52751), .I0(GND_net), .I1(n1_adj_5013[22]), 
            .CO(n52752));
    SB_CARRY add_4514_15 (.CI(n53028), .I0(n12521[12]), .I1(n1026_adj_4681), 
            .CO(n53029));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[21]), 
            .I3(n52750), .O(n46[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_5_lut (.I0(GND_net), .I1(n13100[2]), .I2(n296), .I3(n53678), 
            .O(n11271[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_5 (.CI(n53678), .I0(n13100[2]), .I1(n296), .CO(n53679));
    SB_CARRY add_16_16 (.CI(n52597), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n52598));
    SB_LUT4 add_4514_14_lut (.I0(GND_net), .I1(n12521[11]), .I2(n953_adj_4684), 
            .I3(n53027), .O(n10527[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n52750), .I0(GND_net), .I1(n1_adj_5013[21]), 
            .CO(n52751));
    SB_CARRY add_4514_14 (.CI(n53027), .I0(n12521[11]), .I1(n953_adj_4684), 
            .CO(n53028));
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[20]), 
            .I3(n52749), .O(n46[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4795_4_lut (.I0(GND_net), .I1(n13100[1]), .I2(n223_adj_4686), 
            .I3(n53677), .O(n11271[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_13_lut (.I0(GND_net), .I1(n12521[10]), .I2(n880_adj_4687), 
            .I3(n53026), .O(n10527[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_22 (.CI(n52749), .I0(GND_net), .I1(n1_adj_5013[20]), 
            .CO(n52750));
    SB_CARRY add_4514_13 (.CI(n53026), .I0(n12521[10]), .I1(n880_adj_4687), 
            .CO(n53027));
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[19]), 
            .I3(n52748), .O(n46[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_4 (.CI(n53677), .I0(n13100[1]), .I1(n223_adj_4686), 
            .CO(n53678));
    SB_LUT4 add_4795_3_lut (.I0(GND_net), .I1(n13100[0]), .I2(n150), .I3(n53676), 
            .O(n11271[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_12_lut (.I0(GND_net), .I1(n12521[9]), .I2(n807_adj_4689), 
            .I3(n53025), .O(n10527[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_21 (.CI(n52748), .I0(GND_net), .I1(n1_adj_5013[19]), 
            .CO(n52749));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[18]), 
            .I3(n52747), .O(n46[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n52596), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_15 (.CI(n52596), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n52597));
    SB_CARRY add_4514_12 (.CI(n53025), .I0(n12521[9]), .I1(n807_adj_4689), 
            .CO(n53026));
    SB_CARRY unary_minus_27_add_3_20 (.CI(n52747), .I0(GND_net), .I1(n1_adj_5013[18]), 
            .CO(n52748));
    SB_LUT4 add_4514_11_lut (.I0(GND_net), .I1(n12521[8]), .I2(n734_adj_4693), 
            .I3(n53024), .O(n10527[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[17]), 
            .I3(n52746), .O(n46[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_11 (.CI(n53024), .I0(n12521[8]), .I1(n734_adj_4693), 
            .CO(n53025));
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n52595), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n52746), .I0(GND_net), .I1(n1_adj_5013[17]), 
            .CO(n52747));
    SB_CARRY add_16_14 (.CI(n52595), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n52596));
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n52594), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_10_lut (.I0(GND_net), .I1(n12521[7]), .I2(n661_adj_4695), 
            .I3(n53023), .O(n10527[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[16]), 
            .I3(n52745), .O(n46[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_10 (.CI(n53023), .I0(n12521[7]), .I1(n661_adj_4695), 
            .CO(n53024));
    SB_CARRY unary_minus_27_add_3_18 (.CI(n52745), .I0(GND_net), .I1(n1_adj_5013[16]), 
            .CO(n52746));
    SB_CARRY add_4795_3 (.CI(n53676), .I0(n13100[0]), .I1(n150), .CO(n53677));
    SB_LUT4 add_4514_9_lut (.I0(GND_net), .I1(n12521[6]), .I2(n588_adj_4697), 
            .I3(n53022), .O(n10527[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[15]), 
            .I3(n52744), .O(n46[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_9 (.CI(n53022), .I0(n12521[6]), .I1(n588_adj_4697), 
            .CO(n53023));
    SB_CARRY unary_minus_27_add_3_17 (.CI(n52744), .I0(GND_net), .I1(n1_adj_5013[15]), 
            .CO(n52745));
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[14]), 
            .I3(n52743), .O(n46[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_13 (.CI(n52594), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n52595));
    SB_LUT4 add_4795_2_lut (.I0(GND_net), .I1(n8_adj_4701), .I2(n77), 
            .I3(GND_net), .O(n11271[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4795_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_8_lut (.I0(GND_net), .I1(n12521[5]), .I2(n515_adj_4702), 
            .I3(n53021), .O(n10527[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n52743), .I0(GND_net), .I1(n1_adj_5013[14]), 
            .CO(n52744));
    SB_CARRY add_4514_8 (.CI(n53021), .I0(n12521[5]), .I1(n515_adj_4702), 
            .CO(n53022));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[13]), 
            .I3(n52742), .O(n46[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4795_2 (.CI(GND_net), .I0(n8_adj_4701), .I1(n77), .CO(n53676));
    SB_LUT4 add_4514_7_lut (.I0(GND_net), .I1(n12521[4]), .I2(n442_adj_4704), 
            .I3(n53020), .O(n10527[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_15 (.CI(n52742), .I0(GND_net), .I1(n1_adj_5013[13]), 
            .CO(n52743));
    SB_CARRY add_4514_7 (.CI(n53020), .I0(n12521[4]), .I1(n442_adj_4704), 
            .CO(n53021));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[12]), 
            .I3(n52741), .O(n46[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_22_lut (.I0(GND_net), .I1(n14607[19]), .I2(GND_net), 
            .I3(n53675), .O(n13100[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4514_6_lut (.I0(GND_net), .I1(n12521[3]), .I2(n369_adj_4706), 
            .I3(n53019), .O(n10527[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n52741), .I0(GND_net), .I1(n1_adj_5013[12]), 
            .CO(n52742));
    SB_CARRY add_4514_6 (.CI(n53019), .I0(n12521[3]), .I1(n369_adj_4706), 
            .CO(n53020));
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[11]), 
            .I3(n52740), .O(n46[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_13 (.CI(n52740), .I0(GND_net), .I1(n1_adj_5013[11]), 
            .CO(n52741));
    SB_LUT4 add_4998_21_lut (.I0(GND_net), .I1(n14607[18]), .I2(GND_net), 
            .I3(n53674), .O(n13100[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_21 (.CI(n53674), .I0(n14607[18]), .I1(GND_net), 
            .CO(n53675));
    SB_LUT4 add_4514_5_lut (.I0(GND_net), .I1(n12521[2]), .I2(n296_adj_4708), 
            .I3(n53018), .O(n10527[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[10]), 
            .I3(n52739), .O(n46[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n52739), .I0(GND_net), .I1(n1_adj_5013[10]), 
            .CO(n52740));
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n52593), .O(n233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_12 (.CI(n52593), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n52594));
    SB_CARRY add_4514_5 (.CI(n53018), .I0(n12521[2]), .I1(n296_adj_4708), 
            .CO(n53019));
    SB_LUT4 add_4998_20_lut (.I0(GND_net), .I1(n14607[17]), .I2(GND_net), 
            .I3(n53673), .O(n13100[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_20 (.CI(n53673), .I0(n14607[17]), .I1(GND_net), 
            .CO(n53674));
    SB_LUT4 add_4514_4_lut (.I0(GND_net), .I1(n12521[1]), .I2(n223_adj_4710), 
            .I3(n53017), .O(n10527[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[9]), 
            .I3(n52738), .O(n46[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_11 (.CI(n52738), .I0(GND_net), .I1(n1_adj_5013[9]), 
            .CO(n52739));
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n52592), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n52592), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n52593));
    SB_CARRY add_4514_4 (.CI(n53017), .I0(n12521[1]), .I1(n223_adj_4710), 
            .CO(n53018));
    SB_LUT4 add_4514_3_lut (.I0(GND_net), .I1(n12521[0]), .I2(n150_adj_4712), 
            .I3(n53016), .O(n10527[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[8]), 
            .I3(n52737), .O(n46[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n52591), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_3 (.CI(n53016), .I0(n12521[0]), .I1(n150_adj_4712), 
            .CO(n53017));
    SB_CARRY unary_minus_27_add_3_10 (.CI(n52737), .I0(GND_net), .I1(n1_adj_5013[8]), 
            .CO(n52738));
    SB_LUT4 add_4514_2_lut (.I0(GND_net), .I1(n8_adj_4714), .I2(n77_adj_4715), 
            .I3(GND_net), .O(n10527[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4514_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[7]), 
            .I3(n52736), .O(n46[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n52736), .I0(GND_net), .I1(n1_adj_5013[7]), 
            .CO(n52737));
    SB_LUT4 add_4998_19_lut (.I0(GND_net), .I1(n14607[16]), .I2(GND_net), 
            .I3(n53672), .O(n13100[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4514_2 (.CI(GND_net), .I0(n8_adj_4714), .I1(n77_adj_4715), 
            .CO(n53016));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[6]), 
            .I3(n52735), .O(n46[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_22_lut (.I0(GND_net), .I1(n14096[19]), .I2(GND_net), 
            .I3(n53015), .O(n12521[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n52735), .I0(GND_net), .I1(n1_adj_5013[6]), 
            .CO(n52736));
    SB_CARRY add_4998_19 (.CI(n53672), .I0(n14607[16]), .I1(GND_net), 
            .CO(n53673));
    SB_LUT4 add_4998_18_lut (.I0(GND_net), .I1(n14607[15]), .I2(GND_net), 
            .I3(n53671), .O(n13100[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_21_lut (.I0(GND_net), .I1(n14096[18]), .I2(GND_net), 
            .I3(n53014), .O(n12521[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[5]), 
            .I3(n52734), .O(n46[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_21 (.CI(n53014), .I0(n14096[18]), .I1(GND_net), 
            .CO(n53015));
    SB_CARRY unary_minus_27_add_3_7 (.CI(n52734), .I0(GND_net), .I1(n1_adj_5013[5]), 
            .CO(n52735));
    SB_CARRY add_4998_18 (.CI(n53671), .I0(n14607[15]), .I1(GND_net), 
            .CO(n53672));
    SB_LUT4 add_4972_20_lut (.I0(GND_net), .I1(n14096[17]), .I2(GND_net), 
            .I3(n53013), .O(n12521[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[4]), 
            .I3(n52733), .O(n46[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_20 (.CI(n53013), .I0(n14096[17]), .I1(GND_net), 
            .CO(n53014));
    SB_LUT4 add_4998_17_lut (.I0(GND_net), .I1(n14607[14]), .I2(GND_net), 
            .I3(n53670), .O(n13100[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_19_lut (.I0(GND_net), .I1(n14096[16]), .I2(GND_net), 
            .I3(n53012), .O(n12521[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_17 (.CI(n53670), .I0(n14607[14]), .I1(GND_net), 
            .CO(n53671));
    SB_CARRY add_4972_19 (.CI(n53012), .I0(n14096[16]), .I1(GND_net), 
            .CO(n53013));
    SB_CARRY unary_minus_27_add_3_6 (.CI(n52733), .I0(GND_net), .I1(n1_adj_5013[4]), 
            .CO(n52734));
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[3]), 
            .I3(n52732), .O(n46[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_10 (.CI(n52591), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n52592));
    SB_LUT4 add_4998_16_lut (.I0(GND_net), .I1(n14607[13]), .I2(n1102), 
            .I3(n53669), .O(n13100[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_18_lut (.I0(GND_net), .I1(n14096[15]), .I2(GND_net), 
            .I3(n53011), .O(n12521[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n52590), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_18 (.CI(n53011), .I0(n14096[15]), .I1(GND_net), 
            .CO(n53012));
    SB_CARRY add_16_9 (.CI(n52590), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n52591));
    SB_LUT4 n9980_bdd_4_lut_52161 (.I0(n9980), .I1(n67600), .I2(setpoint[22]), 
            .I3(n4751), .O(n71308));
    defparam n9980_bdd_4_lut_52161.LUT_INIT = 16'he4aa;
    SB_CARRY add_4998_16 (.CI(n53669), .I0(n14607[13]), .I1(n1102), .CO(n53670));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n52589), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_17_lut (.I0(GND_net), .I1(n14096[14]), .I2(GND_net), 
            .I3(n53010), .O(n12521[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n52732), .I0(GND_net), .I1(n1_adj_5013[3]), 
            .CO(n52733));
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[2]), 
            .I3(n52731), .O(n46[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_15_lut (.I0(GND_net), .I1(n14607[12]), .I2(n1029), 
            .I3(n53668), .O(n13100[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_17 (.CI(n53010), .I0(n14096[14]), .I1(GND_net), 
            .CO(n53011));
    SB_CARRY unary_minus_27_add_3_4 (.CI(n52731), .I0(GND_net), .I1(n1_adj_5013[2]), 
            .CO(n52732));
    SB_LUT4 add_4972_16_lut (.I0(GND_net), .I1(n14096[13]), .I2(n1102_adj_4723), 
            .I3(n53009), .O(n12521[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5013[1]), 
            .I3(n52730), .O(n46[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n52730), .I0(GND_net), .I1(n1_adj_5013[1]), 
            .CO(n52731));
    SB_CARRY add_4998_15 (.CI(n53668), .I0(n14607[12]), .I1(n1029), .CO(n53669));
    SB_CARRY add_4972_16 (.CI(n53009), .I0(n14096[13]), .I1(n1102_adj_4723), 
            .CO(n53010));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n41898), .I1(GND_net), .I2(n1_adj_5013[0]), 
            .I3(VCC_net), .O(n67612)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5013[0]), 
            .CO(n52730));
    SB_LUT4 add_4972_15_lut (.I0(GND_net), .I1(n14096[12]), .I2(n1029_adj_4726), 
            .I3(n53008), .O(n12521[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[23]), 
            .I3(n52729), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[22]), 
            .I3(n52728), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_14_lut (.I0(GND_net), .I1(n14607[11]), .I2(n956), 
            .I3(n53667), .O(n13100[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_15 (.CI(n53008), .I0(n14096[12]), .I1(n1029_adj_4726), 
            .CO(n53009));
    SB_CARRY add_4998_14 (.CI(n53667), .I0(n14607[11]), .I1(n956), .CO(n53668));
    SB_LUT4 add_4998_13_lut (.I0(GND_net), .I1(n14607[10]), .I2(n883), 
            .I3(n53666), .O(n13100[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_14_lut (.I0(GND_net), .I1(n14096[11]), .I2(n956_adj_4729), 
            .I3(n53007), .O(n12521[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n52728), .I0(GND_net), .I1(n1_adj_5014[22]), 
            .CO(n52729));
    SB_CARRY add_4972_14 (.CI(n53007), .I0(n14096[11]), .I1(n956_adj_4729), 
            .CO(n53008));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[21]), 
            .I3(n52727), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_8 (.CI(n52589), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n52590));
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n52588), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_13_lut (.I0(GND_net), .I1(n14096[10]), .I2(n883_adj_4731), 
            .I3(n53006), .O(n12521[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n52727), .I0(GND_net), .I1(n1_adj_5014[21]), 
            .CO(n52728));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[20]), 
            .I3(n52726), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_7 (.CI(n52588), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n52589));
    SB_CARRY add_4972_13 (.CI(n53006), .I0(n14096[10]), .I1(n883_adj_4731), 
            .CO(n53007));
    SB_CARRY unary_minus_20_add_3_22 (.CI(n52726), .I0(GND_net), .I1(n1_adj_5014[20]), 
            .CO(n52727));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[19]), 
            .I3(n52725), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n52587), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_13 (.CI(n53666), .I0(n14607[10]), .I1(n883), .CO(n53667));
    SB_LUT4 add_4972_12_lut (.I0(GND_net), .I1(n14096[9]), .I2(n810), 
            .I3(n53005), .O(n12521[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n52725), .I0(GND_net), .I1(n1_adj_5014[19]), 
            .CO(n52726));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[18]), 
            .I3(n52724), .O(n285[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_12 (.CI(n53005), .I0(n14096[9]), .I1(n810), .CO(n53006));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n52724), .I0(GND_net), .I1(n1_adj_5014[18]), 
            .CO(n52725));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[17]), 
            .I3(n52723), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_6 (.CI(n52587), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n52588));
    SB_LUT4 add_4998_12_lut (.I0(GND_net), .I1(n14607[9]), .I2(n810_adj_4737), 
            .I3(n53665), .O(n13100[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_11_lut (.I0(GND_net), .I1(n14096[8]), .I2(n737), 
            .I3(n53004), .O(n12521[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n52723), .I0(GND_net), .I1(n1_adj_5014[17]), 
            .CO(n52724));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[16]), 
            .I3(n52722), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n52586), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_11 (.CI(n53004), .I0(n14096[8]), .I1(n737), .CO(n53005));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n52722), .I0(GND_net), .I1(n1_adj_5014[16]), 
            .CO(n52723));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[15]), 
            .I3(n52721), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_5 (.CI(n52586), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n52587));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n52585), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_12 (.CI(n53665), .I0(n14607[9]), .I1(n810_adj_4737), 
            .CO(n53666));
    SB_LUT4 add_4972_10_lut (.I0(GND_net), .I1(n14096[7]), .I2(n664), 
            .I3(n53003), .O(n12521[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n52721), .I0(GND_net), .I1(n1_adj_5014[15]), 
            .CO(n52722));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[14]), 
            .I3(n52720), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_4 (.CI(n52585), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n52586));
    SB_CARRY add_4972_10 (.CI(n53003), .I0(n14096[7]), .I1(n664), .CO(n53004));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n52720), .I0(GND_net), .I1(n1_adj_5014[14]), 
            .CO(n52721));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[13]), 
            .I3(n52719), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n52584), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_11_lut (.I0(GND_net), .I1(n14607[8]), .I2(n737_adj_4745), 
            .I3(n53664), .O(n13100[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_9_lut (.I0(GND_net), .I1(n14096[6]), .I2(n591), .I3(n53002), 
            .O(n12521[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n52719), .I0(GND_net), .I1(n1_adj_5014[13]), 
            .CO(n52720));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[12]), 
            .I3(n52718), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_3 (.CI(n52584), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n52585));
    SB_CARRY add_4972_9 (.CI(n53002), .I0(n14096[6]), .I1(n591), .CO(n53003));
    SB_CARRY unary_minus_20_add_3_14 (.CI(n52718), .I0(GND_net), .I1(n1_adj_5014[12]), 
            .CO(n52719));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[11]), 
            .I3(n52717), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_11 (.CI(n53664), .I0(n14607[8]), .I1(n737_adj_4745), 
            .CO(n53665));
    SB_LUT4 add_4972_8_lut (.I0(GND_net), .I1(n14096[5]), .I2(n518), .I3(n53001), 
            .O(n12521[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n52717), .I0(GND_net), .I1(n1_adj_5014[11]), 
            .CO(n52718));
    SB_LUT4 add_4998_10_lut (.I0(GND_net), .I1(n14607[7]), .I2(n664_adj_4748), 
            .I3(n53663), .O(n13100[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_8 (.CI(n53001), .I0(n14096[5]), .I1(n518), .CO(n53002));
    SB_CARRY add_4998_10 (.CI(n53663), .I0(n14607[7]), .I1(n664_adj_4748), 
            .CO(n53664));
    SB_LUT4 add_4972_7_lut (.I0(GND_net), .I1(n14096[4]), .I2(n445_adj_4749), 
            .I3(n53000), .O(n12521[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_7 (.CI(n53000), .I0(n14096[4]), .I1(n445_adj_4749), 
            .CO(n53001));
    SB_LUT4 add_4972_6_lut (.I0(GND_net), .I1(n14096[3]), .I2(n372), .I3(n52999), 
            .O(n12521[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_9_lut (.I0(GND_net), .I1(n14607[6]), .I2(n591_adj_4750), 
            .I3(n53662), .O(n13100[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_6 (.CI(n52999), .I0(n14096[3]), .I1(n372), .CO(n53000));
    SB_LUT4 add_4972_5_lut (.I0(GND_net), .I1(n14096[2]), .I2(n299_adj_4751), 
            .I3(n52998), .O(n12521[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_9 (.CI(n53662), .I0(n14607[6]), .I1(n591_adj_4750), 
            .CO(n53663));
    SB_CARRY add_4972_5 (.CI(n52998), .I0(n14096[2]), .I1(n299_adj_4751), 
            .CO(n52999));
    SB_LUT4 add_4998_8_lut (.I0(GND_net), .I1(n14607[5]), .I2(n518_adj_4752), 
            .I3(n53661), .O(n13100[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4972_4_lut (.I0(GND_net), .I1(n14096[1]), .I2(n226_adj_4753), 
            .I3(n52997), .O(n12521[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_4 (.CI(n52997), .I0(n14096[1]), .I1(n226_adj_4753), 
            .CO(n52998));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[10]), 
            .I3(n52716), .O(n285[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n52716), .I0(GND_net), .I1(n1_adj_5014[10]), 
            .CO(n52717));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[9]), 
            .I3(n52715), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n52584));
    SB_LUT4 add_4972_3_lut (.I0(GND_net), .I1(n14096[0]), .I2(n153), .I3(n52996), 
            .O(n12521[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n52715), .I0(GND_net), .I1(n1_adj_5014[9]), 
            .CO(n52716));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[8]), 
            .I3(n52714), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n52583), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n52582), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_3 (.CI(n52996), .I0(n14096[0]), .I1(n153), .CO(n52997));
    SB_CARRY add_4998_8 (.CI(n53661), .I0(n14607[5]), .I1(n518_adj_4752), 
            .CO(n53662));
    SB_LUT4 add_4972_2_lut (.I0(GND_net), .I1(n11_adj_4757), .I2(n80), 
            .I3(GND_net), .O(n12521[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n52714), .I0(GND_net), .I1(n1_adj_5014[8]), 
            .CO(n52715));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[7]), 
            .I3(n52713), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_7_lut (.I0(GND_net), .I1(n14607[4]), .I2(n445_adj_4759), 
            .I3(n53660), .O(n13100[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4972_2 (.CI(GND_net), .I0(n11_adj_4757), .I1(n80), .CO(n52996));
    SB_LUT4 add_5037_21_lut (.I0(GND_net), .I1(n15513[18]), .I2(GND_net), 
            .I3(n52995), .O(n14096[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_7 (.CI(n53660), .I0(n14607[4]), .I1(n445_adj_4759), 
            .CO(n53661));
    SB_CARRY sub_15_add_2_24 (.CI(n52582), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n52583));
    SB_LUT4 add_5037_20_lut (.I0(GND_net), .I1(n15513[17]), .I2(GND_net), 
            .I3(n52994), .O(n14096[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n52713), .I0(GND_net), .I1(n1_adj_5014[7]), 
            .CO(n52714));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[6]), 
            .I3(n52712), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n52581), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_23 (.CI(n52581), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n52582));
    SB_LUT4 add_4998_6_lut (.I0(GND_net), .I1(n14607[3]), .I2(n372_adj_4761), 
            .I3(n53659), .O(n13100[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_6 (.CI(n53659), .I0(n14607[3]), .I1(n372_adj_4761), 
            .CO(n53660));
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n52580), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_20 (.CI(n52994), .I0(n15513[17]), .I1(GND_net), 
            .CO(n52995));
    SB_CARRY unary_minus_20_add_3_8 (.CI(n52712), .I0(GND_net), .I1(n1_adj_5014[6]), 
            .CO(n52713));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[5]), 
            .I3(n52711), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_22 (.CI(n52580), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n52581));
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n52579), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_19_lut (.I0(GND_net), .I1(n15513[16]), .I2(GND_net), 
            .I3(n52993), .O(n14096[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n52711), .I0(GND_net), .I1(n1_adj_5014[5]), 
            .CO(n52712));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[4]), 
            .I3(n52710), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_21 (.CI(n52579), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n52580));
    SB_CARRY add_5037_19 (.CI(n52993), .I0(n15513[16]), .I1(GND_net), 
            .CO(n52994));
    SB_LUT4 add_5037_18_lut (.I0(GND_net), .I1(n15513[15]), .I2(GND_net), 
            .I3(n52992), .O(n14096[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_18 (.CI(n52992), .I0(n15513[15]), .I1(GND_net), 
            .CO(n52993));
    SB_LUT4 add_4998_5_lut (.I0(GND_net), .I1(n14607[2]), .I2(n299_adj_4765), 
            .I3(n53658), .O(n13100[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_17_lut (.I0(GND_net), .I1(n15513[14]), .I2(GND_net), 
            .I3(n52991), .O(n14096[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_17 (.CI(n52991), .I0(n15513[14]), .I1(GND_net), 
            .CO(n52992));
    SB_LUT4 add_5037_16_lut (.I0(GND_net), .I1(n15513[13]), .I2(n1105), 
            .I3(n52990), .O(n14096[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n52578), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_5 (.CI(n53658), .I0(n14607[2]), .I1(n299_adj_4765), 
            .CO(n53659));
    SB_CARRY add_5037_16 (.CI(n52990), .I0(n15513[13]), .I1(n1105), .CO(n52991));
    SB_CARRY unary_minus_20_add_3_6 (.CI(n52710), .I0(GND_net), .I1(n1_adj_5014[4]), 
            .CO(n52711));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[3]), 
            .I3(n52709), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n52578), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n52579));
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n52577), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_15_lut (.I0(GND_net), .I1(n15513[12]), .I2(n1032), 
            .I3(n52989), .O(n14096[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n52709), .I0(GND_net), .I1(n1_adj_5014[3]), 
            .CO(n52710));
    SB_LUT4 add_4998_4_lut (.I0(GND_net), .I1(n14607[1]), .I2(n226_adj_4767), 
            .I3(n53657), .O(n13100[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[2]), 
            .I3(n52708), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_19 (.CI(n52577), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n52578));
    SB_CARRY add_4998_4 (.CI(n53657), .I0(n14607[1]), .I1(n226_adj_4767), 
            .CO(n53658));
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n52576), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_3_lut (.I0(GND_net), .I1(n14607[0]), .I2(n153_adj_4769), 
            .I3(n53656), .O(n13100[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4998_3 (.CI(n53656), .I0(n14607[0]), .I1(n153_adj_4769), 
            .CO(n53657));
    SB_CARRY add_5037_15 (.CI(n52989), .I0(n15513[12]), .I1(n1032), .CO(n52990));
    SB_LUT4 add_5037_14_lut (.I0(GND_net), .I1(n15513[11]), .I2(n959), 
            .I3(n52988), .O(n14096[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_14 (.CI(n52988), .I0(n15513[11]), .I1(n959), .CO(n52989));
    SB_LUT4 add_5037_13_lut (.I0(GND_net), .I1(n15513[10]), .I2(n886), 
            .I3(n52987), .O(n14096[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4998_2_lut (.I0(GND_net), .I1(n11_adj_4770), .I2(n80_adj_4771), 
            .I3(GND_net), .O(n13100[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4998_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_13 (.CI(n52987), .I0(n15513[10]), .I1(n886), .CO(n52988));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n52708), .I0(GND_net), .I1(n1_adj_5014[2]), 
            .CO(n52709));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[1]), 
            .I3(n52707), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n52576), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n52577));
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n52575), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_12_lut (.I0(GND_net), .I1(n15513[9]), .I2(n813), 
            .I3(n52986), .O(n14096[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_12 (.CI(n52986), .I0(n15513[9]), .I1(n813), .CO(n52987));
    SB_CARRY add_4998_2 (.CI(GND_net), .I0(n11_adj_4770), .I1(n80_adj_4771), 
            .CO(n53656));
    SB_LUT4 add_5060_21_lut (.I0(GND_net), .I1(n15960[18]), .I2(GND_net), 
            .I3(n53655), .O(n14607[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_11_lut (.I0(GND_net), .I1(n15513[8]), .I2(n740), 
            .I3(n52985), .O(n14096[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n52707), .I0(GND_net), .I1(n1_adj_5014[1]), 
            .CO(n52708));
    SB_LUT4 add_5060_20_lut (.I0(GND_net), .I1(n15960[17]), .I2(GND_net), 
            .I3(n53654), .O(n14607[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_11 (.CI(n52985), .I0(n15513[8]), .I1(n740), .CO(n52986));
    SB_CARRY add_5060_20 (.CI(n53654), .I0(n15960[17]), .I1(GND_net), 
            .CO(n53655));
    SB_LUT4 add_5037_10_lut (.I0(GND_net), .I1(n15513[7]), .I2(n667), 
            .I3(n52984), .O(n14096[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_10 (.CI(n52984), .I0(n15513[7]), .I1(n667), .CO(n52985));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5014[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n52575), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n52576));
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n52574), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_16 (.CI(n52574), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n52575));
    SB_LUT4 add_5060_19_lut (.I0(GND_net), .I1(n15960[16]), .I2(GND_net), 
            .I3(n53653), .O(n14607[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_9_lut (.I0(GND_net), .I1(n15513[6]), .I2(n594), .I3(n52983), 
            .O(n14096[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5014[0]), 
            .CO(n52707));
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n52573), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n52573), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n52574));
    SB_CARRY add_5037_9 (.CI(n52983), .I0(n15513[6]), .I1(n594), .CO(n52984));
    SB_LUT4 add_5037_8_lut (.I0(GND_net), .I1(n15513[5]), .I2(n521), .I3(n52982), 
            .O(n14096[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_19 (.CI(n53653), .I0(n15960[16]), .I1(GND_net), 
            .CO(n53654));
    SB_CARRY add_5037_8 (.CI(n52982), .I0(n15513[5]), .I1(n521), .CO(n52983));
    SB_LUT4 add_5037_7_lut (.I0(GND_net), .I1(n15513[4]), .I2(n448_adj_4775), 
            .I3(n52981), .O(n14096[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_18_lut (.I0(GND_net), .I1(n15960[15]), .I2(GND_net), 
            .I3(n53652), .O(n14607[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_7 (.CI(n52981), .I0(n15513[4]), .I1(n448_adj_4775), 
            .CO(n52982));
    SB_LUT4 add_5037_6_lut (.I0(GND_net), .I1(n15513[3]), .I2(n375), .I3(n52980), 
            .O(n14096[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_18 (.CI(n53652), .I0(n15960[15]), .I1(GND_net), 
            .CO(n53653));
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n52572), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n52572), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n52573));
    SB_LUT4 add_5060_17_lut (.I0(GND_net), .I1(n15960[14]), .I2(GND_net), 
            .I3(n53651), .O(n14607[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_6 (.CI(n52980), .I0(n15513[3]), .I1(n375), .CO(n52981));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n52571), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n52571), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n52572));
    SB_LUT4 add_5037_5_lut (.I0(GND_net), .I1(n15513[2]), .I2(n302_adj_4776), 
            .I3(n52979), .O(n14096[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_5 (.CI(n52979), .I0(n15513[2]), .I1(n302_adj_4776), 
            .CO(n52980));
    SB_LUT4 add_5037_4_lut (.I0(GND_net), .I1(n15513[1]), .I2(n229), .I3(n52978), 
            .O(n14096[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_17 (.CI(n53651), .I0(n15960[14]), .I1(GND_net), 
            .CO(n53652));
    SB_CARRY add_5037_4 (.CI(n52978), .I0(n15513[1]), .I1(n229), .CO(n52979));
    SB_LUT4 add_5037_3_lut (.I0(GND_net), .I1(n15513[0]), .I2(n156), .I3(n52977), 
            .O(n14096[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_16_lut (.I0(GND_net), .I1(n15960[13]), .I2(n1105_adj_4777), 
            .I3(n53650), .O(n14607[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_3 (.CI(n52977), .I0(n15513[0]), .I1(n156), .CO(n52978));
    SB_CARRY add_5060_16 (.CI(n53650), .I0(n15960[13]), .I1(n1105_adj_4777), 
            .CO(n53651));
    SB_LUT4 add_5037_2_lut (.I0(GND_net), .I1(n14_adj_4778), .I2(n83), 
            .I3(GND_net), .O(n14096[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_15_lut (.I0(GND_net), .I1(n15960[12]), .I2(n1032_adj_4779), 
            .I3(n53649), .O(n14607[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_15 (.CI(n53649), .I0(n15960[12]), .I1(n1032_adj_4779), 
            .CO(n53650));
    SB_CARRY add_5037_2 (.CI(GND_net), .I0(n14_adj_4778), .I1(n83), .CO(n52977));
    SB_LUT4 add_5097_20_lut (.I0(GND_net), .I1(n16781[17]), .I2(GND_net), 
            .I3(n52976), .O(n15513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_14_lut (.I0(GND_net), .I1(n15960[11]), .I2(n959_adj_4780), 
            .I3(n53648), .O(n14607[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_14 (.CI(n53648), .I0(n15960[11]), .I1(n959_adj_4780), 
            .CO(n53649));
    SB_LUT4 add_5060_13_lut (.I0(GND_net), .I1(n15960[10]), .I2(n886_adj_4781), 
            .I3(n53647), .O(n14607[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_19_lut (.I0(GND_net), .I1(n16781[16]), .I2(GND_net), 
            .I3(n52975), .O(n15513[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_19 (.CI(n52975), .I0(n16781[16]), .I1(GND_net), 
            .CO(n52976));
    SB_CARRY add_5060_13 (.CI(n53647), .I0(n15960[10]), .I1(n886_adj_4781), 
            .CO(n53648));
    SB_LUT4 add_5097_18_lut (.I0(GND_net), .I1(n16781[15]), .I2(GND_net), 
            .I3(n52974), .O(n15513[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_18 (.CI(n52974), .I0(n16781[15]), .I1(GND_net), 
            .CO(n52975));
    SB_LUT4 add_5097_17_lut (.I0(GND_net), .I1(n16781[14]), .I2(GND_net), 
            .I3(n52973), .O(n15513[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_17 (.CI(n52973), .I0(n16781[14]), .I1(GND_net), 
            .CO(n52974));
    SB_LUT4 add_5060_12_lut (.I0(GND_net), .I1(n15960[9]), .I2(n813_adj_4782), 
            .I3(n53646), .O(n14607[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_12 (.CI(n53646), .I0(n15960[9]), .I1(n813_adj_4782), 
            .CO(n53647));
    SB_LUT4 add_5097_16_lut (.I0(GND_net), .I1(n16781[13]), .I2(n1108), 
            .I3(n52972), .O(n15513[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_11_lut (.I0(GND_net), .I1(n15960[8]), .I2(n740_adj_4783), 
            .I3(n53645), .O(n14607[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_16 (.CI(n52972), .I0(n16781[13]), .I1(n1108), .CO(n52973));
    SB_LUT4 add_5097_15_lut (.I0(GND_net), .I1(n16781[12]), .I2(n1035), 
            .I3(n52971), .O(n15513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_11 (.CI(n53645), .I0(n15960[8]), .I1(n740_adj_4783), 
            .CO(n53646));
    SB_CARRY add_5097_15 (.CI(n52971), .I0(n16781[12]), .I1(n1035), .CO(n52972));
    SB_LUT4 add_5097_14_lut (.I0(GND_net), .I1(n16781[11]), .I2(n962), 
            .I3(n52970), .O(n15513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_10_lut (.I0(GND_net), .I1(n15960[7]), .I2(n667_adj_4784), 
            .I3(n53644), .O(n14607[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_10 (.CI(n53644), .I0(n15960[7]), .I1(n667_adj_4784), 
            .CO(n53645));
    SB_CARRY add_5097_14 (.CI(n52970), .I0(n16781[11]), .I1(n962), .CO(n52971));
    SB_LUT4 add_5097_13_lut (.I0(GND_net), .I1(n16781[10]), .I2(n889), 
            .I3(n52969), .O(n15513[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_9_lut (.I0(GND_net), .I1(n15960[6]), .I2(n594_adj_4785), 
            .I3(n53643), .O(n14607[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_9 (.CI(n53643), .I0(n15960[6]), .I1(n594_adj_4785), 
            .CO(n53644));
    SB_LUT4 add_5060_8_lut (.I0(GND_net), .I1(n15960[5]), .I2(n521_adj_4786), 
            .I3(n53642), .O(n14607[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_8 (.CI(n53642), .I0(n15960[5]), .I1(n521_adj_4786), 
            .CO(n53643));
    SB_CARRY add_5097_13 (.CI(n52969), .I0(n16781[10]), .I1(n889), .CO(n52970));
    SB_LUT4 add_5060_7_lut (.I0(GND_net), .I1(n15960[4]), .I2(n448_adj_4787), 
            .I3(n53641), .O(n14607[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_7 (.CI(n53641), .I0(n15960[4]), .I1(n448_adj_4787), 
            .CO(n53642));
    SB_LUT4 add_5060_6_lut (.I0(GND_net), .I1(n15960[3]), .I2(n375_adj_4788), 
            .I3(n53640), .O(n14607[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5060_6 (.CI(n53640), .I0(n15960[3]), .I1(n375_adj_4788), 
            .CO(n53641));
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4534));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5060_5_lut (.I0(GND_net), .I1(n15960[2]), .I2(n302_adj_4789), 
            .I3(n53639), .O(n14607[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_5 (.CI(n53639), .I0(n15960[2]), .I1(n302_adj_4789), 
            .CO(n53640));
    SB_LUT4 add_5060_4_lut (.I0(GND_net), .I1(n15960[1]), .I2(n229_adj_4790), 
            .I3(n53638), .O(n14607[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_12_lut (.I0(GND_net), .I1(n16781[9]), .I2(n816), 
            .I3(n52968), .O(n15513[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_12 (.CI(n52968), .I0(n16781[9]), .I1(n816), .CO(n52969));
    SB_CARRY add_5060_4 (.CI(n53638), .I0(n15960[1]), .I1(n229_adj_4790), 
            .CO(n53639));
    SB_LUT4 add_5060_3_lut (.I0(GND_net), .I1(n15960[0]), .I2(n156_adj_4791), 
            .I3(n53637), .O(n14607[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_11_lut (.I0(GND_net), .I1(n16781[8]), .I2(n743_adj_4792), 
            .I3(n52967), .O(n15513[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_11 (.CI(n52967), .I0(n16781[8]), .I1(n743_adj_4792), 
            .CO(n52968));
    SB_CARRY add_5060_3 (.CI(n53637), .I0(n15960[0]), .I1(n156_adj_4791), 
            .CO(n53638));
    SB_LUT4 add_5060_2_lut (.I0(GND_net), .I1(n14_adj_4793), .I2(n83_adj_4794), 
            .I3(GND_net), .O(n14607[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_2 (.CI(GND_net), .I0(n14_adj_4793), .I1(n83_adj_4794), 
            .CO(n53637));
    SB_LUT4 add_5118_20_lut (.I0(GND_net), .I1(n17167[17]), .I2(GND_net), 
            .I3(n53636), .O(n15960[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_19_lut (.I0(GND_net), .I1(n17167[16]), .I2(GND_net), 
            .I3(n53635), .O(n15960[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5118_19 (.CI(n53635), .I0(n17167[16]), .I1(GND_net), 
            .CO(n53636));
    SB_LUT4 add_5118_18_lut (.I0(GND_net), .I1(n17167[15]), .I2(GND_net), 
            .I3(n53634), .O(n15960[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_18 (.CI(n53634), .I0(n17167[15]), .I1(GND_net), 
            .CO(n53635));
    SB_LUT4 add_5118_17_lut (.I0(GND_net), .I1(n17167[14]), .I2(GND_net), 
            .I3(n53633), .O(n15960[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_17 (.CI(n53633), .I0(n17167[14]), .I1(GND_net), 
            .CO(n53634));
    SB_LUT4 add_5118_16_lut (.I0(GND_net), .I1(n17167[13]), .I2(n1108_adj_4795), 
            .I3(n53632), .O(n15960[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_16 (.CI(n53632), .I0(n17167[13]), .I1(n1108_adj_4795), 
            .CO(n53633));
    SB_LUT4 add_5118_15_lut (.I0(GND_net), .I1(n17167[12]), .I2(n1035_adj_4796), 
            .I3(n53631), .O(n15960[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_15 (.CI(n53631), .I0(n17167[12]), .I1(n1035_adj_4796), 
            .CO(n53632));
    SB_LUT4 add_5118_14_lut (.I0(GND_net), .I1(n17167[11]), .I2(n962_adj_4797), 
            .I3(n53630), .O(n15960[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_14 (.CI(n53630), .I0(n17167[11]), .I1(n962_adj_4797), 
            .CO(n53631));
    SB_LUT4 add_5118_13_lut (.I0(GND_net), .I1(n17167[10]), .I2(n889_adj_4798), 
            .I3(n53629), .O(n15960[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_13 (.CI(n53629), .I0(n17167[10]), .I1(n889_adj_4798), 
            .CO(n53630));
    SB_LUT4 add_5118_12_lut (.I0(GND_net), .I1(n17167[9]), .I2(n816_adj_4799), 
            .I3(n53628), .O(n15960[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_12 (.CI(n53628), .I0(n17167[9]), .I1(n816_adj_4799), 
            .CO(n53629));
    SB_LUT4 add_5118_11_lut (.I0(GND_net), .I1(n17167[8]), .I2(n743), 
            .I3(n53627), .O(n15960[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4800));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4801));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4802));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4803));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n233[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4804));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4805));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4806));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4807));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4808));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4809));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4810));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4811));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4812));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45040_2_lut (.I0(counter[13]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n64295));
    defparam i45040_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48563_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n67833));
    defparam i48563_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i9_4_lut (.I0(counter[5]), .I1(counter[2]), .I2(counter[8]), 
            .I3(counter[3]), .O(n23_adj_4813));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(n233[10]), .I1(n285[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4814));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4815));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4816));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4817));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(counter[1]), .I1(counter[6]), .I2(counter[10]), 
            .I3(counter[0]), .O(n22_adj_4818));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4819));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(n23_adj_4813), .I1(counter[4]), .I2(n64295), 
            .I3(counter[9]), .O(n26_adj_4820));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i51700_4_lut (.I0(counter[12]), .I1(n26_adj_4820), .I2(n22_adj_4818), 
            .I3(counter[7]), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i51700_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48575_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n67845));
    defparam i48575_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48664_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(PWMLimit[9]), 
            .I3(n455[9]), .O(n67934));
    defparam i48664_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48737_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(PWMLimit[7]), 
            .I3(n455[7]), .O(n68007));
    defparam i48737_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n335[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4799));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4798));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4797));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4796));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4795));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4794));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4793));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4792));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4791));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4790));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4789));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4788));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4787));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4786));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4785));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4784));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4783));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4782));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4781));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4780));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4779));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4778));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4777));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4821));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4822));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4776));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4775));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4771));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4769));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4765));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4759));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4757));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4753));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4752));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4751));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4750));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n233[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4748));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4745));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4737));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4729));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5014[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4726));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24049_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41898));   // verilog/motorControl.v(61[20:40])
    defparam i24049_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4723));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4715));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4714));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4712));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4710));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4708));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4706));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4704));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4702));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4701));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4695));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4693));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4689));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4823));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4687));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4686));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4684));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4681));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5013[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4677));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4824));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4676));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4825));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4669));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4665));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4663));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4662));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4661));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4660));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4659));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4655));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4652));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4649));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4647));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4646));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5012[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4645));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24032_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41880));   // verilog/motorControl.v(42[14] 73[8])
    defparam i24032_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n36[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4643));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4642));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49190_4_lut (.I0(n21_adj_4804), .I1(n19_adj_4805), .I2(n17_adj_4806), 
            .I3(n9_adj_4800), .O(n68460));
    defparam i49190_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4641));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4639));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4638));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4637));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4636));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4635));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4634));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49177_4_lut (.I0(n27_adj_4823), .I1(n15_adj_4803), .I2(n13_adj_4802), 
            .I3(n11_adj_4801), .O(n68447));
    defparam i49177_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4632));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48961_2_lut_4_lut (.I0(deadband[21]), .I1(n455[21]), .I2(deadband[9]), 
            .I3(n455[9]), .O(n68231));
    defparam i48961_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4826));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4631));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48994_2_lut_4_lut (.I0(deadband[16]), .I1(n455[16]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n68264));
    defparam i48994_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4629));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i38_2_lut (.I0(\Ki[0] ), .I1(n335[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4628));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49039_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n68309));
    defparam i49039_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4625));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4624));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4623));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4622));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4621));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_970 (.I0(\control_mode[7] ), .I1(\control_mode[6] ), 
            .I2(\control_mode[1] ), .I3(\control_mode[0] ), .O(n27602));
    defparam i1_2_lut_4_lut_adj_970.LUT_INIT = 16'h1000;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4620));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4619));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n23080[2]), .I1(n6_adj_4828), .I2(\Ki[4] ), 
            .I3(n335[18]), .O(n23023[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_9_i32_3_lut_3_lut (.I0(setpoint[15]), .I1(setpoint[16]), 
            .I2(PWMLimit[16]), .I3(GND_net), .O(n32_adj_4829));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i138_2_lut (.I0(\Ki[2] ), .I1(n335[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49334_2_lut_4_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), .I2(PWMLimit[17]), 
            .I3(setpoint[17]), .O(n68604));
    defparam i49334_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i34_3_lut_3_lut (.I0(setpoint[17]), .I1(setpoint[21]), 
            .I2(PWMLimit[21]), .I3(GND_net), .O(n34));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i34_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_971 (.I0(n23138[0]), .I1(n52254), .I2(\Ki[2] ), 
            .I3(n335[20]), .O(n23117[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_971.LUT_INIT = 16'h9666;
    SB_LUT4 mult_24_i89_2_lut (.I0(\Ki[1] ), .I1(n335[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i42_2_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4830));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49491_2_lut_4_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(PWMLimit[5]), 
            .I3(setpoint[5]), .O(n68761));
    defparam i49491_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i10_3_lut_3_lut (.I0(setpoint[5]), .I1(setpoint[6]), 
            .I2(PWMLimit[6]), .I3(GND_net), .O(n10_adj_4831));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(setpoint[2]), .I1(setpoint[3]), 
            .I2(PWMLimit[3]), .I3(GND_net), .O(n6_adj_4832));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49427_2_lut_4_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(PWMLimit[4]), 
            .I3(setpoint[4]), .O(n68697));
    defparam i49427_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i8_3_lut_3_lut (.I0(setpoint[4]), .I1(setpoint[8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_4833));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_4802), 
            .I3(GND_net), .O(n10_adj_4834));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4532));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49073_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n68343));
    defparam i49073_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_4826), .I1(n233[17]), .I2(n35_adj_4824), 
            .I3(GND_net), .O(n30_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34477_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n53911));   // verilog/motorControl.v(61[20:26])
    defparam i34477_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34471_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n52279));   // verilog/motorControl.v(61[20:26])
    defparam i34471_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_972 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n335[22]), 
            .I3(n335[23]), .O(n63933));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_973 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(n335[18]), 
            .I3(n335[19]), .O(n63937));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_973.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4531));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_974 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(n335[20]), 
            .I3(n335[21]), .O(n63935));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_974.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_975 (.I0(n63935), .I1(n52224), .I2(n63937), .I3(n63933), 
            .O(n63943));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i34459_4_lut (.I0(n23138[0]), .I1(\Ki[2] ), .I2(n52254), .I3(n335[20]), 
            .O(n4_adj_4836));   // verilog/motorControl.v(61[29:40])
    defparam i34459_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i34597_4_lut (.I0(n23080[2]), .I1(\Ki[4] ), .I2(n6_adj_4828), 
            .I3(n335[18]), .O(n8_adj_4837));   // verilog/motorControl.v(61[29:40])
    defparam i34597_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_976 (.I0(n6_adj_4838), .I1(n8_adj_4837), .I2(n4_adj_4836), 
            .I3(n63943), .O(n62793));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4617));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4616));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4614));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4613));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4611));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4610));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4608));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4607));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4599));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4598));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4596));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49212_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n68482));
    defparam i49212_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4592));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49251_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n68521));
    defparam i49251_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n335[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50199_4_lut (.I0(n13_adj_4802), .I1(n11_adj_4801), .I2(n9_adj_4800), 
            .I3(n68478), .O(n69469));
    defparam i50199_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50191_4_lut (.I0(n19_adj_4805), .I1(n17_adj_4806), .I2(n15_adj_4803), 
            .I3(n69469), .O(n69461));
    defparam i50191_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51307_4_lut (.I0(n25_adj_4808), .I1(n23_adj_4807), .I2(n21_adj_4804), 
            .I3(n69461), .O(n70577));
    defparam i51307_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50714_4_lut (.I0(n31_c), .I1(n29_adj_4825), .I2(n27_adj_4823), 
            .I3(n70577), .O(n69984));
    defparam i50714_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51446_4_lut (.I0(n37), .I1(n35_adj_4824), .I2(n33), .I3(n69984), 
            .O(n70716));
    defparam i51446_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4529));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4839));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i75_2_lut (.I0(\Ki[1] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4587));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4586));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4457));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4456));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4584));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4583));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51004_3_lut (.I0(n6_adj_4840), .I1(n233[10]), .I2(n21_adj_4804), 
            .I3(GND_net), .O(n70274));   // verilog/motorControl.v(56[14:36])
    defparam i51004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51005_3_lut (.I0(n70274), .I1(n233[11]), .I2(n23_adj_4807), 
            .I3(GND_net), .O(n70275));   // verilog/motorControl.v(56[14:36])
    defparam i51005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_4806), 
            .I3(GND_net), .O(n8_adj_4841));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4839), .I1(n233[22]), .I2(n45_adj_4821), 
            .I3(GND_net), .O(n24_adj_4842));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49147_4_lut (.I0(n43), .I1(n25_adj_4808), .I2(n23_adj_4807), 
            .I3(n68460), .O(n68417));
    defparam i49147_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4582));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50512_4_lut (.I0(n24_adj_4842), .I1(n8_adj_4841), .I2(n45_adj_4821), 
            .I3(n68411), .O(n69782));   // verilog/motorControl.v(56[14:36])
    defparam i50512_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49694_3_lut (.I0(n70275), .I1(n233[12]), .I2(n25_adj_4808), 
            .I3(GND_net), .O(n68964));   // verilog/motorControl.v(56[14:36])
    defparam i49694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49141_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n68411));
    defparam i49141_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i34493_2_lut_4_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(\Ki[1] ), 
            .I3(n335[19]), .O(n23080[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34493_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i49165_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n68435));
    defparam i49165_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4843));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i51000_3_lut (.I0(n4_adj_4843), .I1(n233[13]), .I2(n27_adj_4823), 
            .I3(GND_net), .O(n70270));   // verilog/motorControl.v(56[14:36])
    defparam i51000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51001_3_lut (.I0(n70270), .I1(n233[14]), .I2(n29_adj_4825), 
            .I3(GND_net), .O(n70271));   // verilog/motorControl.v(56[14:36])
    defparam i51001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49171_4_lut (.I0(n33), .I1(n31_c), .I2(n29_adj_4825), .I3(n68447), 
            .O(n68441));
    defparam i49171_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n335[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n335[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n310[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i22_3_lut (.I0(n310[21]), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n335[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n335[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n335[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i19_3_lut (.I0(n233[18]), .I1(n285[18]), .I2(n284), 
            .I3(GND_net), .O(n310[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i19_3_lut (.I0(n310[18]), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n335[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n335[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n335[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n335[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n335[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23604_3_lut (.I0(\control_mode[0] ), .I1(control_update), .I2(n27629), 
            .I3(GND_net), .O(n29776));
    defparam i23604_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n335[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4455));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4453));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n335[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4452));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51323_4_lut (.I0(n30_c), .I1(n10_adj_4834), .I2(n35_adj_4824), 
            .I3(n68435), .O(n70593));   // verilog/motorControl.v(56[14:36])
    defparam i51323_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4528));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4451));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49696_3_lut (.I0(n70271), .I1(n233[15]), .I2(n31_c), .I3(GND_net), 
            .O(n68966));   // verilog/motorControl.v(56[14:36])
    defparam i49696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51535_4_lut (.I0(n68966), .I1(n70593), .I2(n35_adj_4824), 
            .I3(n68441), .O(n70805));   // verilog/motorControl.v(56[14:36])
    defparam i51535_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4450));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4449));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4581));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51536_3_lut (.I0(n70805), .I1(n233[18]), .I2(n37), .I3(GND_net), 
            .O(n70806));   // verilog/motorControl.v(56[14:36])
    defparam i51536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51522_3_lut (.I0(n70806), .I1(n233[19]), .I2(n39), .I3(GND_net), 
            .O(n70792));   // verilog/motorControl.v(56[14:36])
    defparam i51522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49151_4_lut (.I0(n43), .I1(n41_adj_4822), .I2(n39), .I3(n70716), 
            .O(n68421));
    defparam i49151_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51167_4_lut (.I0(n68964), .I1(n69782), .I2(n45_adj_4821), 
            .I3(n68417), .O(n70437));   // verilog/motorControl.v(56[14:36])
    defparam i51167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51682_3_lut_4_lut (.I0(n54181), .I1(\control_mode[0] ), .I2(n27629), 
            .I3(\displacement[0] ), .O(motor_state[0]));   // verilog/motorControl.v(53[17:33])
    defparam i51682_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i49702_3_lut (.I0(n70792), .I1(n233[20]), .I2(n41_adj_4822), 
            .I3(GND_net), .O(n68972));   // verilog/motorControl.v(56[14:36])
    defparam i49702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71308_bdd_4_lut (.I0(n71308), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4751), .O(n71311));
    defparam n71308_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4849));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4850));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4851));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4852));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4853));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4854));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4855));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4579));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4578));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4856));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4577));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4857));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4576));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4575));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4858));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24004_2_lut_4_lut (.I0(control_update), .I1(n27602), .I2(n59660), 
            .I3(n41540), .O(n41850));
    defparam i24004_2_lut_4_lut.LUT_INIT = 16'hff5d;
    SB_LUT4 i1_2_lut_4_lut_adj_977 (.I0(control_update), .I1(n27602), .I2(n59660), 
            .I3(n41540), .O(n27506));
    defparam i1_2_lut_4_lut_adj_977.LUT_INIT = 16'h5dff;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4859));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4860));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49037_3_lut_4_lut (.I0(deadband[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(deadband[2]), .O(n68307));   // verilog/motorControl.v(62[14:31])
    defparam i49037_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4861));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48559_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n67557));
    defparam i48559_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4862));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48781_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n67558));
    defparam i48781_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48780_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n67559));
    defparam i48780_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n310[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i13_3_lut (.I0(n310[12]), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n335[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i26_2_lut (.I0(\Ki[0] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48658_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n67563));
    defparam i48658_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4863));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48778_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n67564));
    defparam i48778_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48777_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n67565));
    defparam i48777_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48776_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n67566));
    defparam i48776_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48775_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n67567));
    defparam i48775_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4864));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48706_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[15]), 
            .I3(GND_net), .O(n67568));
    defparam i48706_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4865));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4866));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4867));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48783_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n67801));
    defparam i48783_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4868));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51411_4_lut (.I0(n68972), .I1(n70437), .I2(n45_adj_4821), 
            .I3(n68421), .O(n70681));   // verilog/motorControl.v(56[14:36])
    defparam i51411_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49303_4_lut (.I0(n21_adj_4866), .I1(n19_adj_4865), .I2(n17_adj_4864), 
            .I3(n9_adj_4863), .O(n68573));
    defparam i49303_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51412_3_lut (.I0(n70681), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i51412_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49278_4_lut (.I0(n27_adj_4862), .I1(n15_adj_4867), .I2(n13_adj_4860), 
            .I3(n11_adj_4859), .O(n68548));
    defparam i49278_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4868), 
            .I3(GND_net), .O(n12_adj_4869));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48784_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[4]), 
            .I3(GND_net), .O(n67800));
    defparam i48784_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4574));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4860), 
            .I3(GND_net), .O(n10_adj_4870));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48785_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n67799));
    defparam i48785_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48786_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n67798));
    defparam i48786_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48635_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n67797));
    defparam i48635_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i49508_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[0]), 
            .I3(GND_net), .O(n67796));
    defparam i49508_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4869), .I1(n535[17]), .I2(n35_adj_4858), 
            .I3(GND_net), .O(n30_adj_4871));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48920_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[23]), 
            .I3(GND_net), .O(n67744));
    defparam i48920_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48699_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n67600));
    defparam i48699_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48684_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n67593));
    defparam i48684_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48643_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[20]), 
            .I3(GND_net), .O(n67587));
    defparam i48643_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48956_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n67584));
    defparam i48956_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48987_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n67569));
    defparam i48987_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48774_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n67570));
    defparam i48774_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48662_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n67575));
    defparam i48662_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i49524_2_lut_3_lut (.I0(n7073), .I1(n27508), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n67803));
    defparam i49524_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48656_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n67926));   // verilog/motorControl.v(65[25:41])
    defparam i48656_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50299_4_lut (.I0(n13_adj_4860), .I1(n11_adj_4859), .I2(n9_adj_4863), 
            .I3(n68596), .O(n69569));
    defparam i50299_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4872));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50285_4_lut (.I0(n19_adj_4865), .I1(n17_adj_4864), .I2(n15_adj_4867), 
            .I3(n69569), .O(n69555));
    defparam i50285_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51349_4_lut (.I0(n25_adj_4857), .I1(n23_adj_4856), .I2(n21_adj_4866), 
            .I3(n69555), .O(n70619));
    defparam i51349_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50754_4_lut (.I0(n31_adj_4854), .I1(n29_adj_4853), .I2(n27_adj_4862), 
            .I3(n70619), .O(n70024));
    defparam i50754_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n335[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4573));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4572));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34655_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4874), 
            .I3(GND_net), .O(n23044[0]));   // verilog/motorControl.v(61[20:26])
    defparam i34655_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4874), 
            .I3(n63987), .O(n23044[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i51464_4_lut (.I0(n37_adj_4855), .I1(n35_adj_4858), .I2(n33_adj_4868), 
            .I3(n70024), .O(n70734));
    defparam i51464_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4852), 
            .I3(GND_net), .O(n16_adj_4875));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51014_3_lut (.I0(n6_adj_4876), .I1(n535[10]), .I2(n21_adj_4866), 
            .I3(GND_net), .O(n70284));   // verilog/motorControl.v(47[25:43])
    defparam i51014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51015_3_lut (.I0(n70284), .I1(n535[11]), .I2(n23_adj_4856), 
            .I3(GND_net), .O(n70285));   // verilog/motorControl.v(47[25:43])
    defparam i51015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4571));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_978 (.I0(n70679), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n27538), .O(n7071));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut_adj_978.LUT_INIT = 16'h7100;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4864), 
            .I3(GND_net), .O(n8_adj_4877));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4570));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4875), .I1(n535[22]), .I2(n45_adj_4851), 
            .I3(GND_net), .O(n24_adj_4878));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49214_4_lut (.I0(n43_adj_4852), .I1(n25_adj_4857), .I2(n23_adj_4856), 
            .I3(n68573), .O(n68484));
    defparam i49214_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50510_4_lut (.I0(n24_adj_4878), .I1(n8_adj_4877), .I2(n45_adj_4851), 
            .I3(n68482), .O(n69780));   // verilog/motorControl.v(47[25:43])
    defparam i50510_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_adj_979 (.I0(n70679), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n27538), .O(n27540));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut_adj_979.LUT_INIT = 16'h8e00;
    SB_LUT4 i49684_3_lut (.I0(n70285), .I1(n535[12]), .I2(n25_adj_4857), 
            .I3(GND_net), .O(n68954));   // verilog/motorControl.v(47[25:43])
    defparam i49684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4569));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4879));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51010_3_lut (.I0(n4_adj_4879), .I1(n535[13]), .I2(n27_adj_4862), 
            .I3(GND_net), .O(n70280));   // verilog/motorControl.v(47[25:43])
    defparam i51010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51011_3_lut (.I0(n70280), .I1(n535[14]), .I2(n29_adj_4853), 
            .I3(GND_net), .O(n70281));   // verilog/motorControl.v(47[25:43])
    defparam i51011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49257_4_lut (.I0(n33_adj_4868), .I1(n31_adj_4854), .I2(n29_adj_4853), 
            .I3(n68548), .O(n68527));
    defparam i49257_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51321_4_lut (.I0(n30_adj_4871), .I1(n10_adj_4870), .I2(n35_adj_4858), 
            .I3(n68521), .O(n70591));   // verilog/motorControl.v(47[25:43])
    defparam i51321_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4567));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4880));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9980_bdd_4_lut_52015 (.I0(n9980), .I1(n67593), .I2(setpoint[21]), 
            .I3(n4751), .O(n71290));
    defparam n9980_bdd_4_lut_52015.LUT_INIT = 16'he4aa;
    SB_LUT4 i49686_3_lut (.I0(n70281), .I1(n535[15]), .I2(n31_adj_4854), 
            .I3(GND_net), .O(n68956));   // verilog/motorControl.v(47[25:43])
    defparam i49686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4566));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4565));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51533_4_lut (.I0(n68956), .I1(n70591), .I2(n35_adj_4858), 
            .I3(n68527), .O(n70803));   // verilog/motorControl.v(47[25:43])
    defparam i51533_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n335[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4564));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4563));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n335[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4562));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4561));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4882));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51534_3_lut (.I0(n70803), .I1(n535[18]), .I2(n37_adj_4855), 
            .I3(GND_net), .O(n70804));   // verilog/motorControl.v(47[25:43])
    defparam i51534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4559));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4558));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4557));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51524_3_lut (.I0(n70804), .I1(n535[19]), .I2(n39_adj_4849), 
            .I3(GND_net), .O(n70794));   // verilog/motorControl.v(47[25:43])
    defparam i51524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49217_4_lut (.I0(n43_adj_4852), .I1(n41_adj_4850), .I2(n39_adj_4849), 
            .I3(n70734), .O(n68487));
    defparam i49217_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51165_4_lut (.I0(n68954), .I1(n69780), .I2(n45_adj_4851), 
            .I3(n68484), .O(n70435));   // verilog/motorControl.v(47[25:43])
    defparam i51165_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49692_3_lut (.I0(n70794), .I1(n535[20]), .I2(n41_adj_4850), 
            .I3(GND_net), .O(n68962));   // verilog/motorControl.v(47[25:43])
    defparam i49692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51409_4_lut (.I0(n68962), .I1(n70435), .I2(n45_adj_4851), 
            .I3(n68487), .O(n70679));   // verilog/motorControl.v(47[25:43])
    defparam i51409_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n71290_bdd_4_lut (.I0(n71290), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4751), .O(n71293));
    defparam n71290_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4883));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4884));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4885));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4556));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4555));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49326_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n68596));   // verilog/motorControl.v(47[25:43])
    defparam i49326_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4554));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4553));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(n233[18]), .I1(n285[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4886));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n455[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4887));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4552));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4888));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4550));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4549));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4548));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_c));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4547));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4889));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n335[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4891));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_4876));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4546));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4892));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4893));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4894));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4895));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4896));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4897));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4898));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n455[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4899));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_980 (.I0(n207[23]), .I1(\Kp[2] ), .I2(n52284), 
            .I3(n207[22]), .O(n63987));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_980.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n455[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4900));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4901));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4902));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9980_bdd_4_lut_52001 (.I0(n9980), .I1(n67587), .I2(setpoint[20]), 
            .I3(n4751), .O(n71284));
    defparam n9980_bdd_4_lut_52001.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4903));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_981 (.I0(n207[22]), .I1(n23092[1]), .I2(n4_adj_4904), 
            .I3(\Kp[3] ), .O(n23044[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hc66c;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4905));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_4906));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_982 (.I0(n23092[1]), .I1(n6_adj_4907), .I2(n347_adj_4906), 
            .I3(n60085), .O(n23044[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4908));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4909));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(n63983), .I1(n207[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4904));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34676_4_lut (.I0(n23092[1]), .I1(\Kp[3] ), .I2(n4_adj_4904), 
            .I3(n207[22]), .O(n6_adj_4907));   // verilog/motorControl.v(61[20:26])
    defparam i34676_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i49105_4_lut (.I0(n21_adj_4814), .I1(n19_adj_4815), .I2(n17_adj_4816), 
            .I3(n9_adj_4809), .O(n68375));
    defparam i49105_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n63983));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i45130_3_lut (.I0(n207[23]), .I1(n63983), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n60085));   // verilog/motorControl.v(61[20:26])
    defparam i45130_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i34616_3_lut (.I0(n207[23]), .I1(n52279), .I2(n53911), .I3(GND_net), 
            .O(n23092[1]));   // verilog/motorControl.v(61[20:26])
    defparam i34616_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_23_i46_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_4874));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34607_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n52284));   // verilog/motorControl.v(61[20:26])
    defparam i34607_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_983 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n53911), 
            .I3(n207[22]), .O(n63973));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_983.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_450_2_lut (.I0(n23092[1]), .I1(n60085), .I2(GND_net), 
            .I3(GND_net), .O(n72161));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_450_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_984 (.I0(n52279), .I1(n63973), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n63977));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_984.LUT_INIT = 16'h9666;
    SB_LUT4 i34684_4_lut (.I0(n72161), .I1(\Kp[4] ), .I2(n6_adj_4907), 
            .I3(n207[22]), .O(n8_adj_4910));   // verilog/motorControl.v(61[20:26])
    defparam i34684_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i34630_4_lut (.I0(n23092[1]), .I1(\Kp[3] ), .I2(n63983), .I3(n207[23]), 
            .O(n6_adj_4911));   // verilog/motorControl.v(61[20:26])
    defparam i34630_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_985 (.I0(n6_adj_4911), .I1(n8_adj_4910), .I2(n63977), 
            .I3(n60085), .O(n61693));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4912));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4913));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4544));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i41_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4914));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4543));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49089_4_lut (.I0(n27), .I1(n15_adj_4812), .I2(n13_adj_4811), 
            .I3(n11_adj_4810), .O(n68359));
    defparam i49089_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4541));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4540));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4915));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i15_2_lut (.I0(PWMLimit[7]), .I1(setpoint[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4916));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i13_2_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4917));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i19_2_lut (.I0(PWMLimit[9]), .I1(setpoint[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4918));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n71284_bdd_4_lut (.I0(n71284), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4751), .O(n71287));
    defparam n71284_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_4893), 
            .I3(GND_net), .O(n12_adj_4919));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i17_2_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4920));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i7_2_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4921));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i9_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4922));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i11_2_lut (.I0(PWMLimit[5]), .I1(setpoint[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4923));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i5_2_lut (.I0(PWMLimit[2]), .I1(setpoint[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4924));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49493_4_lut (.I0(n11_adj_4923), .I1(n9_adj_4922), .I2(n7_adj_4921), 
            .I3(n5_adj_4924), .O(n68763));
    defparam i49493_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9980_bdd_4_lut_51996 (.I0(n9980), .I1(n67584), .I2(setpoint[19]), 
            .I3(n4751), .O(n71278));
    defparam n9980_bdd_4_lut_51996.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_9_i16_3_lut (.I0(n8_adj_4833), .I1(setpoint[9]), .I2(n19_adj_4918), 
            .I3(GND_net), .O(n16_adj_4925));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_4926));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_9_i12_3_lut (.I0(n10_adj_4831), .I1(setpoint[7]), .I2(n15_adj_4916), 
            .I3(GND_net), .O(n12_adj_4927));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49485_4_lut (.I0(n17_adj_4920), .I1(n15_adj_4916), .I2(n13_adj_4917), 
            .I3(n68763), .O(n68755));
    defparam i49485_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51319_4_lut (.I0(n16_adj_4925), .I1(n6_adj_4832), .I2(n19_adj_4918), 
            .I3(n68697), .O(n70589));   // verilog/motorControl.v(45[16:33])
    defparam i51319_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50508_4_lut (.I0(n12_adj_4927), .I1(n4_adj_4926), .I2(n15_adj_4916), 
            .I3(n68761), .O(n69778));   // verilog/motorControl.v(45[16:33])
    defparam i50508_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51574_4_lut (.I0(n69778), .I1(n70589), .I2(n19_adj_4918), 
            .I3(n68755), .O(n70844));   // verilog/motorControl.v(45[16:33])
    defparam i51574_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51575_3_lut (.I0(n70844), .I1(setpoint[10]), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n70845));   // verilog/motorControl.v(45[16:33])
    defparam i51575_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51469_3_lut (.I0(n70845), .I1(setpoint[11]), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n70739));   // verilog/motorControl.v(45[16:33])
    defparam i51469_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50855_3_lut (.I0(n70739), .I1(setpoint[12]), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n70125));   // verilog/motorControl.v(45[16:33])
    defparam i50855_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50856_3_lut (.I0(n70125), .I1(setpoint[13]), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n28));   // verilog/motorControl.v(45[16:33])
    defparam i50856_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4811), 
            .I3(GND_net), .O(n10_adj_4928));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71278_bdd_4_lut (.I0(n71278), .I1(n535[19]), .I2(n455[19]), 
            .I3(n4751), .O(n71281));
    defparam n71278_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_9_i33_2_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4929));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4919), .I1(n285[17]), .I2(n35_adj_4905), 
            .I3(GND_net), .O(n30_adj_4930));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i35_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4931));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i37_2_lut (.I0(PWMLimit[18]), .I1(setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4932));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i43_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4933));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49353_4_lut (.I0(n37_adj_4932), .I1(n35_adj_4931), .I2(n33_adj_4929), 
            .I3(n31), .O(n68623));
    defparam i49353_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_9_i42_3_lut (.I0(n34), .I1(setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n42));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51016_3_lut (.I0(n30), .I1(setpoint[18]), .I2(n37_adj_4932), 
            .I3(GND_net), .O(n70286));   // verilog/motorControl.v(45[16:33])
    defparam i51016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51017_3_lut (.I0(n70286), .I1(setpoint[19]), .I2(n39_adj_4915), 
            .I3(GND_net), .O(n70287));   // verilog/motorControl.v(45[16:33])
    defparam i51017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49338_4_lut (.I0(n43_adj_4933), .I1(n41_adj_4914), .I2(n39_adj_4915), 
            .I3(n68623), .O(n68608));
    defparam i49338_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50857_4_lut (.I0(n42), .I1(n32_adj_4829), .I2(n45), .I3(n68604), 
            .O(n70127));   // verilog/motorControl.v(45[16:33])
    defparam i50857_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49682_3_lut (.I0(n70287), .I1(setpoint[20]), .I2(n41_adj_4914), 
            .I3(GND_net), .O(n68952));   // verilog/motorControl.v(45[16:33])
    defparam i49682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51407_4_lut (.I0(n68952), .I1(n70127), .I2(n45), .I3(n68608), 
            .O(n70677));   // verilog/motorControl.v(45[16:33])
    defparam i51407_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51408_3_lut (.I0(n70677), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i51408_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4937));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i39_2_lut (.I0(deadband[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4938));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i45_2_lut (.I0(deadband[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4939));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(deadband[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4940));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(deadband[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4941));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i43_2_lut (.I0(deadband[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4942));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i37_2_lut (.I0(deadband[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4943));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4944));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4945));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4946));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9980_bdd_4_lut_51991 (.I0(n9980), .I1(n67575), .I2(setpoint[18]), 
            .I3(n4751), .O(n71272));
    defparam n9980_bdd_4_lut_51991.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4947));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(deadband[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4948));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(deadband[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4949));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(deadband[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4950));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50133_4_lut (.I0(n13_adj_4811), .I1(n11_adj_4810), .I2(n9_adj_4809), 
            .I3(n68409), .O(n69403));
    defparam i50133_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_26_i33_2_lut (.I0(deadband[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4951));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(deadband[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4952));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4953));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4954));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(deadband[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4955));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50117_4_lut (.I0(n19_adj_4815), .I1(n17_adj_4816), .I2(n15_adj_4812), 
            .I3(n69403), .O(n69387));
    defparam i50117_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48950_4_lut (.I0(n455[6]), .I1(n455[5]), .I2(n46[6]), .I3(n46[5]), 
            .O(n68220));
    defparam i48950_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i49973_3_lut (.I0(n455[7]), .I1(n68220), .I2(n46[7]), .I3(GND_net), 
            .O(n69243));
    defparam i49973_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_28_i27_rep_116_2_lut (.I0(n455[13]), .I1(n46[13]), 
            .I2(GND_net), .I3(GND_net), .O(n71827));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_rep_116_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49939_4_lut (.I0(n455[14]), .I1(n71827), .I2(n46[14]), .I3(n69243), 
            .O(n69209));
    defparam i49939_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i31_rep_111_2_lut (.I0(n455[15]), .I1(n46[15]), 
            .I2(GND_net), .I3(GND_net), .O(n71822));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_rep_111_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48939_4_lut (.I0(n455[8]), .I1(n455[4]), .I2(n46[8]), .I3(n46[4]), 
            .O(n68209));
    defparam i48939_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i49965_3_lut (.I0(n455[9]), .I1(n68209), .I2(n46[9]), .I3(GND_net), 
            .O(n69235));
    defparam i49965_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_28_i21_rep_131_2_lut (.I0(n455[10]), .I1(n46[10]), 
            .I2(GND_net), .I3(GND_net), .O(n71842));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_rep_131_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49959_4_lut (.I0(n455[11]), .I1(n71842), .I2(n46[11]), .I3(n69235), 
            .O(n69229));
    defparam i49959_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i25_rep_126_2_lut (.I0(n455[12]), .I1(n46[12]), 
            .I2(GND_net), .I3(GND_net), .O(n71837));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_rep_126_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51293_4_lut (.I0(n25_adj_4819), .I1(n23_adj_4817), .I2(n21_adj_4814), 
            .I3(n69387), .O(n70563));
    defparam i51293_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n46[9]), .I1(n46[21]), .I2(n455[21]), 
            .I3(GND_net), .O(n16_adj_4956));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48850_4_lut (.I0(n455[21]), .I1(n455[9]), .I2(n46[21]), .I3(n46[9]), 
            .O(n68120));
    defparam i48850_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n46[4]), .I1(n46[8]), .I2(n455[8]), 
            .I3(GND_net), .O(n8_adj_4957));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i24_3_lut (.I0(n16_adj_4956), .I1(n46[22]), .I2(n455[22]), 
            .I3(GND_net), .O(n24_adj_4958));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50678_4_lut (.I0(n31_adj_4889), .I1(n29_adj_4901), .I2(n27), 
            .I3(n70563), .O(n69948));
    defparam i50678_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48959_4_lut (.I0(n455[3]), .I1(n455[2]), .I2(n46[3]), .I3(n46[2]), 
            .O(n68229));
    defparam i48959_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i9_rep_124_2_lut (.I0(n455[4]), .I1(n46[4]), .I2(GND_net), 
            .I3(GND_net), .O(n71835));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_rep_124_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48952_4_lut (.I0(n455[5]), .I1(n71835), .I2(n46[5]), .I3(n68229), 
            .O(n68222));
    defparam i48952_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i13_rep_152_2_lut (.I0(n455[6]), .I1(n46[6]), .I2(GND_net), 
            .I3(GND_net), .O(n71863));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_rep_152_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50618_4_lut (.I0(n455[7]), .I1(n71863), .I2(n46[7]), .I3(n68222), 
            .O(n69888));
    defparam i50618_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i17_rep_149_2_lut (.I0(n455[8]), .I1(n46[8]), .I2(GND_net), 
            .I3(GND_net), .O(n71860));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_rep_149_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51442_4_lut (.I0(n37_adj_4886), .I1(n35_adj_4905), .I2(n33_adj_4893), 
            .I3(n69948), .O(n70712));
    defparam i51442_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_4884), 
            .I3(GND_net), .O(n16_adj_4959));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49969_4_lut (.I0(n455[9]), .I1(n71860), .I2(n46[9]), .I3(n69888), 
            .O(n69239));
    defparam i49969_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i50996_3_lut (.I0(n6_adj_4960), .I1(n285[10]), .I2(n21_adj_4814), 
            .I3(GND_net), .O(n70266));   // verilog/motorControl.v(58[23:46])
    defparam i50996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71272_bdd_4_lut (.I0(n71272), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4751), .O(n71275));
    defparam n71272_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50984_4_lut (.I0(n455[11]), .I1(n71842), .I2(n46[11]), .I3(n69239), 
            .O(n70254));
    defparam i50984_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i50997_3_lut (.I0(n70266), .I1(n285[11]), .I2(n23_adj_4817), 
            .I3(GND_net), .O(n70267));   // verilog/motorControl.v(58[23:46])
    defparam i50997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48924_4_lut (.I0(n455[13]), .I1(n71837), .I2(n46[13]), .I3(n70254), 
            .O(n68194));
    defparam i48924_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_4816), 
            .I3(GND_net), .O(n8_adj_4961));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4959), .I1(n285[22]), .I2(n45_adj_4880), 
            .I3(GND_net), .O(n24_adj_4962));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i29_rep_114_2_lut (.I0(n455[14]), .I1(n46[14]), 
            .I2(GND_net), .I3(GND_net), .O(n71825));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_rep_114_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49045_4_lut (.I0(n43_adj_4884), .I1(n25_adj_4819), .I2(n23_adj_4817), 
            .I3(n68375), .O(n68315));
    defparam i49045_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50592_4_lut (.I0(n455[15]), .I1(n71825), .I2(n46[15]), .I3(n68194), 
            .O(n69862));
    defparam i50592_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i33_rep_143_2_lut (.I0(n455[16]), .I1(n46[16]), 
            .I2(GND_net), .I3(GND_net), .O(n71854));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_rep_143_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51239_4_lut (.I0(n455[17]), .I1(n71854), .I2(n46[17]), .I3(n69862), 
            .O(n70509));
    defparam i51239_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i37_rep_105_2_lut (.I0(n455[18]), .I1(n46[18]), 
            .I2(GND_net), .I3(GND_net), .O(n71816));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i37_rep_105_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50514_4_lut (.I0(n24_adj_4962), .I1(n8_adj_4961), .I2(n45_adj_4880), 
            .I3(n68309), .O(n69784));   // verilog/motorControl.v(58[23:46])
    defparam i50514_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49704_3_lut (.I0(n70267), .I1(n285[12]), .I2(n25_adj_4819), 
            .I3(GND_net), .O(n68974));   // verilog/motorControl.v(58[23:46])
    defparam i49704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51500_4_lut (.I0(n455[19]), .I1(n71816), .I2(n46[19]), .I3(n70509), 
            .O(n70770));
    defparam i51500_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_4963));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_28_i41_rep_102_2_lut (.I0(n455[20]), .I1(n46[20]), 
            .I2(GND_net), .I3(GND_net), .O(n71813));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i41_rep_102_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49008_4_lut (.I0(n27_adj_4955), .I1(n15_adj_4954), .I2(n13_adj_4953), 
            .I3(n11_adj_4952), .O(n68278));
    defparam i49008_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4951), 
            .I3(GND_net), .O(n12_adj_4964));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4953), 
            .I3(GND_net), .O(n10_adj_4965));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50994_3_lut (.I0(n4_adj_4963), .I1(n285[13]), .I2(n27), .I3(GND_net), 
            .O(n70264));   // verilog/motorControl.v(58[23:46])
    defparam i50994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i30_3_lut (.I0(n12_adj_4964), .I1(n455[17]), .I2(n35_adj_4950), 
            .I3(GND_net), .O(n30_adj_4966));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50995_3_lut (.I0(n70264), .I1(n285[14]), .I2(n29_adj_4901), 
            .I3(GND_net), .O(n70265));   // verilog/motorControl.v(58[23:46])
    defparam i50995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50041_4_lut (.I0(n13_adj_4953), .I1(n11_adj_4952), .I2(n9_adj_4949), 
            .I3(n68307), .O(n69311));
    defparam i50041_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50033_4_lut (.I0(n19_adj_4945), .I1(n17_adj_4944), .I2(n15_adj_4954), 
            .I3(n69311), .O(n69303));
    defparam i50033_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51283_4_lut (.I0(n25_adj_4948), .I1(n23_adj_4947), .I2(n21_adj_4946), 
            .I3(n69303), .O(n70553));
    defparam i51283_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50642_4_lut (.I0(n31_adj_4941), .I1(n29_adj_4940), .I2(n27_adj_4955), 
            .I3(n70553), .O(n69912));
    defparam i50642_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51438_4_lut (.I0(n37_adj_4943), .I1(n35_adj_4950), .I2(n33_adj_4951), 
            .I3(n69912), .O(n70708));
    defparam i51438_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4942), 
            .I3(GND_net), .O(n16_adj_4967));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9980_bdd_4_lut_51986 (.I0(n9980), .I1(n67570), .I2(setpoint[17]), 
            .I3(n4751), .O(n71266));
    defparam n9980_bdd_4_lut_51986.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4944), 
            .I3(GND_net), .O(n8_adj_4968));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i24_3_lut (.I0(n16_adj_4967), .I1(n455[22]), .I2(n45_adj_4939), 
            .I3(GND_net), .O(n24_adj_4969));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49081_4_lut (.I0(n33_adj_4893), .I1(n31_adj_4889), .I2(n29_adj_4901), 
            .I3(n68359), .O(n68351));
    defparam i49081_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50990_3_lut (.I0(n6_adj_4861), .I1(n455[10]), .I2(n21_adj_4946), 
            .I3(GND_net), .O(n70260));   // verilog/motorControl.v(62[14:31])
    defparam i50990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50991_3_lut (.I0(n70260), .I1(n455[11]), .I2(n23_adj_4947), 
            .I3(GND_net), .O(n70261));   // verilog/motorControl.v(62[14:31])
    defparam i50991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49016_4_lut (.I0(n21_adj_4946), .I1(n19_adj_4945), .I2(n17_adj_4944), 
            .I3(n9_adj_4949), .O(n68286));
    defparam i49016_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48966_4_lut (.I0(n43_adj_4942), .I1(n25_adj_4948), .I2(n23_adj_4947), 
            .I3(n68286), .O(n68236));
    defparam i48966_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50516_4_lut (.I0(n24_adj_4969), .I1(n8_adj_4968), .I2(n45_adj_4939), 
            .I3(n68231), .O(n69786));   // verilog/motorControl.v(62[14:31])
    defparam i50516_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51325_4_lut (.I0(n30_adj_4930), .I1(n10_adj_4928), .I2(n35_adj_4905), 
            .I3(n68343), .O(n70595));   // verilog/motorControl.v(58[23:46])
    defparam i51325_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49706_3_lut (.I0(n70265), .I1(n285[15]), .I2(n31_adj_4889), 
            .I3(GND_net), .O(n68976));   // verilog/motorControl.v(58[23:46])
    defparam i49706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49714_3_lut (.I0(n70261), .I1(n455[12]), .I2(n25_adj_4948), 
            .I3(GND_net), .O(n68984));   // verilog/motorControl.v(62[14:31])
    defparam i49714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n67612), .I1(n46[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_4970));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50604_3_lut (.I0(n4_adj_4970), .I1(n46[13]), .I2(n455[13]), 
            .I3(GND_net), .O(n69874));   // verilog/motorControl.v(62[35:55])
    defparam i50604_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51539_4_lut (.I0(n68976), .I1(n70595), .I2(n35_adj_4905), 
            .I3(n68351), .O(n70809));   // verilog/motorControl.v(58[23:46])
    defparam i51539_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50605_3_lut (.I0(n69874), .I1(n46[14]), .I2(n455[14]), .I3(GND_net), 
            .O(n69875));   // verilog/motorControl.v(62[35:55])
    defparam i50605_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n46[7]), .I1(n46[16]), .I2(n455[16]), 
            .I3(GND_net), .O(n12_adj_4971));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48881_4_lut (.I0(n455[16]), .I1(n455[7]), .I2(n46[16]), .I3(n46[7]), 
            .O(n68151));
    defparam i48881_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i35_rep_137_2_lut (.I0(n455[17]), .I1(n46[17]), 
            .I2(GND_net), .I3(GND_net), .O(n71848));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_rep_137_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n46[5]), .I1(n46[6]), .I2(n455[6]), 
            .I3(GND_net), .O(n10_adj_4972));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_4971), .I1(n46[17]), .I2(n455[17]), 
            .I3(GND_net), .O(n30_adj_4973));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48895_4_lut (.I0(n455[16]), .I1(n71822), .I2(n46[16]), .I3(n69209), 
            .O(n68165));
    defparam i48895_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i51540_3_lut (.I0(n70809), .I1(n285[18]), .I2(n37_adj_4886), 
            .I3(GND_net), .O(n70810));   // verilog/motorControl.v(58[23:46])
    defparam i51540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51520_3_lut (.I0(n70810), .I1(n285[19]), .I2(n39_adj_4882), 
            .I3(GND_net), .O(n70790));   // verilog/motorControl.v(58[23:46])
    defparam i51520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51092_4_lut (.I0(n30_adj_4973), .I1(n10_adj_4972), .I2(n71848), 
            .I3(n68151), .O(n70362));   // verilog/motorControl.v(62[35:55])
    defparam i51092_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 n71266_bdd_4_lut (.I0(n71266), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4751), .O(n71269));
    defparam n71266_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49726_3_lut (.I0(n69875), .I1(n46[15]), .I2(n455[15]), .I3(GND_net), 
            .O(n68996));   // verilog/motorControl.v(62[35:55])
    defparam i49726_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49049_4_lut (.I0(n43_adj_4884), .I1(n41_adj_4883), .I2(n39_adj_4882), 
            .I3(n70712), .O(n68319));
    defparam i49049_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51448_4_lut (.I0(n68996), .I1(n70362), .I2(n71848), .I3(n68165), 
            .O(n70718));   // verilog/motorControl.v(62[35:55])
    defparam i51448_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51169_4_lut (.I0(n68974), .I1(n69784), .I2(n45_adj_4880), 
            .I3(n68315), .O(n70439));   // verilog/motorControl.v(58[23:46])
    defparam i51169_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51449_3_lut (.I0(n70718), .I1(n46[18]), .I2(n455[18]), .I3(GND_net), 
            .O(n70719));   // verilog/motorControl.v(62[35:55])
    defparam i51449_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51435_3_lut (.I0(n70719), .I1(n46[19]), .I2(n455[19]), .I3(GND_net), 
            .O(n70705));   // verilog/motorControl.v(62[35:55])
    defparam i51435_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i6_3_lut (.I0(n46[2]), .I1(n46[3]), .I2(n455[3]), 
            .I3(GND_net), .O(n6_adj_4974));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49712_3_lut (.I0(n70790), .I1(n285[20]), .I2(n41_adj_4883), 
            .I3(GND_net), .O(n68982));   // verilog/motorControl.v(58[23:46])
    defparam i49712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50608_3_lut (.I0(n6_adj_4974), .I1(n46[10]), .I2(n455[10]), 
            .I3(GND_net), .O(n69878));   // verilog/motorControl.v(62[35:55])
    defparam i50608_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50609_3_lut (.I0(n69878), .I1(n46[11]), .I2(n455[11]), .I3(GND_net), 
            .O(n69879));   // verilog/motorControl.v(62[35:55])
    defparam i50609_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48852_4_lut (.I0(n455[21]), .I1(n71837), .I2(n46[21]), .I3(n69229), 
            .O(n68122));
    defparam i48852_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i51413_4_lut (.I0(n68982), .I1(n70439), .I2(n45_adj_4880), 
            .I3(n68319), .O(n70683));   // verilog/motorControl.v(58[23:46])
    defparam i51413_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51414_3_lut (.I0(n70683), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i51414_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i45_rep_99_2_lut (.I0(n455[22]), .I1(n46[22]), .I2(GND_net), 
            .I3(GND_net), .O(n71810));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_rep_99_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n335[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50518_4_lut (.I0(n24_adj_4958), .I1(n8_adj_4957), .I2(n71810), 
            .I3(n68120), .O(n69788));   // verilog/motorControl.v(62[35:55])
    defparam i50518_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49724_3_lut (.I0(n69879), .I1(n46[12]), .I2(n455[12]), .I3(GND_net), 
            .O(n68994));   // verilog/motorControl.v(62[35:55])
    defparam i49724_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48863_4_lut (.I0(n455[21]), .I1(n71813), .I2(n46[21]), .I3(n70770), 
            .O(n68133));
    defparam i48863_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i51173_4_lut (.I0(n68994), .I1(n69788), .I2(n71810), .I3(n68122), 
            .O(n70443));   // verilog/motorControl.v(62[35:55])
    defparam i51173_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49732_3_lut (.I0(n70705), .I1(n46[20]), .I2(n455[20]), .I3(GND_net), 
            .O(n69002));   // verilog/motorControl.v(62[35:55])
    defparam i49732_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51417_4_lut (.I0(n69002), .I1(n70443), .I2(n71810), .I3(n68133), 
            .O(n70687));   // verilog/motorControl.v(62[35:55])
    defparam i51417_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_4975));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50988_3_lut (.I0(n4_adj_4975), .I1(n455[13]), .I2(n27_adj_4955), 
            .I3(GND_net), .O(n70258));   // verilog/motorControl.v(62[14:31])
    defparam i50988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50989_3_lut (.I0(n70258), .I1(n455[14]), .I2(n29_adj_4940), 
            .I3(GND_net), .O(n70259));   // verilog/motorControl.v(62[14:31])
    defparam i50989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49000_4_lut (.I0(n33_adj_4951), .I1(n31_adj_4941), .I2(n29_adj_4940), 
            .I3(n68278), .O(n68270));
    defparam i49000_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51329_4_lut (.I0(n30_adj_4966), .I1(n10_adj_4965), .I2(n35_adj_4950), 
            .I3(n68264), .O(n70599));   // verilog/motorControl.v(62[14:31])
    defparam i51329_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49716_3_lut (.I0(n70259), .I1(n455[15]), .I2(n31_adj_4941), 
            .I3(GND_net), .O(n68986));   // verilog/motorControl.v(62[14:31])
    defparam i49716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51541_4_lut (.I0(n68986), .I1(n70599), .I2(n35_adj_4950), 
            .I3(n68270), .O(n70811));   // verilog/motorControl.v(62[14:31])
    defparam i51541_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9980_bdd_4_lut_51981 (.I0(n9980), .I1(n67569), .I2(setpoint[16]), 
            .I3(n4751), .O(n71260));
    defparam n9980_bdd_4_lut_51981.LUT_INIT = 16'he4aa;
    SB_LUT4 i51542_3_lut (.I0(n70811), .I1(n455[18]), .I2(n37_adj_4943), 
            .I3(GND_net), .O(n70812));   // verilog/motorControl.v(62[14:31])
    defparam i51542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51518_3_lut (.I0(n70812), .I1(n455[19]), .I2(n39_adj_4938), 
            .I3(GND_net), .O(n70788));   // verilog/motorControl.v(62[14:31])
    defparam i51518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48981_4_lut (.I0(n43_adj_4942), .I1(n41_adj_4937), .I2(n39_adj_4938), 
            .I3(n70708), .O(n68251));
    defparam i48981_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51171_4_lut (.I0(n68984), .I1(n69786), .I2(n45_adj_4939), 
            .I3(n68236), .O(n70441));   // verilog/motorControl.v(62[14:31])
    defparam i51171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49722_3_lut (.I0(n70788), .I1(n455[20]), .I2(n41_adj_4937), 
            .I3(GND_net), .O(n68992));   // verilog/motorControl.v(62[14:31])
    defparam i49722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51418_3_lut (.I0(n70687), .I1(n455[23]), .I2(n47_adj_4678), 
            .I3(GND_net), .O(n70688));   // verilog/motorControl.v(62[35:55])
    defparam i51418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71260_bdd_4_lut (.I0(n71260), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4751), .O(n71263));
    defparam n71260_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51415_4_lut (.I0(n68992), .I1(n70441), .I2(n45_adj_4939), 
            .I3(n68251), .O(n70685));   // verilog/motorControl.v(62[14:31])
    defparam i51415_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i23694_4_lut (.I0(n70685), .I1(n70688), .I2(deadband[23]), 
            .I3(n455[23]), .O(n41540));
    defparam i23694_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 i34417_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n23138[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34417_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i34419_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n52224));   // verilog/motorControl.v(61[29:40])
    defparam i34419_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i34446_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n23117[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34446_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i34448_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n52254));   // verilog/motorControl.v(61[29:40])
    defparam i34448_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i34589_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4976), 
            .I3(n23080[1]), .O(n6_adj_4828));   // verilog/motorControl.v(61[29:40])
    defparam i34589_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_986 (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4976), 
            .I3(n23080[1]), .O(n23023[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_986.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_987 (.I0(\Ki[2] ), .I1(n335[18]), .I2(n52388), 
            .I3(n23080[0]), .O(n23023[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_987.LUT_INIT = 16'h8778;
    SB_LUT4 i34581_3_lut_4_lut (.I0(\Ki[2] ), .I1(n335[18]), .I2(n52388), 
            .I3(n23080[0]), .O(n4_adj_4976));   // verilog/motorControl.v(61[29:40])
    defparam i34581_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4526));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34568_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n23023[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34568_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i34570_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n52388));   // verilog/motorControl.v(61[29:40])
    defparam i34570_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut_4_lut_adj_988 (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4977), 
            .I3(n23117[1]), .O(n23080[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_988.LUT_INIT = 16'h8778;
    SB_LUT4 i34514_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4977), 
            .I3(n23117[1]), .O(n6_adj_4838));   // verilog/motorControl.v(61[29:40])
    defparam i34514_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34506_3_lut_4_lut (.I0(n62_adj_4830), .I1(n131), .I2(n204), 
            .I3(n23117[0]), .O(n4_adj_4977));   // verilog/motorControl.v(61[29:40])
    defparam i34506_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_989 (.I0(n62_adj_4830), .I1(n131), .I2(n204), 
            .I3(n23117[0]), .O(n23080[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_989.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4978));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4979));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4525));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i45_2_lut (.I0(PWMLimit[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4980));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i43_2_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4981));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4982));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4983));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4984));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i23_2_lut (.I0(PWMLimit[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4985));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i25_2_lut (.I0(PWMLimit[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4986));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4987));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4988));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4989));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9980_bdd_4_lut_51976 (.I0(n9980), .I1(n67568), .I2(setpoint[15]), 
            .I3(n4751), .O(n71254));
    defparam n9980_bdd_4_lut_51976.LUT_INIT = 16'he4aa;
    SB_LUT4 n71254_bdd_4_lut (.I0(n71254), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4751), .O(n71257));
    defparam n71254_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9980_bdd_4_lut_51971 (.I0(n9980), .I1(n67567), .I2(setpoint[14]), 
            .I3(n4751), .O(n71248));
    defparam n9980_bdd_4_lut_51971.LUT_INIT = 16'he4aa;
    SB_LUT4 n71248_bdd_4_lut (.I0(n71248), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4751), .O(n71251));
    defparam n71248_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4990));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9980_bdd_4_lut_51966 (.I0(n9980), .I1(n67566), .I2(setpoint[13]), 
            .I3(n4751), .O(n71242));
    defparam n9980_bdd_4_lut_51966.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4991));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4992));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i9_2_lut (.I0(PWMLimit[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4993));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4994));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4995));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n71242_bdd_4_lut (.I0(n71242), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4751), .O(n71245));
    defparam n71242_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i21_2_lut (.I0(PWMLimit[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4996));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48802_4_lut (.I0(n21_adj_4996), .I1(n19_adj_4995), .I2(n17_adj_4994), 
            .I3(n9_adj_4993), .O(n68072));
    defparam i48802_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9980_bdd_4_lut_51961 (.I0(n9980), .I1(n67565), .I2(setpoint[12]), 
            .I3(n4751), .O(n71236));
    defparam n9980_bdd_4_lut_51961.LUT_INIT = 16'he4aa;
    SB_LUT4 n71236_bdd_4_lut (.I0(n71236), .I1(n535[12]), .I2(n455[12]), 
            .I3(n4751), .O(n71239));
    defparam n71236_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9980_bdd_4_lut_51956 (.I0(n9980), .I1(n67564), .I2(setpoint[11]), 
            .I3(n4751), .O(n71230));
    defparam n9980_bdd_4_lut_51956.LUT_INIT = 16'he4aa;
    SB_LUT4 n71230_bdd_4_lut (.I0(n71230), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4751), .O(n71233));
    defparam n71230_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48766_4_lut (.I0(n27_adj_4992), .I1(n15_adj_4991), .I2(n13_adj_4990), 
            .I3(n11_adj_4989), .O(n68036));
    defparam i48766_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4988), 
            .I3(GND_net), .O(n12_adj_4997));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4990), 
            .I3(GND_net), .O(n10_adj_4998));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n12_adj_4997), .I1(n455[17]), .I2(n35_adj_4987), 
            .I3(GND_net), .O(n30_adj_4999));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49796_4_lut (.I0(n13_adj_4990), .I1(n11_adj_4989), .I2(n9_adj_4993), 
            .I3(n68118), .O(n69066));
    defparam i49796_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49792_4_lut (.I0(n19_adj_4995), .I1(n17_adj_4994), .I2(n15_adj_4991), 
            .I3(n69066), .O(n69062));
    defparam i49792_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51199_4_lut (.I0(n25_adj_4986), .I1(n23_adj_4985), .I2(n21_adj_4996), 
            .I3(n69062), .O(n70469));
    defparam i51199_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n9980_bdd_4_lut_51951 (.I0(n9980), .I1(n67563), .I2(setpoint[10]), 
            .I3(n4751), .O(n71224));
    defparam n9980_bdd_4_lut_51951.LUT_INIT = 16'he4aa;
    SB_LUT4 i50534_4_lut (.I0(n31_adj_4984), .I1(n29_adj_4983), .I2(n27_adj_4992), 
            .I3(n70469), .O(n69804));
    defparam i50534_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51419_4_lut (.I0(n37_adj_4982), .I1(n35_adj_4987), .I2(n33_adj_4988), 
            .I3(n69804), .O(n70689));
    defparam i51419_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4981), 
            .I3(GND_net), .O(n16_adj_5000));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71224_bdd_4_lut (.I0(n71224), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4751), .O(n71227));
    defparam n71224_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50596_3_lut (.I0(n6), .I1(n455[10]), .I2(n21_adj_4996), .I3(GND_net), 
            .O(n69866));   // verilog/motorControl.v(63[16:31])
    defparam i50596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9980_bdd_4_lut_51946 (.I0(n9980), .I1(n67559), .I2(setpoint[9]), 
            .I3(n4751), .O(n71218));
    defparam n9980_bdd_4_lut_51946.LUT_INIT = 16'he4aa;
    SB_LUT4 i50597_3_lut (.I0(n69866), .I1(n455[11]), .I2(n23_adj_4985), 
            .I3(GND_net), .O(n69867));   // verilog/motorControl.v(63[16:31])
    defparam i50597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4994), 
            .I3(GND_net), .O(n8_adj_5001));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71218_bdd_4_lut (.I0(n71218), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4751), .O(n71221));
    defparam n71218_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_30_i24_3_lut (.I0(n16_adj_5000), .I1(n455[22]), .I2(n45_adj_4980), 
            .I3(GND_net), .O(n24_adj_5002));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9980_bdd_4_lut_51941 (.I0(n9980), .I1(n67558), .I2(setpoint[8]), 
            .I3(n4751), .O(n71212));
    defparam n9980_bdd_4_lut_51941.LUT_INIT = 16'he4aa;
    SB_LUT4 n71212_bdd_4_lut (.I0(n71212), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4751), .O(n71215));
    defparam n71212_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48676_4_lut (.I0(n43_adj_4981), .I1(n25_adj_4986), .I2(n23_adj_4985), 
            .I3(n68072), .O(n67946));
    defparam i48676_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9980_bdd_4_lut_51936 (.I0(n9980), .I1(n67557), .I2(setpoint[7]), 
            .I3(n4751), .O(n71206));
    defparam n9980_bdd_4_lut_51936.LUT_INIT = 16'he4aa;
    SB_LUT4 i50520_4_lut (.I0(n24_adj_5002), .I1(n8_adj_5001), .I2(n45_adj_4980), 
            .I3(n67934), .O(n69790));   // verilog/motorControl.v(63[16:31])
    defparam i50520_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49734_3_lut (.I0(n69867), .I1(n455[12]), .I2(n25_adj_4986), 
            .I3(GND_net), .O(n69004));   // verilog/motorControl.v(63[16:31])
    defparam i49734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_5003));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i50594_3_lut (.I0(n4_adj_5003), .I1(n455[13]), .I2(n27_adj_4992), 
            .I3(GND_net), .O(n69864));   // verilog/motorControl.v(63[16:31])
    defparam i50594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50595_3_lut (.I0(n69864), .I1(n455[14]), .I2(n29_adj_4983), 
            .I3(GND_net), .O(n69865));   // verilog/motorControl.v(63[16:31])
    defparam i50595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48739_4_lut (.I0(n33_adj_4988), .I1(n31_adj_4984), .I2(n29_adj_4983), 
            .I3(n68036), .O(n68009));
    defparam i48739_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n71206_bdd_4_lut (.I0(n71206), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4751), .O(n71209));
    defparam n71206_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51450_4_lut (.I0(n30_adj_4999), .I1(n10_adj_4998), .I2(n35_adj_4987), 
            .I3(n68007), .O(n70720));   // verilog/motorControl.v(63[16:31])
    defparam i51450_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49736_3_lut (.I0(n69865), .I1(n455[15]), .I2(n31_adj_4984), 
            .I3(GND_net), .O(n69006));   // verilog/motorControl.v(63[16:31])
    defparam i49736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51599_4_lut (.I0(n69006), .I1(n70720), .I2(n35_adj_4987), 
            .I3(n68009), .O(n70869));   // verilog/motorControl.v(63[16:31])
    defparam i51599_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51600_3_lut (.I0(n70869), .I1(n455[18]), .I2(n37_adj_4982), 
            .I3(GND_net), .O(n70870));   // verilog/motorControl.v(63[16:31])
    defparam i51600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51562_3_lut (.I0(n70870), .I1(n455[19]), .I2(n39_adj_4978), 
            .I3(GND_net), .O(n70832));   // verilog/motorControl.v(63[16:31])
    defparam i51562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48678_4_lut (.I0(n43_adj_4981), .I1(n41_adj_4979), .I2(n39_adj_4978), 
            .I3(n70689), .O(n67948));
    defparam i48678_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51177_4_lut (.I0(n69004), .I1(n69790), .I2(n45_adj_4980), 
            .I3(n67946), .O(n70447));   // verilog/motorControl.v(63[16:31])
    defparam i51177_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51487_3_lut (.I0(n70832), .I1(n455[20]), .I2(n41_adj_4979), 
            .I3(GND_net), .O(n40_adj_5004));   // verilog/motorControl.v(63[16:31])
    defparam i51487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51179_4_lut (.I0(n40_adj_5004), .I1(n70447), .I2(n45_adj_4980), 
            .I3(n67948), .O(n70449));   // verilog/motorControl.v(63[16:31])
    defparam i51179_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49139_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n68409));   // verilog/motorControl.v(58[23:46])
    defparam i49139_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4960));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49208_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n68478));   // verilog/motorControl.v(56[14:36])
    defparam i49208_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_adj_4840));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i3_4_lut (.I0(n59660), .I1(n27602), .I2(control_update), .I3(n105), 
            .O(n7073));
    defparam i3_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i3_4_lut_adj_990 (.I0(n7071), .I1(n7073), .I2(n27508), .I3(n41850), 
            .O(n4751));
    defparam i3_4_lut_adj_990.LUT_INIT = 16'hefff;
    SB_LUT4 i48589_4_lut (.I0(n27_adj_4913), .I1(n15_adj_4912), .I2(n13_adj_4909), 
            .I3(n11_adj_4908), .O(n67859));
    defparam i48589_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4903), 
            .I3(GND_net), .O(n12_adj_5005));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4909), 
            .I3(GND_net), .O(n10_adj_5006));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_5005), .I1(n535[17]), .I2(n35_adj_4902), 
            .I3(GND_net), .O(n30_adj_5007));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49619_4_lut (.I0(n13_adj_4909), .I1(n11_adj_4908), .I2(n9_adj_4900), 
            .I3(n67926), .O(n68889));
    defparam i49619_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49613_4_lut (.I0(n19_adj_4896), .I1(n17_adj_4895), .I2(n15_adj_4912), 
            .I3(n68889), .O(n68883));
    defparam i49613_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51145_4_lut (.I0(n25_adj_4899), .I1(n23_adj_4898), .I2(n21_adj_4897), 
            .I3(n68883), .O(n70415));
    defparam i51145_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50450_4_lut (.I0(n31_adj_4892), .I1(n29_adj_4891), .I2(n27_adj_4913), 
            .I3(n70415), .O(n69720));
    defparam i50450_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51401_4_lut (.I0(n37_adj_4894), .I1(n35_adj_4902), .I2(n33_adj_4903), 
            .I3(n69720), .O(n70671));
    defparam i51401_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51090_3_lut (.I0(n6_adj_4872), .I1(n535[10]), .I2(n21_adj_4897), 
            .I3(GND_net), .O(n70360));   // verilog/motorControl.v(65[25:41])
    defparam i51090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51091_3_lut (.I0(n70360), .I1(n535[11]), .I2(n23_adj_4898), 
            .I3(GND_net), .O(n70361));   // verilog/motorControl.v(65[25:41])
    defparam i51091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4888), 
            .I3(GND_net), .O(n16_adj_5008));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4895), 
            .I3(GND_net), .O(n8_adj_5009));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_5008), .I1(n535[22]), .I2(n45_c), 
            .I3(GND_net), .O(n24_adj_5010));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48616_4_lut (.I0(n21_adj_4897), .I1(n19_adj_4896), .I2(n17_adj_4895), 
            .I3(n9_adj_4900), .O(n67886));
    defparam i48616_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48565_4_lut (.I0(n43_adj_4888), .I1(n25_adj_4899), .I2(n23_adj_4898), 
            .I3(n67886), .O(n67835));
    defparam i48565_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50522_4_lut (.I0(n24_adj_5010), .I1(n8_adj_5009), .I2(n45_c), 
            .I3(n67833), .O(n69792));   // verilog/motorControl.v(65[25:41])
    defparam i50522_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50862_3_lut (.I0(n70361), .I1(n535[12]), .I2(n25_adj_4899), 
            .I3(GND_net), .O(n70132));   // verilog/motorControl.v(65[25:41])
    defparam i50862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_5011));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51086_3_lut (.I0(n4_adj_5011), .I1(n535[13]), .I2(n27_adj_4913), 
            .I3(GND_net), .O(n70356));   // verilog/motorControl.v(65[25:41])
    defparam i51086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51087_3_lut (.I0(n70356), .I1(n535[14]), .I2(n29_adj_4891), 
            .I3(GND_net), .O(n70357));   // verilog/motorControl.v(65[25:41])
    defparam i51087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48577_4_lut (.I0(n33_adj_4903), .I1(n31_adj_4892), .I2(n29_adj_4891), 
            .I3(n67859), .O(n67847));
    defparam i48577_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51452_4_lut (.I0(n30_adj_5007), .I1(n10_adj_5006), .I2(n35_adj_4902), 
            .I3(n67845), .O(n70722));   // verilog/motorControl.v(65[25:41])
    defparam i51452_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50864_3_lut (.I0(n70357), .I1(n535[15]), .I2(n31_adj_4892), 
            .I3(GND_net), .O(n70134));   // verilog/motorControl.v(65[25:41])
    defparam i50864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51601_4_lut (.I0(n70134), .I1(n70722), .I2(n35_adj_4902), 
            .I3(n67847), .O(n70871));   // verilog/motorControl.v(65[25:41])
    defparam i51601_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51602_3_lut (.I0(n70871), .I1(n535[18]), .I2(n37_adj_4894), 
            .I3(GND_net), .O(n70872));   // verilog/motorControl.v(65[25:41])
    defparam i51602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51560_3_lut (.I0(n70872), .I1(n535[19]), .I2(n39_adj_4887), 
            .I3(GND_net), .O(n70830));   // verilog/motorControl.v(65[25:41])
    defparam i51560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48569_4_lut (.I0(n43_adj_4888), .I1(n41_adj_4885), .I2(n39_adj_4887), 
            .I3(n70671), .O(n67839));
    defparam i48569_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50867_4_lut (.I0(n70132), .I1(n69792), .I2(n45_c), .I3(n67835), 
            .O(n70137));   // verilog/motorControl.v(65[25:41])
    defparam i50867_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51489_3_lut (.I0(n70830), .I1(n535[20]), .I2(n41_adj_4885), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(65[25:41])
    defparam i51489_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (enable_slow_N_4213, clk16MHz, n29874, data, ID, GND_net, 
            baudrate, n31646, n31645, n31644, n31643, n31642, n31641, 
            n31640, n31639, \state_7__N_3918[0] , data_ready, \state_7__N_4110[0] , 
            \state[0] , scl_enable, VCC_net, sda_enable, n32362, n32360, 
            n32356, n32339, n32338, n32337, n32335, n32065, n8, 
            n6722, scl, sda_out, \state_7__N_4126[3] , n41430, n6, 
            n4, n4_adj_3, n41590, n10, n27672, n27624) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output enable_slow_N_4213;
    input clk16MHz;
    output n29874;
    output [7:0]data;
    output [7:0]ID;
    input GND_net;
    output [31:0]baudrate;
    input n31646;
    input n31645;
    input n31644;
    input n31643;
    input n31642;
    input n31641;
    input n31640;
    input n31639;
    input \state_7__N_3918[0] ;
    output data_ready;
    output \state_7__N_4110[0] ;
    output \state[0] ;
    output scl_enable;
    input VCC_net;
    output sda_enable;
    input n32362;
    input n32360;
    input n32356;
    input n32339;
    input n32338;
    input n32337;
    input n32335;
    input n32065;
    input n8;
    output n6722;
    output scl;
    output sda_out;
    input \state_7__N_4126[3] ;
    output n41430;
    output n6;
    output n4;
    output n4_adj_3;
    output n41590;
    output n10;
    output n27672;
    output n27624;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire n3, n50803, n29791;
    wire [7:0]state_7__N_3885;
    
    wire ready_prev;
    wire [0:0]n5942;
    
    wire enable, n41452;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    wire [2:0]n17;
    
    wire n23732, n62518;
    wire [15:0]delay_counter_15__N_3956;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n15, n31466, n31671, n6946, n6948, n6949, n6950, n6951, 
        n6952, n31672, n31673, n31674, n31675, n31676, n31677, 
        n50789, n64383, n41842, n54769, n29983, n31409, n31670, 
        n31669, n31668, n31667, n31666, n31665, n31664, n31663, 
        n31662, n31661, n31660, n31659, n59022, n59026, n59024, 
        n59020, n31654, n31653, n31652, n31651, n31650, n31649, 
        n31648, n31647, n4_c, n64433, n27499;
    wire [7:0]state_adj_4447;   // verilog/i2c_controller.v(33[12:17])
    
    wire n67788, n59032, rw, n31470, n32383, n59192;
    wire [15:0]n5408;
    
    wire n52803, n52802, n52801, n52800, n52799, n52798, n50775, 
        n52797, n52796, n52795, n52794, n52793, n52792, n52791, 
        n52790, n52789, n62688, n16, n22, n20, n24, n54190, 
        n4_adj_4441, n12, n67779, n29797, n4_adj_4442, n10_c;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n59552;
    
    SB_LUT4 i1_4_lut_4_lut (.I0(state[2]), .I1(n3), .I2(state[0]), .I3(state[1]), 
            .O(n50803));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0052;
    SB_LUT4 i25_4_lut_4_lut (.I0(state[2]), .I1(n3), .I2(state[1]), .I3(state[0]), 
            .O(n29791));   // verilog/eeprom.v(27[11:16])
    defparam i25_4_lut_4_lut.LUT_INIT = 16'h0552;
    SB_LUT4 i1_4_lut_4_lut_adj_955 (.I0(state[2]), .I1(n3), .I2(state[1]), 
            .I3(state[0]), .O(state_7__N_3885[1]));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_4_lut_adj_955.LUT_INIT = 16'ha5f2;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5942[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i34539_3_lut_4_lut (.I0(n41452), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i34539_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i3_4_lut (.I0(byte_counter[1]), .I1(n23732), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n29874));
    defparam i3_4_lut.LUT_INIT = 16'h0010;
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n62518), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n29791), 
            .D(delay_counter_15__N_3956[1]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13521_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(ID[0]), .O(n31466));
    defparam i13521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n29791), 
            .D(delay_counter_15__N_3956[2]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i33381_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(ID[7]), .O(n31671));
    defparam i33381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n29791), 
            .D(delay_counter_15__N_3956[3]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n29791), 
            .D(n6946), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n29791), 
            .D(delay_counter_15__N_3956[5]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n29791), 
            .D(n6948), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n29791), 
            .D(n6949), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n29791), 
            .D(n6950), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n29791), 
            .D(n6951), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n29791), .D(n6952), .S(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n29791), .D(delay_counter_15__N_3956[11]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n29791), .D(delay_counter_15__N_3956[12]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n29791), .D(delay_counter_15__N_3956[13]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13727_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(ID[6]), .O(n31672));
    defparam i13727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n29791), .D(delay_counter_15__N_3956[14]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n29791), .D(delay_counter_15__N_3956[15]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13728_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(ID[5]), .O(n31673));
    defparam i13728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13729_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(ID[4]), .O(n31674));
    defparam i13729_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13730_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(ID[3]), .O(n31675));
    defparam i13730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13731_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(ID[2]), .O(n31676));
    defparam i13731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13732_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(ID[1]), .O(n31677));
    defparam i13732_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(byte_counter[2]), .I1(n23732), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n50789));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_956 (.I0(byte_counter[2]), .I1(n23732), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n15));
    defparam i1_2_lut_3_lut_adj_956.LUT_INIT = 16'hfefe;
    SB_LUT4 i45124_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n64383));
    defparam i45124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(state[2]), .I1(n41842), .I2(ready_prev), .I3(n64383), 
            .O(n23732));
    defparam i4_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFESR byte_counter_2048__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n29983), .D(n54769), .R(n31409));   // verilog/eeprom.v(68[25:39])
    SB_LUT4 i13725_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(baudrate[0]), .O(n31670));   // verilog/eeprom.v(68[25:39])
    defparam i13725_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13724_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(baudrate[1]), .O(n31669));   // verilog/eeprom.v(68[25:39])
    defparam i13724_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESR byte_counter_2048__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n29983), .D(n17[2]), .R(n31409));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2048__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n29983), .D(n17[1]), .R(n31409));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n31677));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n31676));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n31675));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n31674));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n31673));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n31672));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n31671));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n31670));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n31669));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n31668));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n31667));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n31666));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n31665));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n31664));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n31663));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n31662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n31661));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n31660));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n31659));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n59022));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n59026));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n59024));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n59020));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n31654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n31653));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n31652));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n31651));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n31650));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n31649));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n31648));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n31647));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n31646));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n31645));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n31644));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n31643));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n31642));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n31641));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n31640));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n31639));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13723_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(baudrate[2]), .O(n31668));   // verilog/eeprom.v(68[25:39])
    defparam i13723_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13722_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(baudrate[3]), .O(n31667));   // verilog/eeprom.v(68[25:39])
    defparam i13722_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13721_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(baudrate[4]), .O(n31666));   // verilog/eeprom.v(68[25:39])
    defparam i13721_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13720_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(baudrate[5]), .O(n31665));   // verilog/eeprom.v(68[25:39])
    defparam i13720_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13719_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(baudrate[6]), .O(n31664));   // verilog/eeprom.v(68[25:39])
    defparam i13719_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13718_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(baudrate[7]), .O(n31663));   // verilog/eeprom.v(68[25:39])
    defparam i13718_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n29791), 
            .D(delay_counter_15__N_3956[0]), .R(n50803));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i23607_2_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n41452));
    defparam i23607_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n3));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut (.I0(state[2]), .I1(state[1]), .I2(\state_7__N_3918[0] ), 
            .I3(state[0]), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'hbbba;
    SB_LUT4 i49478_4_lut (.I0(n64433), .I1(n27499), .I2(state[1]), .I3(state_adj_4447[3]), 
            .O(n67788));
    defparam i49478_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n67788), .I1(n4_c), .I2(n41452), .I3(state[0]), 
            .O(n62518));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n59032));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n31470));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n32383));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n31466));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n59192));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1200_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5408[9]), 
            .I3(n52803), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1200_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5408[9]), 
            .I3(n52802), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_16 (.CI(n52802), .I0(delay_counter[14]), .I1(n5408[9]), 
            .CO(n52803));
    SB_LUT4 add_1200_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5408[9]), 
            .I3(n52801), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_15 (.CI(n52801), .I0(delay_counter[13]), .I1(n5408[9]), 
            .CO(n52802));
    SB_LUT4 add_1200_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5408[9]), 
            .I3(n52800), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_14 (.CI(n52800), .I0(delay_counter[12]), .I1(n5408[9]), 
            .CO(n52801));
    SB_LUT4 add_1200_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5408[9]), 
            .I3(n52799), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_13 (.CI(n52799), .I0(delay_counter[11]), .I1(n5408[9]), 
            .CO(n52800));
    SB_LUT4 add_1200_12_lut (.I0(n50775), .I1(delay_counter[10]), .I2(n5408[9]), 
            .I3(n52798), .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_12 (.CI(n52798), .I0(delay_counter[10]), .I1(n5408[9]), 
            .CO(n52799));
    SB_LUT4 add_1200_11_lut (.I0(n50775), .I1(delay_counter[9]), .I2(n5408[9]), 
            .I3(n52797), .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_11 (.CI(n52797), .I0(delay_counter[9]), .I1(n5408[9]), 
            .CO(n52798));
    SB_LUT4 add_1200_10_lut (.I0(n50775), .I1(delay_counter[8]), .I2(n5408[9]), 
            .I3(n52796), .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_10 (.CI(n52796), .I0(delay_counter[8]), .I1(n5408[9]), 
            .CO(n52797));
    SB_LUT4 add_1200_9_lut (.I0(n50775), .I1(delay_counter[7]), .I2(n5408[9]), 
            .I3(n52795), .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_9 (.CI(n52795), .I0(delay_counter[7]), .I1(n5408[9]), 
            .CO(n52796));
    SB_LUT4 add_1200_8_lut (.I0(n50775), .I1(delay_counter[6]), .I2(n5408[9]), 
            .I3(n52794), .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_8 (.CI(n52794), .I0(delay_counter[6]), .I1(n5408[9]), 
            .CO(n52795));
    SB_LUT4 add_1200_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5408[9]), 
            .I3(n52793), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_7 (.CI(n52793), .I0(delay_counter[5]), .I1(n5408[9]), 
            .CO(n52794));
    SB_LUT4 add_1200_6_lut (.I0(n50775), .I1(delay_counter[4]), .I2(n5408[9]), 
            .I3(n52792), .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1200_6 (.CI(n52792), .I0(delay_counter[4]), .I1(n5408[9]), 
            .CO(n52793));
    SB_LUT4 add_1200_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5408[9]), 
            .I3(n52791), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_5 (.CI(n52791), .I0(delay_counter[3]), .I1(n5408[9]), 
            .CO(n52792));
    SB_LUT4 add_1200_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5408[9]), 
            .I3(n52790), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_4 (.CI(n52790), .I0(delay_counter[2]), .I1(n5408[9]), 
            .CO(n52791));
    SB_LUT4 add_1200_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5408[9]), 
            .I3(n52789), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_3 (.CI(n52789), .I0(delay_counter[1]), .I1(n5408[9]), 
            .CO(n52790));
    SB_LUT4 add_1200_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5408[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1200_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1200_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5408[9]), 
            .CO(n52789));
    SB_LUT4 i3_4_lut_adj_957 (.I0(delay_counter[4]), .I1(delay_counter[10]), 
            .I2(delay_counter[5]), .I3(delay_counter[8]), .O(n62688));   // verilog/eeprom.v(55[12:28])
    defparam i3_4_lut_adj_957.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(delay_counter[12]), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/eeprom.v(55[12:28])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(delay_counter[9]), .I1(delay_counter[11]), .I2(delay_counter[7]), 
            .I3(delay_counter[14]), .O(n22));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(delay_counter[3]), .I1(n62688), .I2(delay_counter[13]), 
            .I3(GND_net), .O(n20));   // verilog/eeprom.v(55[12:28])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[0]), .I1(n22), .I2(n16), .I3(delay_counter[2]), 
            .O(n24));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(delay_counter[15]), .I1(n24), .I2(n20), .I3(delay_counter[1]), 
            .O(n27499));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n27499), .I1(state[0]), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n54190));
    defparam i2_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_4_lut_adj_958 (.I0(state[0]), .I1(state[2]), .I2(\state_7__N_3918[0] ), 
            .I3(state[1]), .O(n31409));   // verilog/eeprom.v(68[25:39])
    defparam i2_4_lut_adj_958.LUT_INIT = 16'h0010;
    SB_LUT4 i1_4_lut_adj_959 (.I0(state[2]), .I1(\state_7__N_3918[0] ), 
            .I2(state[1]), .I3(state[0]), .O(n29983));
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h5004;
    SB_LUT4 i13_2_lut (.I0(state[2]), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n50775));
    defparam i13_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i51691_2_lut (.I0(n27499), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5408[9]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i51691_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30_4_lut (.I0(\state_7__N_3918[0] ), .I1(n27499), .I2(state[1]), 
            .I3(n4_adj_4441), .O(n12));
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12), .I1(n67779), .I2(state[0]), .I3(state[2]), 
            .O(n59192));
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i49443_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(state[1]), .I3(GND_net), .O(n67779));
    defparam i49443_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_960 (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n54769));
    defparam i1_2_lut_3_lut_adj_960.LUT_INIT = 16'hd2d2;
    SB_LUT4 mux_1517_Mux_0_i3_3_lut_4_lut (.I0(state[0]), .I1(n27499), .I2(enable_slow_N_4213), 
            .I3(state[1]), .O(n5942[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1517_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h10aa;
    SB_LUT4 i1_4_lut_adj_961 (.I0(state[1]), .I1(state[0]), .I2(n41452), 
            .I3(state[2]), .O(n32383));
    defparam i1_4_lut_adj_961.LUT_INIT = 16'hee08;
    SB_LUT4 i2_4_lut_adj_962 (.I0(state[0]), .I1(n3), .I2(state[1]), .I3(state[2]), 
            .O(n29797));
    defparam i2_4_lut_adj_962.LUT_INIT = 16'h0405;
    SB_LUT4 i1_2_lut (.I0(state[2]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4442));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i14_4_lut (.I0(n29797), .I1(state[1]), .I2(data_ready), .I3(n4_adj_4442), 
            .O(n31470));   // verilog/eeprom.v(27[11:16])
    defparam i14_4_lut.LUT_INIT = 16'h5072;
    SB_LUT4 i1_4_lut_adj_963 (.I0(state[1]), .I1(rw), .I2(n54190), .I3(state[2]), 
            .O(n10_c));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h888a;
    SB_LUT4 i1_4_lut_adj_964 (.I0(n10_c), .I1(rw), .I2(state[0]), .I3(state[2]), 
            .O(n59032));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_964.LUT_INIT = 16'heeae;
    SB_LUT4 i1_4_lut_adj_965 (.I0(\state_7__N_4110[0] ), .I1(saved_addr[0]), 
            .I2(rw), .I3(n41842), .O(n59552));   // verilog/i2c_controller.v(34[12:22])
    defparam i1_4_lut_adj_965.LUT_INIT = 16'hcce4;
    SB_LUT4 i13714_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[3]), 
            .I3(baudrate[11]), .O(n31659));   // verilog/eeprom.v(68[25:39])
    defparam i13714_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13717_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[0]), 
            .I3(baudrate[8]), .O(n31662));   // verilog/eeprom.v(68[25:39])
    defparam i13717_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13715_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[2]), 
            .I3(baudrate[10]), .O(n31660));   // verilog/eeprom.v(68[25:39])
    defparam i13715_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13716_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[1]), 
            .I3(baudrate[9]), .O(n31661));   // verilog/eeprom.v(68[25:39])
    defparam i13716_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[4]), 
            .I3(baudrate[12]), .O(n59022));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_966 (.I0(byte_counter[0]), .I1(n50789), 
            .I2(data[5]), .I3(baudrate[13]), .O(n59026));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_966.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_967 (.I0(byte_counter[0]), .I1(n50789), 
            .I2(data[6]), .I3(baudrate[14]), .O(n59024));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_967.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_968 (.I0(byte_counter[0]), .I1(n50789), 
            .I2(data[7]), .I3(baudrate[15]), .O(n59020));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_968.LUT_INIT = 16'hfb40;
    SB_LUT4 i13709_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[0]), 
            .I3(baudrate[16]), .O(n31654));   // verilog/eeprom.v(68[25:39])
    defparam i13709_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13708_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[1]), 
            .I3(baudrate[17]), .O(n31653));   // verilog/eeprom.v(68[25:39])
    defparam i13708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13707_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[2]), 
            .I3(baudrate[18]), .O(n31652));   // verilog/eeprom.v(68[25:39])
    defparam i13707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13706_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[3]), 
            .I3(baudrate[19]), .O(n31651));   // verilog/eeprom.v(68[25:39])
    defparam i13706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13705_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[4]), 
            .I3(baudrate[20]), .O(n31650));   // verilog/eeprom.v(68[25:39])
    defparam i13705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13704_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[5]), 
            .I3(baudrate[21]), .O(n31649));   // verilog/eeprom.v(68[25:39])
    defparam i13704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13703_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[6]), 
            .I3(baudrate[22]), .O(n31648));   // verilog/eeprom.v(68[25:39])
    defparam i13703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13702_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50789), .I2(data[7]), 
            .I3(baudrate[23]), .O(n31647));   // verilog/eeprom.v(68[25:39])
    defparam i13702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i34532_2_lut_3_lut_4_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i34532_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    i2c_controller i2c (.GND_net(GND_net), .\state[3] (state_adj_4447[3]), 
            .\state[0] (\state[0] ), .n4(n4_adj_4441), .n64433(n64433), 
            .clk16MHz(clk16MHz), .scl_enable(scl_enable), .\state_7__N_4110[0] (\state_7__N_4110[0] ), 
            .VCC_net(VCC_net), .n41842(n41842), .sda_enable(sda_enable), 
            .n59552(n59552), .\saved_addr[0] (saved_addr[0]), .n32362(n32362), 
            .data({data}), .n32360(n32360), .n32356(n32356), .n32339(n32339), 
            .n32338(n32338), .n32337(n32337), .n32335(n32335), .n32065(n32065), 
            .n8(n8), .n6722(n6722), .scl(scl), .sda_out(sda_out), .enable_slow_N_4213(enable_slow_N_4213), 
            .\state_7__N_4126[3] (\state_7__N_4126[3] ), .enable(enable), 
            .n41430(n41430), .n6(n6), .n4_adj_1(n4), .n4_adj_2(n4_adj_3), 
            .n41590(n41590), .n10(n10), .n27672(n27672), .n27624(n27624)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (GND_net, \state[3] , \state[0] , n4, n64433, 
            clk16MHz, scl_enable, \state_7__N_4110[0] , VCC_net, n41842, 
            sda_enable, n59552, \saved_addr[0] , n32362, data, n32360, 
            n32356, n32339, n32338, n32337, n32335, n32065, n8, 
            n6722, scl, sda_out, enable_slow_N_4213, \state_7__N_4126[3] , 
            enable, n41430, n6, n4_adj_1, n4_adj_2, n41590, n10, 
            n27672, n27624) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output \state[3] ;
    output \state[0] ;
    output n4;
    output n64433;
    input clk16MHz;
    output scl_enable;
    output \state_7__N_4110[0] ;
    input VCC_net;
    output n41842;
    output sda_enable;
    input n59552;
    output \saved_addr[0] ;
    input n32362;
    output [7:0]data;
    input n32360;
    input n32356;
    input n32339;
    input n32338;
    input n32337;
    input n32335;
    input n32065;
    input n8;
    output n6722;
    output scl;
    output sda_out;
    output enable_slow_N_4213;
    input \state_7__N_4126[3] ;
    input enable;
    output n41430;
    output n6;
    output n4_adj_1;
    output n4_adj_2;
    output n41590;
    output n10;
    output n27672;
    output n27624;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n6715, n67753, i2c_clk_N_4199, scl_enable_N_4200, enable_slow_N_4212, 
        n29851;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n31165, n53511, n53510, n53509, n53508, n53507, n62552, 
        n29846, n59222, n62101, n29844, sda_out_adj_4430;
    wire [7:0]n119;
    
    wire n29896;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n31102, n10_c, n5, n62960, n41728, n41905, n62860, n62586, 
        n52810, n52809, n52808, n52807, n52806, n52805, n52804, 
        n11, n11_adj_4431, n11_adj_4432, n11_adj_4433, n4_adj_4434, 
        n4_adj_4435, n11_adj_4436, n29722, n9, n12, n61039, n28, 
        n70913, n60932;
    wire [1:0]n6791;
    
    wire n10_adj_4440;
    
    SB_LUT4 i49357_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(n6715), 
            .I3(GND_net), .O(n67753));
    defparam i49357_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n4));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45172_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(\state[0] ), 
            .I3(GND_net), .O(n64433));
    defparam i45172_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n29851), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFSR counter2_2058_2059__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 counter2_2058_2059_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n53511), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2058_2059_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n53510), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2058_2059_add_4_6 (.CI(n53510), .I0(GND_net), .I1(counter2[4]), 
            .CO(n53511));
    SB_LUT4 counter2_2058_2059_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n53509), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2058_2059_add_4_5 (.CI(n53509), .I0(GND_net), .I1(counter2[3]), 
            .CO(n53510));
    SB_LUT4 counter2_2058_2059_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n53508), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2058_2059_add_4_4 (.CI(n53508), .I0(GND_net), .I1(counter2[2]), 
            .CO(n53509));
    SB_LUT4 counter2_2058_2059_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n53507), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2058_2059_add_4_3 (.CI(n53507), .I0(GND_net), .I1(counter2[1]), 
            .CO(n53508));
    SB_LUT4 counter2_2058_2059_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2058_2059_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2058_2059_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n53507));
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[3] ), .I2(state[2]), 
            .I3(state[1]), .O(n41842));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n29846), 
            .D(n62552), .S(n59222));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4430), .C(i2c_clk), .E(n29844), 
            .D(n62101), .S(n59222));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n29896), .D(n119[0]), 
            .S(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n31165));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n31165), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4199));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n59552));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n32362));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n32360));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n32356));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n32339));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n32338));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n32337));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n32335));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n32065));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n29896), .D(n119[1]), 
            .S(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n29896), .D(n119[2]), 
            .S(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n29896), .D(n119[3]), 
            .R(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n29896), .D(n119[4]), 
            .R(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n29896), .D(n119[5]), 
            .R(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n29896), .D(n119[6]), 
            .R(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n29896), .D(n119[7]), 
            .R(n31102));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n6722), .D(n5), 
            .S(n62960));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(state[2]), .C(i2c_clk), .E(n6722), .D(n41728), 
            .S(n41905));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6722), .D(n62860), 
            .S(n62586));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2058_2059__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2058_2059__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2058_2059__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2058_2059__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2058_2059__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n31165));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n52810), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n52809), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n52809), .I0(counter[6]), .I1(VCC_net), 
            .CO(n52810));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n52808), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n52808), .I0(counter[5]), .I1(VCC_net), 
            .CO(n52809));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n52807), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n52807), .I0(counter[4]), .I1(VCC_net), 
            .CO(n52808));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n52806), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n52806), .I0(counter[3]), .I1(VCC_net), 
            .CO(n52807));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n52805), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n52805), .I0(counter[2]), .I1(VCC_net), 
            .CO(n52806));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n52804), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n52804), .I0(counter[1]), .I1(VCC_net), 
            .CO(n52805));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n52804));
    SB_LUT4 i23628_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i23628_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2558_2_lut (.I0(sda_out_adj_4430), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2558_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51661_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(state[1]), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i51661_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(state[1]), .O(n11));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i23690_4_lut_4_lut_4_lut (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(state[1]), .O(scl_enable_N_4200));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i23690_4_lut_4_lut_4_lut.LUT_INIT = 16'hffea;
    SB_LUT4 i51654_2_lut (.I0(enable_slow_N_4213), .I1(\state_7__N_4110[0] ), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));
    defparam i51654_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(state[1]), .O(n11_adj_4431));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i2_3_lut_4_lut_adj_944 (.I0(\state[3] ), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[2]), .O(n62552));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_944.LUT_INIT = 16'h1110;
    SB_LUT4 equal_1564_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(state[2]), .I3(\state[3] ), .O(n11_adj_4432));
    defparam equal_1564_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4433), .I2(n11_adj_4432), 
            .I3(enable), .O(n4_adj_4434));
    defparam i1_4_lut.LUT_INIT = 16'h2a2f;
    SB_LUT4 i51808_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_4433), 
            .I2(GND_net), .I3(GND_net), .O(n41728));
    defparam i51808_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_945 (.I0(n6722), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4435));
    defparam i1_2_lut_adj_945.LUT_INIT = 16'hdddd;
    SB_LUT4 i51779_4_lut (.I0(\state[3] ), .I1(n4_adj_4435), .I2(\state[0] ), 
            .I3(state[1]), .O(n62960));
    defparam i51779_4_lut.LUT_INIT = 16'h0130;
    SB_LUT4 i1_4_lut_adj_946 (.I0(n11_adj_4436), .I1(n11_adj_4433), .I2(\state_7__N_4126[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h5755;
    SB_LUT4 i51667_4_lut (.I0(n29722), .I1(n6715), .I2(n11), .I3(n41430), 
            .O(n6722));
    defparam i51667_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i2_2_lut_4_lut_4_lut (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(state[1]), .O(n6));
    defparam i2_2_lut_4_lut_4_lut.LUT_INIT = 16'hfebf;
    SB_LUT4 i23619_2_lut_3_lut (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n41430));
    defparam i23619_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 state_7__I_0_145_i11_2_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[2]), .I3(\state[3] ), .O(n11_adj_4436));   // verilog/i2c_controller.v(161[5:14])
    defparam state_7__I_0_145_i11_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i51775_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), .I2(state[1]), 
            .I3(n6722), .O(n62586));
    defparam i51775_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(enable_slow_N_4213), .I2(\state_7__N_4110[0] ), 
            .I3(GND_net), .O(n29851));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i23744_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n41590));
    defparam i23744_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), .I2(state[2]), 
            .I3(\state[3] ), .O(n29722));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(\state[3] ), .I3(state[2]), .O(n11_adj_4433));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6715));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n29896), .I1(state[2]), .I2(\state[0] ), .I3(GND_net), 
            .O(n31102));
    defparam i3_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i41816_3_lut (.I0(state[2]), .I1(\state_7__N_4126[3] ), .I2(state[1]), 
            .I3(GND_net), .O(n61039));
    defparam i41816_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_947 (.I0(\state[3] ), .I1(n67753), .I2(n61039), 
            .I3(\state[0] ), .O(n29896));
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h0544;
    SB_LUT4 i1_4_lut_adj_948 (.I0(\state[3] ), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[2]), .O(n28));
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h5110;
    SB_LUT4 i51643_2_lut (.I0(\state[3] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n70913));
    defparam i51643_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n11_adj_4432), .I1(n70913), .I2(n28), 
            .I3(n60932), .O(n29844));
    defparam i1_4_lut_adj_949.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1832_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6791[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1832_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 state_7__I_0_144_i10_2_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4440));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i41711_2_lut (.I0(\state[0] ), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n60932));
    defparam i41711_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n11_adj_4432), .I1(n60932), .I2(\state[3] ), 
            .I3(state[1]), .O(n59222));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n11_adj_4432), .I1(state[1]), .I2(\state[3] ), 
            .I3(n60932), .O(n29846));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_2_lut_3_lut_adj_951 (.I0(n9), .I1(n10_adj_4440), .I2(counter[0]), 
            .I3(GND_net), .O(n27672));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_951.LUT_INIT = 16'hfefe;
    SB_LUT4 i51777_3_lut_4_lut (.I0(n9), .I1(n10_adj_4440), .I2(n11_adj_4431), 
            .I3(n6722), .O(n41905));   // verilog/i2c_controller.v(151[5:14])
    defparam i51777_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut_adj_952 (.I0(n9), .I1(n10_adj_4440), .I2(counter[0]), 
            .I3(GND_net), .O(n27624));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_952.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_953 (.I0(state[2]), .I1(\state[3] ), .I2(n4_adj_4434), 
            .I3(n9), .O(n62860));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_953.LUT_INIT = 16'hf0f4;
    SB_LUT4 i2_3_lut_4_lut_adj_954 (.I0(state[2]), .I1(\state[3] ), .I2(n6791[1]), 
            .I3(state[1]), .O(n62101));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_954.LUT_INIT = 16'h1000;
    
endmodule
