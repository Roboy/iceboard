// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Oct  4 23:07:54 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    input PIN_3 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    output PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    output PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    output PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    output PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    output PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    inout PIN_20 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    inout PIN_21 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    inout PIN_22 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire GND_net, VCC_net, CLK_c, LED_c, PIN_6_c_0, PIN_7_c_1, PIN_8_c_2, 
        PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, PIN_13_c, PIN_14_c, PIN_18_c_1, 
        PIN_19_c_0, PIN_23_c_1, PIN_24_c_0;
    wire [23:0]color;   // verilog/TinyFPGA_B.v(42[14:19])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(73[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(74[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(75[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(76[22:30])
    
    wire n47465, n47461;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(77[22:24])
    
    wire n48126, n48613;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(78[22:24])
    
    wire n48383;
    wire [23:0]Kd;   // verilog/TinyFPGA_B.v(79[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(80[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(81[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(82[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(83[22:30])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(84[22:34])
    
    wire hall1, hall2, hall3;
    wire [23:0]pwm;   // verilog/TinyFPGA_B.v(92[10:13])
    wire [31:0]motor_state;   // verilog/TinyFPGA_B.v(152[22:33])
    wire [23:0]color_23__N_1;
    
    wire PIN_13_N_50;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_51;
    wire [24:0]displacement_23__N_118;
    wire [23:0]displacement_23__N_25;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n34858;
    wire [3:0]state_3__N_248;
    
    wire n35151, n47451, n35150, n34857, n18466, n18470, n18469, 
        n18468, n18467, n34856, n18459, n48879, n35149, n35148, 
        n34855, n16688, n15, n35147, n34854, n25, n35146, n35145, 
        n47440, n35144, n34853, n18464, n18463, n18462, n2666, 
        n2665, n2664, n47434, n18458, n40180, n34852, n2663, n2662, 
        n2593, n2594, n2661, n2660, n2659, n2658, n2657, n2656, 
        n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, 
        n2647, n2646, n2645, n2644, n2643, n2616, n2615, n2614, 
        n2613, n2612, n2611, n2610, n2609, n2608, n34851, n35143, 
        n35142, n47430, n34850, n34849, n35141, n23171, n44294, 
        n47428, n18460, n534, n533, n532, n531, n530, n529, 
        n528, n527, n526, n525, n524, n523, n522, n521, n520, 
        n519, n518, n517, n516, n515, n514, n513, n512, n511, 
        n510, n17863, n17862, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n47396;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n16683, n16680, n16675, n47394, n34848;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n48397, n34847, n16672, n47392, n123, n34846, n40968, 
        n34845, n16678, n44276, n48404, n2607, n2606, n2605, n2604, 
        n2603, n2596, n2595, n35118, n35117, n35116, n35115, n35114, 
        n35113, n35112, n35111, n35110, n740, n35109, n35108, 
        n35107, n35106, n35105, n35104, n35103, n35102, n35101, 
        n35100, n35099, n35098, n35097, n18457, n18456, n35096, 
        n35095, n35094, n48433, n16669, n16666, n35093, n35092, 
        n35091, n118, n35090, n49070, n6, n35089, n35088, n16663, 
        n50704, n35087, n43362, n20911, n29, n35086, n35085, n35084, 
        n35083, n16660, n35082, n35081, n35080, n16657, n16654, 
        n16651, n16648, n16645, n16642, n16639, n16636, n18369, 
        n18368, n16633, n16630, n2484, n2602, n2601, n2600, n24, 
        n23, n22, n21, n20, n19, n18, n17, n2244, n2857, n18367, 
        n18366, n18365, n18364, n18363, n18362, n16627, n16624, 
        n48188, n8, n35056, n6_adj_4559, n4, n35055, n15_adj_4560, 
        n35054, n35053, n35052, Kp_23__N_679, n35051, n35050, n35049, 
        n35048, n35047, n2, n35046, n35045, n35044, n35043, n35042, 
        n35041, n48247, n35040, n35039, n35038, n49067, n35037, 
        n35036, n35035, n35034, n35033, n35032, n41336, n19921, 
        n35031, n35030, n35029, n35028, n35027, n16621, n48461, 
        n4_adj_4561, n2_adj_4562, n16617, n40184, n40176, n40172, 
        n40208, n40204, n40200, n40196, n18329, n18328, n18327, 
        n18326, n18325, n18324, n18323, n18322, n18305, n18304, 
        n18303, n40192, n18302, n18301, n18300, n18299, n18298, 
        n18266, n18265, n18264, n18263, n18262, n18261, n18260, 
        n18259, n18258, n18257, n18256, n18255, n18254, n18253, 
        n18252, n18251, n18250, n18249, n18248, n18247, n18246, 
        n18245, n18244, n18243, n18242, n18241, n18240, n18239, 
        n18238, n18237, n18236, n18235, n18234, n18233, n18232, 
        n18231, n18230, n18229, n18228, n18227, n18226, n18225, 
        n18224, n18223, n18222, n18221, n18220, n18219, n18218, 
        n18217, n18216, n18215, n18214, n18213, n18212, n18211, 
        n18210, n18209, n18208, n18207, n18206, n18205, n18204, 
        n18203, n18202, n18201, n18200, n18199, n18198, n18197, 
        n18196, n18195, n18194, n18193, n18192, n18191, n18190, 
        n18189, n18188, n18187, n18186, n18185, n18184, n18183, 
        n18182, n18181, n18180, n18179, n18178, n18177, n18176, 
        n18175, n18174, n18173, n18172, n18171, n18170, n18169, 
        n18168, n18167, n18166, n18165, n18164, n18163, n18162, 
        n18161, n18160, n18159, n18158, n18157, n18156, n18155, 
        n18154, n18153, n18152, n18151, n18150, n18149, n18148, 
        n18147, n18146, n18145, n18144, n18143, n18142, n18141, 
        n18140, n18139, n18135, n18134, n18133, n18132, n18131, 
        n18130, n18129, n18128, n18127, n18126, n18125, n18124, 
        n18123, n18122, n18121, n18120, n18119, n18118, n18117, 
        n18116, n18115, n18114, n18113, n18112, n18111, n18110, 
        n18109, n18108, n18107, n18106, n18105, n18104, n18103, 
        n18102, n18101, n18100, n18099, n18098, n18097, n18096, 
        n18095, n393, n392, n369, n18094, n249, n248, n18093, 
        n18092, n18091, n18090, n18089, n18088, n18087, n18086, 
        n18085, n18084, n18083, n18082, n18081, n18080, n18079, 
        n18078, n18077, n18076, n18075, n18074, n18073, n18072, 
        n18071, n18070, n224, n41857, n16614, n48212, n18433, 
        n49062, n18432, n29_adj_4563, n18431, n18430, n16, n18069, 
        n4469, n4468, n4467, n4466, n4465, n4464, n4463, n4462, 
        n4461, n4460, n4459, n4458, n4457, n4456, n4455, n4454, 
        n4453, n4452, n4451, n4450, n4449, n4448, n4447, n4446, 
        n18429, n18068;
    wire [31:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(30[23:26])
    wire [31:0]\PID_CONTROLLER.err_prev ;   // verilog/motorControl.v(31[23:31])
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    wire [8:0]pwm_count;   // verilog/motorControl.v(62[13:22])
    
    wire n40188, n18451, n18450, n18449, n18448, n18447, n48482, 
        n25_adj_4564, n24_adj_4565, n23_adj_4566, n22_adj_4567, n21_adj_4568, 
        n20_adj_4569, n19_adj_4570, n18_adj_4571, n17_adj_4572, n16_adj_4573, 
        n15_adj_4574, n14, n13, n12, n11, n10, n9, n8_adj_4575, 
        n7, n6_adj_4576, n4497, n41348;
    wire [31:0]pwm_23__N_3310;
    
    wire pwm_23__N_3307, n387, n401, n403, n407, n410, n414, n416, 
        n448, n449, n450, n451, n453, n455, n456, n457, n459, 
        n460, n462, n463, n464, n466, n48977, n468, n469, n470, 
        n471, n15_adj_4577, n14_adj_4578, n13_adj_4579, n12_adj_4580, 
        n11_adj_4581, n10_adj_4582, n9_adj_4583, n8_adj_4584, n7_adj_4585, 
        n6_adj_4586, n5, n4_adj_4587, n3, n99, n98, n97, n96, 
        n2599, n2598, GATES_5__N_3405, n4694;
    wire [5:0]GATES_5__N_3398;
    
    wire n853, n855, n856, n857, n859, n860, n861, n862, n863, 
        n864, n865, n866, n867, n868, n869, n870, n871, n872, 
        n873, n874, n875, n2597, n35002, quadA_debounced, quadB_debounced, 
        count_enable, n48478, n4_adj_4588, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, 
        n81, n80, n79, n78, n77, n75, n74, n73, n72, n71, 
        n35001, quadA_debounced_adj_4589, quadB_debounced_adj_4590, count_enable_adj_4591, 
        n16572, n4_adj_4592, n70, n69, n68, n67, n66, n65, n64, 
        n63, n62, n61, n60, n59, n58, n57, n56, n55, n54, 
        n53, n18428, n2677, n48658, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n35000, n221, n225, n226;
    wire [2:0]r_SM_Main_2__N_3032;
    
    wire n18067, n18066, n18065, n18064, n18063, n18062, n18061, 
        n18060, n18059;
    wire [2:0]r_SM_Main_adj_5024;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_5025;   // verilog/uart_tx.v(32[16:29])
    
    wire n34999, n18058, n18057, n18056, n18055, n18054, n18053, 
        n18052, n18051, n18050;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    wire [1:0]reg_B_adj_5037;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n34998, n34997, n34996, n34995, n48236, n34994, n35333, 
        n35332, n34993, n35331, n35330, n34992, n35329, n34991, 
        n35328, n35327, n34990, n34989, n35326, n35325, n4_adj_4596, 
        n35324, n34988, n35323, n3_adj_4597, n35322, n48940, n35321, 
        n35320, n35319, n35318, n35317, n35316, n3_adj_4598, n15_adj_4599, 
        n35315, n558, n35314, n35313, n35312, n648, n649, n671, 
        n672, n35311, n40168, n35310, n37696, n35309, n783, n784, 
        n785, n806, n807, n35308, n40156, n41851, n914, n915, 
        n916, n917, n918, n938, n939, n35307, n35306, n35305, 
        n14276, n1043, n1044, n1045, n1046, n1047, n1048, n1067, 
        n1068, n35304, n35303, n35302, n40144, n1169, n1170, n1171, 
        n1172, n1173, n1174, n1175, n35301, n34962, n1193, n1194, 
        n35300, n34961, n35299, n35298, n35297, n35296, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n35295, 
        n40164, n1316, n1317, n48877, n40160, n6481, n6482, n6483, 
        n6484, n6485, n40136, n34960, n41862, n35294, n34959, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n1436, n1437, n34958, n35293, n8_adj_4600, n50009, 
        n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
        n1537, n1538, n1553, n1554, n6443, n6442, n6441, n6440, 
        n6439, n6438, n40152, n6502, n6503, n6504, n6505, n6506, 
        n6507, n6508, n6509, n6510, n6511, n6512, n40148, n42459, 
        n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
        n1651, n1652, n1653, n6452, n6451, n6450, n6449, n6448, 
        n6447, n1667, n1668, n47079, n35292, n34957, n35291, n16687, 
        n34956, n41848, n1754, n1755, n1756, n1757, n1758, n1759, 
        n1760, n1761, n1762, n1763, n1764, n1765, n35290, n1778, 
        n1779, n34955, n35289, n35288, n40120, n1862, n1863, n1864, 
        n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
        n1873, n1874, n35287, n6462, n6461, n6460, n6459, n6458, 
        n1886, n1887, n35286, n6456, n6455, n40140, n6546, n6547, 
        n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
        n6556, n6557, n6558, n6559, n6471, n6472, n6473, n1967, 
        n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
        n1976, n1977, n1978, n1979, n1980, n6470, n6469, n6468, 
        n6467, n6466, n35285, n1991, n1992, n18446, n34954, n6572, 
        n6573, n6574, n6575, n6576, n6577, n6578, n2069, n2070, 
        n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
        n2079, n2080, n2081, n2082, n2083, n2093, n2094, n47071, 
        n6597, n40116, n35284, n34953, n2168, n2169, n2170, n2171, 
        n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
        n2180, n2181, n2182, n2183, n2192, n2193, n6608, n6609, 
        n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, 
        n6638, n6660, n6477, n6478, n6479, n6480, n35283, n2264, 
        n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
        n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
        n6476, n40132, n2288, n2289, n34952, n6620, n6621, n6622, 
        n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, 
        n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6497, 
        n6498, n35282, n40128, n2357, n2358, n2359, n2360, n2361, 
        n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
        n2370, n2371, n2372, n2373, n2374, n6496, n6495, n6494, 
        n6493, n6492, n6491, n2381, n2382, n6489, n6488, n6641, 
        n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, 
        n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
        n6658, n6659, n2447, n2448, n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
        n2461, n2462, n2463, n2464, n2465, n2471, n2472, n6665, 
        n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
        n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
        n6682, n6683, n10_adj_4601, n16550, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n2558, n2559, n47061, n6692, n6693, n6694, n6695, 
        n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
        n6704, n6705, n6706, n6707, n2618, n2619, n2620, n2621, 
        n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
        n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
        n2638, n2642, n2643_adj_4602, n35281, n6714, n6715, n6716, 
        n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, 
        n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, 
        n47055, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
        n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
        n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2723, 
        n2724, n35280, n2777, n2798, n2799, n2801, n2802, n18049, 
        n18048, n18047, n18046, n18045, n18044, n18043, n18042, 
        n18041, n35279, n18040, n18039, n18038, n35278, n18034, 
        n18033, n18032, n40124, n5_adj_4603, n6527, n6526, n6525, 
        n6524, n6523, n6522, n6521, n6520, n6519, n6518, n6517, 
        n6516, n6515, n48399, n6560, n6543, n6542, n6541, n6540, 
        n6539, n6538, n6537, n6536, n6535, n6534, n6533, n6532, 
        n6531, n47041, n18442, n4_adj_4604, n35277, n41860, n35276, 
        n35275, n35274, n35273, n35272, n35271, n35270, n6571, 
        n6570, n35269, n6569, n6568, n6567, n35268, n6566, n6565, 
        n6564, n6563, n35267, n6596, n6595, n6594, n6593, n35266, 
        n6592, n6591, n6590, n6589, n6588, n6587, n6586, n6585, 
        n6584, n6583, n6582, n6581, n6607, n6606, n6605, n6604, 
        n6603, n6602, n6601, n35265, n35264, n35263, n35262, n35261, 
        n35260, n35259, n35258, n47021, n35257, n35256, n6664, 
        n6663, n6691, n6690, n6689, n6688, n6687, n6686, n6713, 
        n6712, n35255, n35254, n48445, n35253, n35252, n9_adj_4605, 
        n13_adj_4606, n21_adj_4607, n27, n35, n39, n48403, n9_adj_4608, 
        n13_adj_4609, n22_adj_4610, n9_adj_4611, n13_adj_4612, n21_adj_4613, 
        n27_adj_4614, n44088, n9_adj_4615, n13_adj_4616, n21_adj_4617, 
        n27_adj_4618, n35_adj_4619, n39_adj_4620, n48474, n35251, 
        n4_adj_4621, n6_adj_4622, n8_adj_4623, n9_adj_4624, n11_adj_4625, 
        n13_adj_4626, n15_adj_4627, n18013, n18012, n35250, n18011, 
        n18010, n18009, n18008, n18007, n18006, n18005, n18004, 
        n18003, n18002, n18001, n18000, n17999, n17998, n17997, 
        n17996, n17995, n17994, n17993, n35249, n17992, n17991, 
        n41916, n17984, n17983, n17980, n17977, n17974, n17973, 
        n17971, n17970, n17969, n17967, n17966, n17965, n47019, 
        n17963, n17962, n17961, n35248, n17960, n17959, n17958, 
        n17955, n35247, n38230, n6711, n6710, n48158, n18427, 
        n47000, n5_adj_4628, n7_adj_4629, n18701, n4_adj_4630, n6_adj_4631, 
        n8_adj_4632, n9_adj_4633, n16_adj_4634, n18698, n18697, n18696, 
        n18695, n18694, n18693, n18692, n18691, n18690, n18689, 
        n46995, n18688, n18687, n18686, n18685, n18684, n18683, 
        n18682, n18681, n18680, n18679, n18678, n18677, n18676, 
        n18675, n18674, n18673, n18672, n46992, n48160, n18671, 
        n18670, n40242, n17897, n17896, n17895, n17894, n17893, 
        n17892, n17891, n46980, n17890, n18669, n18668, n18667, 
        n18666, n18665, n18664, n18663, n18662, n18661, n18660, 
        n18659, n18658, n18657, n18656, n18655, n18654, n18653, 
        n18652, n18651, n18650, n18649, n18648, n18647, n18646, 
        n18645, n18644, n18643, n18642, n18641, n18639, n18637, 
        n2_adj_4635, n3_adj_4636, n4_adj_4637, n5_adj_4638, n6_adj_4639, 
        n7_adj_4640, n8_adj_4641, n9_adj_4642, n10_adj_4643, n11_adj_4644, 
        n12_adj_4645, n13_adj_4646, n14_adj_4647, n15_adj_4648, n16_adj_4649, 
        n17_adj_4650, n18_adj_4651, n19_adj_4652, n20_adj_4653, n21_adj_4654, 
        n22_adj_4655, n23_adj_4656, n24_adj_4657, n25_adj_4658, n2_adj_4659, 
        n3_adj_4660, n4_adj_4661, n5_adj_4662, n6_adj_4663, n7_adj_4664, 
        n8_adj_4665, n9_adj_4666, n10_adj_4667, n11_adj_4668, n12_adj_4669, 
        n13_adj_4670, n14_adj_4671, n15_adj_4672, n16_adj_4673, n17_adj_4674, 
        n18_adj_4675, n19_adj_4676, n20_adj_4677, n21_adj_4678, n22_adj_4679, 
        n23_adj_4680, n24_adj_4681, n25_adj_4682, n17283, n46, n18636, 
        n18635, n18633, n18632, n18630, n18629, n18628, n18626, 
        n18624, n18623, n18622, n18618, n44, n48480, n18616, n18615, 
        n18614, n18613, n18612, n18611, n18610, n18609, n18608, 
        n18607, n18606, n18605, n18604, n18603, n18602, n18601, 
        n18600, n18599, n18598, n42, n18597, n18596, n46971, n18595, 
        n18594, n18593, n18587, n18583, n42216, n40, n42_adj_4683, 
        n44_adj_4684, n45, n18575, n18574, n18567, n38, n40_adj_4685, 
        n42_adj_4686, n43, n48489, n48744, n18555, n18552, n18550, 
        n18548, n18547, n36, n38_adj_4687, n40_adj_4688, n41, n18545, 
        n18544, n18542, n18541, n18539, n18538, n18536, n18535, 
        n18533, n18532, n34, n36_adj_4689, n38_adj_4690, n39_adj_4691, 
        n41_adj_4692, n43_adj_4693, n44_adj_4694, n45_adj_4695, n48232, 
        n18531, n18530, n18529, n18528, n18527, n18526, n18525, 
        n18524, n18523, n18522, n18521, n18520, n18519, n18518, 
        n32, n34_adj_4696, n37, n39_adj_4697, n41_adj_4698, n48660, 
        n43_adj_4699, n18517, n18516, n18515, n18514, n18513, n18512, 
        n18511, n18510, n18509, n18507, n46965, n30, n31, n32_adj_4700, 
        n33, n34_adj_4701, n35_adj_4702, n37_adj_4703, n39_adj_4704, 
        n48656, n41_adj_4705, n42_adj_4706, n43_adj_4707, n45_adj_4708, 
        n48841, n18497, n18495, n18494, n18493, n28, n29_adj_4709, 
        n30_adj_4710, n31_adj_4711, n32_adj_4712, n33_adj_4713, n35_adj_4714, 
        n37_adj_4715, n48654, n39_adj_4716, n40_adj_4717, n41_adj_4718, 
        n43_adj_4719, n48652, n18492, n18491, n18490, n18489, n18488, 
        n18487, n18486, n18485, n18484, n18483, n18482, n26, n27_adj_4720, 
        n28_adj_4721, n29_adj_4722, n30_adj_4723, n31_adj_4724, n33_adj_4725, 
        n35_adj_4726, n48650, n37_adj_4727, n38_adj_4728, n39_adj_4729, 
        n41_adj_4730, n48932, n18481, n18480, n18479, n18478, n18477, 
        n18476, n18475, n18474, n18473, n18472, n18471, n24_adj_4731, 
        n25_adj_4732, n26_adj_4733, n27_adj_4734, n28_adj_4735, n29_adj_4736, 
        n30_adj_4737, n31_adj_4738, n32_adj_4739, n33_adj_4740, n35_adj_4741, 
        n36_adj_4742, n37_adj_4743, n39_adj_4744, n41_adj_4745, n48506, 
        n43_adj_4746, n44_adj_4747, n45_adj_4748, n48508, n17887, 
        n6457, n22_adj_4749, n23_adj_4750, n24_adj_4751, n25_adj_4752, 
        n26_adj_4753, n27_adj_4754, n28_adj_4755, n29_adj_4756, n30_adj_4757, 
        n31_adj_4758, n33_adj_4759, n34_adj_4760, n35_adj_4761, n37_adj_4762, 
        n39_adj_4763, n41_adj_4764, n42_adj_4765, n43_adj_4766, n48642, 
        n20_adj_4767, n21_adj_4768, n22_adj_4769, n23_adj_4770, n24_adj_4771, 
        n25_adj_4772, n26_adj_4773, n27_adj_4774, n28_adj_4775, n29_adj_4776, 
        n31_adj_4777, n32_adj_4778, n33_adj_4779, n35_adj_4780, n37_adj_4781, 
        n39_adj_4782, n41_adj_4783, n48636, n49016, n17707, n18_adj_4784, 
        n19_adj_4785, n20_adj_4786, n21_adj_4787, n22_adj_4788, n23_adj_4789, 
        n24_adj_4790, n25_adj_4791, n26_adj_4792, n27_adj_4793, n29_adj_4794, 
        n30_adj_4795, n31_adj_4796, n33_adj_4797, n35_adj_4798, n37_adj_4799, 
        n48942, n39_adj_4800, n41_adj_4801, n42_adj_4802, n43_adj_4803, 
        n45_adj_4804, n48244, n16_adj_4805, n17_adj_4806, n18_adj_4807, 
        n19_adj_4808, n20_adj_4809, n21_adj_4810, n22_adj_4811, n23_adj_4812, 
        n25_adj_4813, n27_adj_4814, n28_adj_4815, n29_adj_4816, n31_adj_4817, 
        n33_adj_4818, n35_adj_4819, n36_adj_4820, n37_adj_4821, n39_adj_4822, 
        n40_adj_4823, n41_adj_4824, n43_adj_4825, n48880, n14_adj_4826, 
        n16_adj_4827, n17_adj_4828, n18_adj_4829, n19_adj_4830, n20_adj_4831, 
        n21_adj_4832, n22_adj_4833, n23_adj_4834, n25_adj_4835, n26_adj_4836, 
        n27_adj_4837, n29_adj_4838, n31_adj_4839, n33_adj_4840, n48770, 
        n35_adj_4841, n37_adj_4842, n48628, n39_adj_4843, n40_adj_4844, 
        n41_adj_4845, n43_adj_4846, n45_adj_4847, n48772, n6490, n12_adj_4848, 
        n14_adj_4849, n15_adj_4850, n16_adj_4851, n17_adj_4852, n18_adj_4853, 
        n19_adj_4854, n20_adj_4855, n21_adj_4856, n23_adj_4857, n24_adj_4858, 
        n25_adj_4859, n27_adj_4860, n29_adj_4861, n31_adj_4862, n48948, 
        n33_adj_4863, n35_adj_4864, n48624, n37_adj_4865, n38_adj_4866, 
        n39_adj_4867, n41_adj_4868, n43_adj_4869, n48622, n10_adj_4870, 
        n12_adj_4871, n13_adj_4872, n14_adj_4873, n15_adj_4874, n16_adj_4875, 
        n17_adj_4876, n18_adj_4877, n19_adj_4878, n21_adj_4879, n22_adj_4880, 
        n23_adj_4881, n25_adj_4882, n27_adj_4883, n29_adj_4884, n48950, 
        n31_adj_4885, n33_adj_4886, n48618, n35_adj_4887, n36_adj_4888, 
        n37_adj_4889, n39_adj_4890, n41_adj_4891, n48952, n49071, 
        n14246, n8_adj_4892, n10_adj_4893, n11_adj_4894, n12_adj_4895, 
        n13_adj_4896, n14_adj_4897, n15_adj_4898, n16_adj_4899, n17_adj_4900, 
        n19_adj_4901, n20_adj_4902, n21_adj_4903, n23_adj_4904, n25_adj_4905, 
        n48614, n27_adj_4906, n29_adj_4907, n31_adj_4908, n48612, 
        n33_adj_4909, n34_adj_4910, n35_adj_4911, n37_adj_4912, n39_adj_4913, 
        n48554, n48556, n48558, n6_adj_4914, n8_adj_4915, n9_adj_4916, 
        n10_adj_4917, n11_adj_4918, n12_adj_4919, n13_adj_4920, n14_adj_4921, 
        n15_adj_4922, n17_adj_4923, n19_adj_4924, n21_adj_4925, n23_adj_4926, 
        n48387, n25_adj_4927, n27_adj_4928, n29_adj_4929, n31_adj_4930, 
        n32_adj_4931, n33_adj_4932, n35_adj_4933, n37_adj_4934, n48878, 
        n48861, n4_adj_4935, n6_adj_4936, n7_adj_4937, n8_adj_4938, 
        n9_adj_4939, n10_adj_4940, n11_adj_4941, n12_adj_4942, n13_adj_4943, 
        n15_adj_4944, n16_adj_4945, n17_adj_4946, n19_adj_4947, n21_adj_4948, 
        n48668, n23_adj_4949, n24_adj_4950, n25_adj_4951, n27_adj_4952, 
        n29_adj_4953, n30_adj_4954, n31_adj_4955, n33_adj_4956, n35_adj_4957, 
        n37_adj_4958, n39_adj_4959, n41_adj_4960, n43_adj_4961, n45_adj_4962, 
        n48910, n46951, n46949, n46947, n46913, n17849, n46908, 
        n46896, n46892, n46889, n46887, n46881, n48190, n16563, 
        n17665, n46877, n46871, n17657, n46865, n43079, n41444, 
        n48245, n17872, n17632, n46849, n46847, n46845, n35225, 
        n46841, n46839, n41446, n17869, n17866, n35224, n46830, 
        n35223, n48216, n46828, n88_adj_4963, n17802, n35222, n48230, 
        n35221, n35220, n46812, n46808, n46806, n43352, n46804, 
        n46802, n48234, n46800, n48242, n35219, n47844, n46781, 
        n46779, n42577, n35218, n35217, n46775, n46772, n35216, 
        n35215, n46759, n35214, n46743, n35213, n35212, n46741, 
        n6_adj_4964, n35211, n4_adj_4965, n49075, n49074, n49053, 
        n49045, n49043, n49042, n49065, n49020, n49044, n46739, 
        n46737, n46735, n46733, n49017, n46723, n17574, n18393, 
        n18392, n18426, n49005, n49046, n35_adj_4966, n30_adj_4967, 
        n49052, n28_adj_4968, n46719, n26_adj_4969, n25_adj_4970, 
        n17503, n49048, n48924, n48978, n49014, n48955, n48949, 
        n48947, n48945, n48943, n48941, n48937, n48935, n48933, 
        n46705, n48908, n48876, n46703, n48869, n48862, n46701, 
        n48858, n48842, n48838, n48836, n48834, n48938, n48830, 
        n48828, n48826, n48824, n48822, n35210, n46697, n40240, 
        n40236, n40232, n40228, n40224, n40220, n40216, n40212, 
        n18455, n18391, n18454, n48776, n18453, n18390, n3_adj_4971, 
        n2_adj_4972, n18389, n18452, n48774, n48946, n35209, n48769, 
        n48944, n19_adj_4973, n48765, n48757, n48936, n35208, n6446, 
        n48934, n35207, n48748, n48745, n6465, n48930, n6501, 
        n37_adj_4974, n35206, n35205, n28_adj_4975, n6530, n6600, 
        n48857, n48701, n48859, n35204, n48695, n48690, n48669, 
        n48667, n48666, n48661, n48659, n35203, n48657, n48655, 
        n48651, n46660, n48637, n35202, n46659, n48633, n48629, 
        n35201, n35200, n35199, n48625, n46658, n46657, n35198, 
        n48560, n46656, n46655, n48551, n46654, n48549, n46653, 
        n48545, n46652, n35197, n48539, n35196, n18445, n18388, 
        n18444, n18387, n35195, n18443, n18386, n48535, n48632, 
        n35194, n35588, n35587, n46651, n35586, n35585, n48530, 
        n35584, n35583, n35582, n35581, n46650, n35580, n35579, 
        n35578, n35577, n35576, n35575, n35574, n35573, n35572, 
        n35571, n46649, n35570, n35569, n35568, n35567, n35566, 
        n35565, n35564, n35563, n35562, n35561, n35560, n35559, 
        n35558, n35557, n35556, n35555, n35554, n46648, n46647, 
        n48501, n35193, n25520, n35553, n35552, n35192, n35551, 
        n46646, n35550, n35191, n48497, n48495, n46645, n35190, 
        n23694, n35189, n35188, n35549, n46644, n35548, n35187, 
        n35547, n35546, n35545, n35544, n35186, n35543, n35185, 
        n35184, n35183, n35182, n46643, n35181, n35180, n35179, 
        n35178, n35177, n46642, n35176, n48122, n35175, n35174, 
        n46641, n48118, n35173, n35172, n35171, n46640, n35170, 
        n35169, n48096, n48092, n35168, n35167, n46639, n2_adj_4976, 
        n46638, n46637, n46636, n46635, n35166, n42079, n25329, 
        n46634, n16566, n46633, n46632, n35165, n35164, n35163, 
        n35162, n34867, n42066, n35161, n46631, n44245, n34866, 
        n46630, n34865, n35160, n34864, n37561, n35159, n35158, 
        n34863, n35157, n35156, n34862, n34861, n35155, n42125, 
        n37512, n35154, n35153, n34860, n34859, n27708, n43056, 
        n16432, n35152, n46629, n46628, n48619, n47866, n47841, 
        n47835, n47833, n47821, n47819, n48395, n47796, n43650, 
        n47779, n47765, n47738, n48413, n49780, n48449, n41781, 
        n16_adj_4977, n47649, n15_adj_4978, n42357, n14_adj_4979, 
        n13_adj_4980, n49063, n42429, n43448, n42330, n42342, n47581, 
        n5_adj_4981, n41074, n5_adj_4982, n47561, n48396, n48388, 
        n41130, n42140, n41150, n48386, n48926, n48361, n47478, 
        n47511, n47492, n47499, n47503, n47531, n41224, n47533, 
        n47474, n42219, n42432, n48615, n46549, n46548, n48956, 
        n41442, n48960, n42610, n42696, n48684, n42503, n42501, 
        n42499, n4_adj_4983, n48680, n48875, n5_adj_4984, n8_adj_4985, 
        n7_adj_4986, n48385;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF color_i1 (.Q(color[0]), .C(clk32MHz), .D(color_23__N_1[0]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_IO hall1_input (.PACKAGE_PIN(PIN_20), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall2_input (.PACKAGE_PIN(PIN_21), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_22), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3140_12 (.CI(n35320), .I0(n49780), .I1(n1886), .CO(n35321));
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3140_11_lut (.I0(n1992), .I1(n49780), .I2(n1991), .I3(n35319), 
            .O(displacement_23__N_118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_11_lut.LUT_INIT = 16'h8BB8;
    neopixel nx (.clk32MHz(clk32MHz), .timer({timer}), .bit_ctr({bit_ctr}), 
            .VCC_net(VCC_net), .n40240(n40240), .n40236(n40236), .n40232(n40232), 
            .n40228(n40228), .n40224(n40224), .n40220(n40220), .n46646(n46646), 
            .GND_net(GND_net), .n41781(n41781), .n40216(n40216), .n40212(n40212), 
            .n40208(n40208), .n40204(n40204), .n40200(n40200), .n40196(n40196), 
            .n46634(n46634), .n40192(n40192), .n40188(n40188), .n40184(n40184), 
            .n40180(n40180), .n40176(n40176), .n40172(n40172), .n40168(n40168), 
            .n40164(n40164), .n40160(n40160), .n40156(n40156), .n40152(n40152), 
            .n40148(n40148), .n40144(n40144), .n40140(n40140), .n40136(n40136), 
            .n40132(n40132), .n18698(n18698), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n18697(n18697), .n18696(n18696), .n18695(n18695), .n18694(n18694), 
            .n18693(n18693), .n18692(n18692), .n18691(n18691), .n18690(n18690), 
            .n18689(n18689), .n18688(n18688), .n18687(n18687), .n18686(n18686), 
            .n18685(n18685), .n18684(n18684), .n18683(n18683), .n18682(n18682), 
            .n18681(n18681), .n18680(n18680), .n18679(n18679), .n18678(n18678), 
            .n18677(n18677), .n18676(n18676), .n18675(n18675), .n18674(n18674), 
            .n18673(n18673), .n18672(n18672), .n18671(n18671), .n18670(n18670), 
            .n18669(n18669), .n18668(n18668), .n40242(n40242), .start(start), 
            .n40116(n40116), .n18552(n18552), .\state[1] (state[1]), .n40120(n40120), 
            .n40124(n40124), .n40128(n40128), .n46645(n46645), .\state[0] (state[0]), 
            .n46644(n46644), .n46633(n46633), .n46643(n46643), .n35(n35_adj_4966), 
            .n46642(n46642), .n29(n29), .\state_3__N_248[1] (state_3__N_248[1]), 
            .n16572(n16572), .n20911(n20911), .n43079(n43079), .n46632(n46632), 
            .n46641(n46641), .n46631(n46631), .n46640(n46640), .n46639(n46639), 
            .n46630(n46630), .n17665(n17665), .n17802(n17802), .n46629(n46629), 
            .n46659(n46659), .n46658(n46658), .n46638(n46638), .n46657(n46657), 
            .n46656(n46656), .n46655(n46655), .n46654(n46654), .n46637(n46637), 
            .n46653(n46653), .n17984(n17984), .n46652(n46652), .n46651(n46651), 
            .n46636(n46636), .n46650(n46650), .n46628(n46628), .PIN_14_c(PIN_14_c), 
            .n46649(n46649), .n46635(n46635), .n46648(n46648), .n46647(n46647), 
            .n17574(n17574), .\color[2] (color[2]), .\color[3] (color[3]), 
            .n4(n4_adj_4983), .n43650(n43650), .\color[1] (color[1]), 
            .\color[0] (color[0]), .\color[6] (color[6]), .\color[7] (color[7]), 
            .\color[5] (color[5]), .\color[4] (color[4]), .\color[10] (color[10]), 
            .\color[11] (color[11]), .\color[9] (color[9]), .\color[8] (color[8]), 
            .\color[18] (color[18]), .\color[19] (color[19]), .\color[17] (color[17]), 
            .\color[16] (color[16]), .\color[14] (color[14]), .\color[15] (color[15]), 
            .\color[13] (color[13]), .\color[12] (color[12])) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(52[12] 58[4])
    SB_CARRY add_3140_11 (.CI(n35319), .I0(n49780), .I1(n1991), .CO(n35320));
    SB_LUT4 add_3140_10_lut (.I0(n2094), .I1(n49780), .I2(n2093), .I3(n35318), 
            .O(displacement_23__N_118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_10 (.CI(n35318), .I0(n49780), .I1(n2093), .CO(n35319));
    SB_LUT4 add_3140_9_lut (.I0(n2193), .I1(n49780), .I2(n2192), .I3(n35317), 
            .O(displacement_23__N_118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_9 (.CI(n35317), .I0(n49780), .I1(n2192), .CO(n35318));
    SB_LUT4 add_3140_8_lut (.I0(n2289), .I1(n49780), .I2(n2288), .I3(n35316), 
            .O(displacement_23__N_118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_8 (.CI(n35316), .I0(n49780), .I1(n2288), .CO(n35317));
    SB_IO PIN_10_pad (.PACKAGE_PIN(PIN_10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_10_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_10_pad.PIN_TYPE = 6'b011001;
    defparam PIN_10_pad.PULLUP = 1'b0;
    defparam PIN_10_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3140_7_lut (.I0(n2382), .I1(n49780), .I2(n2381), .I3(n35315), 
            .O(displacement_23__N_118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_7 (.CI(n35315), .I0(n49780), .I1(n2381), .CO(n35316));
    SB_LUT4 add_3140_6_lut (.I0(n2472), .I1(n49780), .I2(n2471), .I3(n35314), 
            .O(displacement_23__N_118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_6 (.CI(n35314), .I0(n49780), .I1(n2471), .CO(n35315));
    SB_LUT4 add_3140_5_lut (.I0(n2559), .I1(n49780), .I2(n2558), .I3(n35313), 
            .O(displacement_23__N_118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_5 (.CI(n35313), .I0(n49780), .I1(n2558), .CO(n35314));
    SB_LUT4 add_3140_4_lut (.I0(n2643_adj_4602), .I1(n49780), .I2(n2642), 
            .I3(n35312), .O(displacement_23__N_118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7_2_lut (.I0(deadband[19]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(32[23:29])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3140_4 (.CI(n35312), .I0(n49780), .I1(n2642), .CO(n35313));
    SB_LUT4 i5_2_lut (.I0(deadband[17]), .I1(\PID_CONTROLLER.result [17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(32[23:29])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3140_3_lut (.I0(n2724), .I1(n49780), .I2(n2723), .I3(n35311), 
            .O(displacement_23__N_118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_3 (.CI(n35311), .I0(n49780), .I1(n2723), .CO(n35312));
    SB_LUT4 add_3140_2_lut (.I0(n2802), .I1(n49780), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_2 (.CI(VCC_net), .I0(n49780), .I1(n2801), .CO(n35311));
    SB_LUT4 add_3139_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n35310), 
            .O(n6710)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3139_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n35309), 
            .O(n6711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_24 (.CI(n35309), .I0(n2700), .I1(n79), .CO(n35310));
    SB_LUT4 add_3139_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n35308), 
            .O(n6712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_23 (.CI(n35308), .I0(n2701), .I1(n80), .CO(n35309));
    SB_LUT4 add_3139_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n35307), 
            .O(n6713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_22 (.CI(n35307), .I0(n2702), .I1(n81), .CO(n35308));
    SB_LUT4 add_3139_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n35306), 
            .O(n6714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_21 (.CI(n35306), .I0(n2703), .I1(n82), .CO(n35307));
    SB_LUT4 add_3139_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n35305), 
            .O(n6715)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_20 (.CI(n35305), .I0(n2704), .I1(n83), .CO(n35306));
    SB_LUT4 add_3139_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n35304), 
            .O(n6716)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_19 (.CI(n35304), .I0(n2705), .I1(n84), .CO(n35305));
    SB_LUT4 add_3139_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n35303), 
            .O(n6717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_18 (.CI(n35303), .I0(n2706), .I1(n85), .CO(n35304));
    SB_LUT4 add_3139_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n35302), 
            .O(n6718)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_17 (.CI(n35302), .I0(n2707), .I1(n86), .CO(n35303));
    SB_LUT4 add_3139_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n35301), 
            .O(n6719)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_16 (.CI(n35301), .I0(n2708), .I1(n87), .CO(n35302));
    SB_LUT4 add_3139_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n35300), 
            .O(n6720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_15 (.CI(n35300), .I0(n2709), .I1(n88), .CO(n35301));
    SB_LUT4 add_3139_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n35299), 
            .O(n6721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_14 (.CI(n35299), .I0(n2710), .I1(n89), .CO(n35300));
    SB_LUT4 add_3139_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n35298), 
            .O(n6722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_13 (.CI(n35298), .I0(n2711), .I1(n90), .CO(n35299));
    SB_LUT4 add_3139_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n35297), 
            .O(n6723)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_12 (.CI(n35297), .I0(n2712), .I1(n91), .CO(n35298));
    SB_LUT4 add_3139_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n35296), 
            .O(n6724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_11 (.CI(n35296), .I0(n2713), .I1(n92), .CO(n35297));
    SB_LUT4 add_3139_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n35295), 
            .O(n6725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_10 (.CI(n35295), .I0(n2714), .I1(n93), .CO(n35296));
    SB_LUT4 add_3139_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n35294), 
            .O(n6726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_9 (.CI(n35294), .I0(n2715), .I1(n94), .CO(n35295));
    SB_LUT4 add_3139_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n35293), 
            .O(n6727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_8 (.CI(n35293), .I0(n2716), .I1(n95), .CO(n35294));
    SB_LUT4 add_3139_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n35292), 
            .O(n6728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_7 (.CI(n35292), .I0(n2717), .I1(n96), .CO(n35293));
    SB_LUT4 add_3139_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n35291), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_6 (.CI(n35291), .I0(n2718), .I1(n97), .CO(n35292));
    SB_LUT4 add_3139_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n35290), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_5 (.CI(n35290), .I0(n2719), .I1(n98), .CO(n35291));
    SB_LUT4 add_3139_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n35289), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_4 (.CI(n35289), .I0(n2720), .I1(n99), .CO(n35290));
    SB_LUT4 add_3139_3_lut (.I0(GND_net), .I1(n531), .I2(n558), .I3(n35288), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3139_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3139_3 (.CI(n35288), .I0(n531), .I1(n558), .CO(n35289));
    SB_CARRY add_3139_2 (.CI(VCC_net), .I0(n532), .I1(VCC_net), .CO(n35288));
    SB_LUT4 add_3138_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n35287), 
            .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n35286), 
            .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_22 (.CI(n35286), .I0(n2619), .I1(n80), .CO(n35287));
    SB_LUT4 add_3138_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n35285), 
            .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_21 (.CI(n35285), .I0(n2620), .I1(n81), .CO(n35286));
    SB_LUT4 add_3138_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n35284), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_20 (.CI(n35284), .I0(n2621), .I1(n82), .CO(n35285));
    SB_LUT4 add_3138_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n35283), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_19 (.CI(n35283), .I0(n2622), .I1(n83), .CO(n35284));
    SB_LUT4 add_3138_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n35282), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_18 (.CI(n35282), .I0(n2623), .I1(n84), .CO(n35283));
    SB_LUT4 add_3123_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n34962), 
            .O(n6446)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n35281), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3123_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n34961), 
            .O(n6447)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_17 (.CI(n35281), .I0(n2624), .I1(n85), .CO(n35282));
    SB_CARRY add_3123_7 (.CI(n34961), .I0(n1044), .I1(n95), .CO(n34962));
    SB_LUT4 add_3138_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n35280), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_16 (.CI(n35280), .I0(n2625), .I1(n86), .CO(n35281));
    SB_LUT4 add_3123_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n34960), 
            .O(n6448)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_2_lut (.I0(deadband[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4606));   // verilog/motorControl.v(32[23:29])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3138_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n35279), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_15 (.CI(n35279), .I0(n2626), .I1(n87), .CO(n35280));
    SB_CARRY add_3123_6 (.CI(n34960), .I0(n1045), .I1(n96), .CO(n34961));
    SB_LUT4 add_3138_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n35278), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_14 (.CI(n35278), .I0(n2627), .I1(n88), .CO(n35279));
    SB_LUT4 add_3123_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n34959), 
            .O(n6449)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n35277), 
            .O(n6696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_13 (.CI(n35277), .I0(n2628), .I1(n89), .CO(n35278));
    SB_CARRY add_3123_5 (.CI(n34959), .I0(n1046), .I1(n97), .CO(n34960));
    SB_LUT4 i13_2_lut (.I0(deadband[13]), .I1(\PID_CONTROLLER.result [13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(32[23:29])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3138_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n35276), 
            .O(n6697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_12 (.CI(n35276), .I0(n2629), .I1(n90), .CO(n35277));
    SB_LUT4 add_3123_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n34958), 
            .O(n6450)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n35275), 
            .O(n6698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_11 (.CI(n35275), .I0(n2630), .I1(n91), .CO(n35276));
    SB_CARRY add_3123_4 (.CI(n34958), .I0(n1047), .I1(n98), .CO(n34959));
    SB_LUT4 add_3138_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n35274), 
            .O(n6699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_10 (.CI(n35274), .I0(n2631), .I1(n92), .CO(n35275));
    SB_LUT4 add_3123_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n34957), 
            .O(n6451)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n35273), 
            .O(n6700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_9 (.CI(n35273), .I0(n2632), .I1(n93), .CO(n35274));
    SB_CARRY add_3123_3 (.CI(n34957), .I0(n1048), .I1(n99), .CO(n34958));
    SB_LUT4 add_3138_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n35272), 
            .O(n6701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3123_2_lut (.I0(GND_net), .I1(n515), .I2(n558), .I3(VCC_net), 
            .O(n6452)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3123_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_8 (.CI(n35272), .I0(n2633), .I1(n94), .CO(n35273));
    SB_CARRY add_3123_2 (.CI(VCC_net), .I0(n515), .I1(n558), .CO(n34957));
    SB_LUT4 add_3138_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n35271), 
            .O(n6702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3122_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n34956), 
            .O(n6438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_7 (.CI(n35271), .I0(n2634), .I1(n95), .CO(n35272));
    SB_LUT4 add_3122_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n34955), 
            .O(n6439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n35270), 
            .O(n6703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3122_6 (.CI(n34955), .I0(n915), .I1(n96), .CO(n34956));
    SB_CARRY add_3138_6 (.CI(n35270), .I0(n2635), .I1(n96), .CO(n35271));
    SB_LUT4 add_3122_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n34954), 
            .O(n6440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n35269), 
            .O(n6704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3122_5 (.CI(n34954), .I0(n916), .I1(n97), .CO(n34955));
    SB_CARRY add_3138_5 (.CI(n35269), .I0(n2636), .I1(n97), .CO(n35270));
    SB_LUT4 add_3122_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n34953), 
            .O(n6441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3138_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n35268), 
            .O(n6705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3122_4 (.CI(n34953), .I0(n917), .I1(n98), .CO(n34954));
    SB_CARRY add_3138_4 (.CI(n35268), .I0(n2637), .I1(n98), .CO(n35269));
    SB_LUT4 i22_2_lut (.I0(deadband[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4605));   // verilog/motorControl.v(32[23:29])
    defparam i22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3122_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n34952), 
            .O(n6442)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3122_3 (.CI(n34952), .I0(n918), .I1(n99), .CO(n34953));
    SB_LUT4 add_3138_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n35267), 
            .O(n6706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3122_2_lut (.I0(GND_net), .I1(n514), .I2(n558), .I3(VCC_net), 
            .O(n6443)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3122_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_3 (.CI(n35267), .I0(n2638), .I1(n99), .CO(n35268));
    SB_CARRY add_3122_2 (.CI(VCC_net), .I0(n514), .I1(n558), .CO(n34952));
    SB_LUT4 i24_2_lut (.I0(PWMLimit[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4611));   // verilog/motorControl.v(32[23:29])
    defparam i24_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3138_2_lut (.I0(GND_net), .I1(n530), .I2(n558), .I3(VCC_net), 
            .O(n6707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3138_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3138_2 (.CI(VCC_net), .I0(n530), .I1(n558), .CO(n35267));
    SB_LUT4 i18_2_lut (.I0(PWMLimit[10]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4613));   // verilog/motorControl.v(32[23:29])
    defparam i18_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11_2_lut (.I0(PWMLimit[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4612));   // verilog/motorControl.v(32[23:29])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_2_lut_adj_1568 (.I0(PWMLimit[13]), .I1(\PID_CONTROLLER.result [13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4614));   // verilog/motorControl.v(32[23:29])
    defparam i14_2_lut_adj_1568.LUT_INIT = 16'h6666;
    SB_LUT4 add_3137_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n35266), 
            .O(n6663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3137_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n35265), 
            .O(n6664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1417_i18_4_lut (.I0(n525), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4784));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40733_3_lut (.I0(n18_adj_4784), .I1(n87), .I2(n41_adj_4801), 
            .I3(GND_net), .O(n48636));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40733_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3137_21 (.CI(n35265), .I0(n2535), .I1(n81), .CO(n35266));
    SB_LUT4 i15_2_lut (.I0(deadband[10]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4607));   // verilog/motorControl.v(32[23:29])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_LessThan_1417_i30_3_lut (.I0(n22_adj_4788), .I1(n91), 
            .I2(n33_adj_4797), .I3(GND_net), .O(n30_adj_4795));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3137_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n35264), 
            .O(n6665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40734_3_lut (.I0(n48636), .I1(n86), .I2(n43_adj_4803), .I3(GND_net), 
            .O(n48637));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40734_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3137_20 (.CI(n35264), .I0(n2536), .I1(n82), .CO(n35265));
    SB_LUT4 i41037_4_lut (.I0(n30_adj_4795), .I1(n20_adj_4786), .I2(n33_adj_4797), 
            .I3(n46737), .O(n48940));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41037_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3137_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n35263), 
            .O(n6666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_19 (.CI(n35263), .I0(n2537), .I1(n83), .CO(n35264));
    SB_IO PIN_18_pad (.PACKAGE_PIN(PIN_18), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_18_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_18_pad.PIN_TYPE = 6'b000001;
    defparam PIN_18_pad.PULLUP = 1'b0;
    defparam PIN_18_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3137_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n35262), 
            .O(n6667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_18 (.CI(n35262), .I0(n2538), .I1(n84), .CO(n35263));
    SB_LUT4 add_3137_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n35261), 
            .O(n6668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_17 (.CI(n35261), .I0(n2539), .I1(n85), .CO(n35262));
    SB_LUT4 add_3137_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n35260), 
            .O(n6669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_16 (.CI(n35260), .I0(n2540), .I1(n86), .CO(n35261));
    SB_LUT4 add_3137_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n35259), 
            .O(n6670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_15 (.CI(n35259), .I0(n2541), .I1(n87), .CO(n35260));
    SB_LUT4 i41038_3_lut (.I0(n48940), .I1(n90), .I2(n35_adj_4798), .I3(GND_net), 
            .O(n48941));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41038_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3137_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n35258), 
            .O(n6671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_14 (.CI(n35258), .I0(n2542), .I1(n88), .CO(n35259));
    SB_LUT4 add_3137_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n35257), 
            .O(n6672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_13 (.CI(n35257), .I0(n2543), .I1(n89), .CO(n35258));
    SB_LUT4 add_3137_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n35256), 
            .O(n6673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17624_3_lut (.I0(pwm_23__N_3310[10]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(n29_adj_4563), .I3(GND_net), .O(n22_adj_4610));   // verilog/motorControl.v(32[23:29])
    defparam i17624_3_lut.LUT_INIT = 16'hb2b2;
    SB_CARRY add_3137_12 (.CI(n35256), .I0(n2544), .I1(n90), .CO(n35257));
    SB_LUT4 add_3137_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n35255), 
            .O(n6674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_11 (.CI(n35255), .I0(n2545), .I1(n91), .CO(n35256));
    SB_LUT4 add_3137_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n35254), 
            .O(n6675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_10 (.CI(n35254), .I0(n2546), .I1(n92), .CO(n35255));
    SB_LUT4 add_3137_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n35253), 
            .O(n6676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_9 (.CI(n35253), .I0(n2547), .I1(n93), .CO(n35254));
    SB_LUT4 add_3137_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n35252), 
            .O(n6677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_8 (.CI(n35252), .I0(n2548), .I1(n94), .CO(n35253));
    SB_LUT4 add_3137_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n35251), 
            .O(n6678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_7 (.CI(n35251), .I0(n2549), .I1(n95), .CO(n35252));
    SB_LUT4 add_3137_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n35250), 
            .O(n6679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_25[1]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_LUT4 i40927_3_lut (.I0(n48941), .I1(n89), .I2(n37_adj_4799), .I3(GND_net), 
            .O(n48830));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40927_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_25[0]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_CARRY add_3137_6 (.CI(n35250), .I0(n2550), .I1(n96), .CO(n35251));
    SB_LUT4 add_3137_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n35249), 
            .O(n6680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_5 (.CI(n35249), .I0(n2551), .I1(n97), .CO(n35250));
    SB_LUT4 add_3137_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n35248), 
            .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_4 (.CI(n35248), .I0(n2552), .I1(n98), .CO(n35249));
    SB_LUT4 add_3137_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n35247), 
            .O(n6682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_3 (.CI(n35247), .I0(n2553), .I1(n99), .CO(n35248));
    SB_LUT4 add_3137_2_lut (.I0(GND_net), .I1(n529), .I2(n558), .I3(VCC_net), 
            .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3137_2 (.CI(VCC_net), .I0(n529), .I1(n558), .CO(n35247));
    SB_LUT4 i39630_4_lut (.I0(n43_adj_4803), .I1(n41_adj_4801), .I2(n39_adj_4800), 
            .I3(n48399), .O(n47533));
    defparam i39630_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40339_4_lut (.I0(n42_adj_4802), .I1(n26_adj_4792), .I2(n45_adj_4804), 
            .I3(n47531), .O(n48242));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40339_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40862_3_lut (.I0(n48830), .I1(n88), .I2(n39_adj_4800), .I3(GND_net), 
            .O(n48765));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40862_3_lut.LUT_INIT = 16'h3a3a;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3136_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n35225), 
            .O(n6641)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3136_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n35224), 
            .O(n6642)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_20 (.CI(n35224), .I0(n2448), .I1(n82), .CO(n35225));
    SB_LUT4 add_3136_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n35223), 
            .O(n6643)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_19 (.CI(n35223), .I0(n2449), .I1(n83), .CO(n35224));
    SB_LUT4 add_3136_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n35222), 
            .O(n6644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_18 (.CI(n35222), .I0(n2450), .I1(n84), .CO(n35223));
    SB_LUT4 add_3136_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n35221), 
            .O(n6645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_17 (.CI(n35221), .I0(n2451), .I1(n85), .CO(n35222));
    SB_LUT4 add_3136_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n35220), 
            .O(n6646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_16 (.CI(n35220), .I0(n2452), .I1(n86), .CO(n35221));
    SB_LUT4 add_3136_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n35219), 
            .O(n6647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_15 (.CI(n35219), .I0(n2453), .I1(n87), .CO(n35220));
    SB_LUT4 add_3136_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n35218), 
            .O(n6648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_14 (.CI(n35218), .I0(n2454), .I1(n88), .CO(n35219));
    SB_LUT4 add_3136_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n35217), 
            .O(n6649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_13 (.CI(n35217), .I0(n2455), .I1(n89), .CO(n35218));
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_14_pad (.PACKAGE_PIN(PIN_14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_14_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_14_pad.PIN_TYPE = 6'b011001;
    defparam PIN_14_pad.PULLUP = 1'b0;
    defparam PIN_14_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c_5)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_23_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b000001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3136_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n35216), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_12 (.CI(n35216), .I0(n2456), .I1(n90), .CO(n35217));
    SB_LUT4 add_3136_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n35215), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_11 (.CI(n35215), .I0(n2457), .I1(n91), .CO(n35216));
    SB_LUT4 add_3136_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n35214), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_10 (.CI(n35214), .I0(n2458), .I1(n92), .CO(n35215));
    SB_LUT4 add_3136_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n35213), 
            .O(n6653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_9 (.CI(n35213), .I0(n2459), .I1(n93), .CO(n35214));
    SB_LUT4 add_3136_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n35212), 
            .O(n6654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_8 (.CI(n35212), .I0(n2460), .I1(n94), .CO(n35213));
    SB_LUT4 add_3136_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n35211), 
            .O(n6655)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_7 (.CI(n35211), .I0(n2461), .I1(n95), .CO(n35212));
    SB_LUT4 add_3136_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n35210), 
            .O(n6656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_6 (.CI(n35210), .I0(n2462), .I1(n96), .CO(n35211));
    SB_LUT4 add_3136_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n35209), 
            .O(n6657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_5 (.CI(n35209), .I0(n2463), .I1(n97), .CO(n35210));
    SB_LUT4 add_3136_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n35208), 
            .O(n6658)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_4 (.CI(n35208), .I0(n2464), .I1(n98), .CO(n35209));
    SB_LUT4 add_3136_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n35207), 
            .O(n6659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_3 (.CI(n35207), .I0(n2465), .I1(n99), .CO(n35208));
    SB_LUT4 add_3136_2_lut (.I0(GND_net), .I1(n528), .I2(n558), .I3(VCC_net), 
            .O(n6660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3136_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3136_2 (.CI(VCC_net), .I0(n528), .I1(n558), .CO(n35207));
    SB_LUT4 add_3135_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n35206), 
            .O(n6620)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3135_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n35205), 
            .O(n6621)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_19 (.CI(n35205), .I0(n2358), .I1(n83), .CO(n35206));
    SB_LUT4 add_3135_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n35204), 
            .O(n6622)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_18 (.CI(n35204), .I0(n2359), .I1(n84), .CO(n35205));
    SB_LUT4 i40341_4_lut (.I0(n48765), .I1(n48242), .I2(n45_adj_4804), 
            .I3(n47533), .O(n48244));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40341_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3135_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n35203), 
            .O(n6623)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_17 (.CI(n35203), .I0(n2360), .I1(n85), .CO(n35204));
    SB_LUT4 i39628_4_lut (.I0(n43_adj_4803), .I1(n41_adj_4801), .I2(n29_adj_4794), 
            .I3(n46741), .O(n47531));
    defparam i39628_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_15_LessThan_1417_i26_3_lut (.I0(n24_adj_4790), .I1(n93), 
            .I2(n29_adj_4794), .I3(GND_net), .O(n26_adj_4792));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40622_3_lut (.I0(n48637), .I1(n85), .I2(n45_adj_4804), .I3(GND_net), 
            .O(n42_adj_4802));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40622_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3135_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n35202), 
            .O(n6624)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_16 (.CI(n35202), .I0(n2361), .I1(n86), .CO(n35203));
    SB_LUT4 add_3135_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n35201), 
            .O(n6625)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_15 (.CI(n35201), .I0(n2362), .I1(n87), .CO(n35202));
    SB_LUT4 add_3135_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n35200), 
            .O(n6626)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1137_i38_3_lut (.I0(n30_adj_4723), .I1(n91), 
            .I2(n41_adj_4730), .I3(GND_net), .O(n38_adj_4728));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3135_14 (.CI(n35200), .I0(n2363), .I1(n88), .CO(n35201));
    SB_LUT4 add_3135_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n35199), 
            .O(n6627)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_13 (.CI(n35199), .I0(n2364), .I1(n89), .CO(n35200));
    SB_LUT4 i13360_4_lut (.I0(pwm_23__N_3307), .I1(n448), .I2(PWMLimit[23]), 
            .I3(n387), .O(n18644));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13360_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 add_3135_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n35198), 
            .O(n6628)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13361_3_lut (.I0(setpoint[1]), .I1(n4447), .I2(n43448), .I3(GND_net), 
            .O(n18645));   // verilog/coms.v(126[12] 289[6])
    defparam i13361_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3135_12 (.CI(n35198), .I0(n2365), .I1(n90), .CO(n35199));
    SB_LUT4 add_3135_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n35197), 
            .O(n6629)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13362_3_lut (.I0(setpoint[2]), .I1(n4448), .I2(n43448), .I3(GND_net), 
            .O(n18646));   // verilog/coms.v(126[12] 289[6])
    defparam i13362_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3135_11 (.CI(n35197), .I0(n2366), .I1(n91), .CO(n35198));
    SB_LUT4 add_3135_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n35196), 
            .O(n6630)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_10 (.CI(n35196), .I0(n2367), .I1(n92), .CO(n35197));
    SB_LUT4 add_3135_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n35195), 
            .O(n6631)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13363_3_lut (.I0(setpoint[3]), .I1(n4449), .I2(n43448), .I3(GND_net), 
            .O(n18647));   // verilog/coms.v(126[12] 289[6])
    defparam i13363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13364_3_lut (.I0(setpoint[4]), .I1(n4450), .I2(n43448), .I3(GND_net), 
            .O(n18648));   // verilog/coms.v(126[12] 289[6])
    defparam i13364_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3135_9 (.CI(n35195), .I0(n2368), .I1(n93), .CO(n35196));
    SB_LUT4 i13365_3_lut (.I0(setpoint[5]), .I1(n4451), .I2(n43448), .I3(GND_net), 
            .O(n18649));   // verilog/coms.v(126[12] 289[6])
    defparam i13365_3_lut.LUT_INIT = 16'hacac;
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_9_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b011001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c_2)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3135_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n35194), 
            .O(n6632)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_8 (.CI(n35194), .I0(n2369), .I1(n94), .CO(n35195));
    SB_LUT4 i13366_3_lut (.I0(setpoint[6]), .I1(n4452), .I2(n43448), .I3(GND_net), 
            .O(n18650));   // verilog/coms.v(126[12] 289[6])
    defparam i13366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3135_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n35193), 
            .O(n6633)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13367_3_lut (.I0(setpoint[7]), .I1(n4453), .I2(n43448), .I3(GND_net), 
            .O(n18651));   // verilog/coms.v(126[12] 289[6])
    defparam i13367_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13368_3_lut (.I0(setpoint[8]), .I1(n4454), .I2(n43448), .I3(GND_net), 
            .O(n18652));   // verilog/coms.v(126[12] 289[6])
    defparam i13368_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3135_7 (.CI(n35193), .I0(n2370), .I1(n95), .CO(n35194));
    SB_LUT4 i13369_3_lut (.I0(setpoint[9]), .I1(n4455), .I2(n43448), .I3(GND_net), 
            .O(n18653));   // verilog/coms.v(126[12] 289[6])
    defparam i13369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3135_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n35192), 
            .O(n6634)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_6 (.CI(n35192), .I0(n2371), .I1(n96), .CO(n35193));
    SB_LUT4 add_3135_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n35191), 
            .O(n6635)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_5 (.CI(n35191), .I0(n2372), .I1(n97), .CO(n35192));
    SB_LUT4 add_3135_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n35190), 
            .O(n6636)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_4 (.CI(n35190), .I0(n2373), .I1(n98), .CO(n35191));
    SB_LUT4 i13370_3_lut (.I0(setpoint[10]), .I1(n4456), .I2(n43448), 
            .I3(GND_net), .O(n18654));   // verilog/coms.v(126[12] 289[6])
    defparam i13370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3135_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n35189), 
            .O(n6637)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_3 (.CI(n35189), .I0(n2374), .I1(n99), .CO(n35190));
    SB_LUT4 add_3135_2_lut (.I0(GND_net), .I1(n527), .I2(n558), .I3(VCC_net), 
            .O(n6638)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3135_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3135_2 (.CI(VCC_net), .I0(n527), .I1(n558), .CO(n35189));
    SB_LUT4 add_3134_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n35188), 
            .O(n6600)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3134_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n35187), 
            .O(n6601)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_18 (.CI(n35187), .I0(n2265), .I1(n84), .CO(n35188));
    SB_LUT4 add_3134_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n35186), 
            .O(n6602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13371_3_lut (.I0(setpoint[11]), .I1(n4457), .I2(n43448), 
            .I3(GND_net), .O(n18655));   // verilog/coms.v(126[12] 289[6])
    defparam i13371_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3134_17 (.CI(n35186), .I0(n2266), .I1(n85), .CO(n35187));
    SB_LUT4 i13372_3_lut (.I0(setpoint[12]), .I1(n4458), .I2(n43448), 
            .I3(GND_net), .O(n18656));   // verilog/coms.v(126[12] 289[6])
    defparam i13372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13373_3_lut (.I0(setpoint[13]), .I1(n4459), .I2(n43448), 
            .I3(GND_net), .O(n18657));   // verilog/coms.v(126[12] 289[6])
    defparam i13373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13374_3_lut (.I0(setpoint[14]), .I1(n4460), .I2(n43448), 
            .I3(GND_net), .O(n18658));   // verilog/coms.v(126[12] 289[6])
    defparam i13374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3134_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n35185), 
            .O(n6603)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_16 (.CI(n35185), .I0(n2267), .I1(n86), .CO(n35186));
    SB_LUT4 i13375_3_lut (.I0(setpoint[15]), .I1(n4461), .I2(n43448), 
            .I3(GND_net), .O(n18659));   // verilog/coms.v(126[12] 289[6])
    defparam i13375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3134_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n35184), 
            .O(n6604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13376_3_lut (.I0(setpoint[16]), .I1(n4462), .I2(n43448), 
            .I3(GND_net), .O(n18660));   // verilog/coms.v(126[12] 289[6])
    defparam i13376_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3134_15 (.CI(n35184), .I0(n2268), .I1(n87), .CO(n35185));
    SB_LUT4 add_3134_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n35183), 
            .O(n6605)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13377_3_lut (.I0(setpoint[17]), .I1(n4463), .I2(n43448), 
            .I3(GND_net), .O(n18661));   // verilog/coms.v(126[12] 289[6])
    defparam i13377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13378_3_lut (.I0(setpoint[18]), .I1(n4464), .I2(n43448), 
            .I3(GND_net), .O(n18662));   // verilog/coms.v(126[12] 289[6])
    defparam i13378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n48244), .I1(n16657), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_CARRY add_3134_14 (.CI(n35183), .I0(n2269), .I1(n88), .CO(n35184));
    SB_LUT4 add_3134_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n35182), 
            .O(n6606)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13379_3_lut (.I0(setpoint[19]), .I1(n4465), .I2(n43448), 
            .I3(GND_net), .O(n18663));   // verilog/coms.v(126[12] 289[6])
    defparam i13379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13380_3_lut (.I0(setpoint[20]), .I1(n4466), .I2(n43448), 
            .I3(GND_net), .O(n18664));   // verilog/coms.v(126[12] 289[6])
    defparam i13380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13165_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[7] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18449));   // verilog/coms.v(126[12] 289[6])
    defparam i13165_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3134_13 (.CI(n35182), .I0(n2270), .I1(n89), .CO(n35183));
    SB_LUT4 add_3134_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n35181), 
            .O(n6607)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_12 (.CI(n35181), .I0(n2271), .I1(n90), .CO(n35182));
    SB_LUT4 i13166_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[7] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18450));   // verilog/coms.v(126[12] 289[6])
    defparam i13166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13167_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[7] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18451));   // verilog/coms.v(126[12] 289[6])
    defparam i13167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17156_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[7] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18452));
    defparam i17156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13169_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[7] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18453));   // verilog/coms.v(126[12] 289[6])
    defparam i13169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17274_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[7] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18454));
    defparam i17274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13171_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[7] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18455));   // verilog/coms.v(126[12] 289[6])
    defparam i13171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13172_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[6] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18456));   // verilog/coms.v(126[12] 289[6])
    defparam i13172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4578), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1199_3_lut (.I0(n521), .I1(n6527), .I2(n1778), .I3(GND_net), 
            .O(n1874));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13381_3_lut (.I0(setpoint[21]), .I1(n4467), .I2(n43448), 
            .I3(GND_net), .O(n18665));   // verilog/coms.v(126[12] 289[6])
    defparam i13381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3134_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n35180), 
            .O(n6608)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_11 (.CI(n35180), .I0(n2272), .I1(n91), .CO(n35181));
    SB_LUT4 div_15_i1270_3_lut (.I0(n1874), .I1(n6542), .I2(n1886), .I3(GND_net), 
            .O(n1979));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13382_3_lut (.I0(setpoint[22]), .I1(n4468), .I2(n43448), 
            .I3(GND_net), .O(n18666));   // verilog/coms.v(126[12] 289[6])
    defparam i13382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3134_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n35179), 
            .O(n6609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_10 (.CI(n35179), .I0(n2273), .I1(n92), .CO(n35180));
    SB_LUT4 div_15_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n16672));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 add_3134_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n35178), 
            .O(n6610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_9 (.CI(n35178), .I0(n2274), .I1(n93), .CO(n35179));
    SB_LUT4 div_15_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(n81), .I1(n16666), .I2(GND_net), .I3(GND_net), 
            .O(n16663));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'hdddd;
    SB_LUT4 div_15_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1570 (.I0(n84), .I1(n16657), .I2(GND_net), .I3(GND_net), 
            .O(n16654));
    defparam i1_2_lut_adj_1570.LUT_INIT = 16'hdddd;
    SB_LUT4 div_15_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4783));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3134_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n35177), 
            .O(n6611)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_8 (.CI(n35177), .I0(n2275), .I1(n94), .CO(n35178));
    SB_LUT4 div_15_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4781));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4782));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4780));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3134_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n35176), 
            .O(n6612)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_7 (.CI(n35176), .I0(n2276), .I1(n95), .CO(n35177));
    SB_LUT4 add_3134_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n35175), 
            .O(n6613)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_6 (.CI(n35175), .I0(n2277), .I1(n96), .CO(n35176));
    SB_LUT4 add_3134_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n35174), 
            .O(n6614)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4582), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i891_3_lut (.I0(n517), .I1(n6473), .I2(n1316), .I3(GND_net), 
            .O(n1420));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i970_3_lut (.I0(n1420), .I1(n6484), .I2(n1436), .I3(GND_net), 
            .O(n1537));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1047_3_lut (.I0(n1537), .I1(n6496), .I2(n1553), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1122_3_lut (.I0(n1651), .I1(n6509), .I2(n1667), .I3(GND_net), 
            .O(n1762));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1195_3_lut (.I0(n1762), .I1(n6523), .I2(n1778), .I3(GND_net), 
            .O(n1870));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1266_3_lut (.I0(n1870), .I1(n6538), .I2(n1886), .I3(GND_net), 
            .O(n1975));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4581), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i971_3_lut (.I0(n518), .I1(n6485), .I2(n1436), .I3(GND_net), 
            .O(n1538));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1048_3_lut (.I0(n1538), .I1(n6497), .I2(n1553), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1123_3_lut (.I0(n1652), .I1(n6510), .I2(n1667), .I3(GND_net), 
            .O(n1763));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1196_3_lut (.I0(n1763), .I1(n6524), .I2(n1778), .I3(GND_net), 
            .O(n1871));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1196_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3134_5 (.CI(n35174), .I0(n2278), .I1(n97), .CO(n35175));
    SB_LUT4 add_3134_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n35173), 
            .O(n6615)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_4 (.CI(n35173), .I0(n2279), .I1(n98), .CO(n35174));
    SB_LUT4 add_3134_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n35172), 
            .O(n6616)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3134_3 (.CI(n35172), .I0(n2280), .I1(n99), .CO(n35173));
    SB_LUT4 div_15_i1267_3_lut (.I0(n1871), .I1(n6539), .I2(n1886), .I3(GND_net), 
            .O(n1976));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4776));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4777));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4779));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4770));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4772));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4774));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4768));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3134_2_lut (.I0(GND_net), .I1(n526), .I2(n558), .I3(VCC_net), 
            .O(n6617)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3134_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38879_4_lut (.I0(n27_adj_4774), .I1(n25_adj_4772), .I2(n23_adj_4770), 
            .I3(n21_adj_4768), .O(n46781));
    defparam i38879_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38873_4_lut (.I0(n33_adj_4779), .I1(n31_adj_4777), .I2(n29_adj_4776), 
            .I3(n46781), .O(n46775));
    defparam i38873_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1350_i20_4_lut (.I0(n524), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4767));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_1350_i28_3_lut (.I0(n26_adj_4773), .I1(n93), 
            .I2(n31_adj_4777), .I3(GND_net), .O(n28_adj_4775));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3134_2 (.CI(VCC_net), .I0(n526), .I1(n558), .CO(n35172));
    SB_LUT4 add_3133_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n35171), 
            .O(n6581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1350_i32_3_lut (.I0(n24_adj_4771), .I1(n91), 
            .I2(n35_adj_4780), .I3(GND_net), .O(n32_adj_4778));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41033_4_lut (.I0(n32_adj_4778), .I1(n22_adj_4769), .I2(n35_adj_4780), 
            .I3(n46772), .O(n48936));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41033_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3133_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n35170), 
            .O(n6582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_17 (.CI(n35170), .I0(n2169), .I1(n85), .CO(n35171));
    SB_LUT4 i41034_3_lut (.I0(n48936), .I1(n90), .I2(n37_adj_4781), .I3(GND_net), 
            .O(n48937));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41034_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40931_3_lut (.I0(n48937), .I1(n89), .I2(n39_adj_4782), .I3(GND_net), 
            .O(n48834));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40931_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40510_4_lut (.I0(n39_adj_4782), .I1(n37_adj_4781), .I2(n35_adj_4780), 
            .I3(n46775), .O(n48413));
    defparam i40510_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i41035_4_lut (.I0(n28_adj_4775), .I1(n20_adj_4767), .I2(n31_adj_4777), 
            .I3(n46779), .O(n48938));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41035_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40854_3_lut (.I0(n48834), .I1(n88), .I2(n41_adj_4783), .I3(GND_net), 
            .O(n48757));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40854_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41113_4_lut (.I0(n48757), .I1(n48938), .I2(n41_adj_4783), 
            .I3(n48413), .O(n49016));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41113_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41114_3_lut (.I0(n49016), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n49017));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41114_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i41052_3_lut (.I0(n49017), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n48955));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41052_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n48955), .I1(n16654), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'hceef;
    SB_LUT4 i13173_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[6] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18457));   // verilog/coms.v(126[12] 289[6])
    defparam i13173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17630_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[6] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18458));
    defparam i17630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13175_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[6] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18459));   // verilog/coms.v(126[12] 289[6])
    defparam i13175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13176_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[6] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18460));   // verilog/coms.v(126[12] 289[6])
    defparam i13176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13383_3_lut (.I0(setpoint[23]), .I1(n4469), .I2(n43448), 
            .I3(GND_net), .O(n18667));   // verilog/coms.v(126[12] 289[6])
    defparam i13383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n35169), 
            .O(n6583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13384_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18668));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13384_3_lut.LUT_INIT = 16'hacac;
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_7_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b011001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_15_i1258_3_lut (.I0(n1862), .I1(n6530), .I2(n1886), .I3(GND_net), 
            .O(n1967));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1259_3_lut (.I0(n1863), .I1(n6531), .I2(n1886), .I3(GND_net), 
            .O(n1968));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4580), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1049_3_lut (.I0(n519), .I1(n6498), .I2(n1553), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1124_3_lut (.I0(n1653), .I1(n6511), .I2(n1667), .I3(GND_net), 
            .O(n1764));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1197_3_lut (.I0(n1764), .I1(n6525), .I2(n1778), .I3(GND_net), 
            .O(n1872));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1268_3_lut (.I0(n1872), .I1(n6540), .I2(n1886), .I3(GND_net), 
            .O(n1977));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4754));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i549_4_lut (.I0(n784), .I1(n4), .I2(n806), .I3(n98), 
            .O(n916));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i549_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_i636_3_lut (.I0(n916), .I1(n6440), .I2(n938), .I3(GND_net), 
            .O(n1045));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i721_3_lut (.I0(n1045), .I1(n6448), .I2(n1067), .I3(GND_net), 
            .O(n1171));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i804_3_lut (.I0(n1171), .I1(n6457), .I2(n1193), .I3(GND_net), 
            .O(n1294));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13385_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18669));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13385_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3133_16 (.CI(n35169), .I0(n2170), .I1(n86), .CO(n35170));
    SB_LUT4 div_15_i885_3_lut (.I0(n1294), .I1(n6467), .I2(n1316), .I3(GND_net), 
            .O(n1414));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i964_3_lut (.I0(n1414), .I1(n6478), .I2(n1436), .I3(GND_net), 
            .O(n1531));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13386_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18670));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1041_3_lut (.I0(n1531), .I1(n6490), .I2(n1553), .I3(GND_net), 
            .O(n1645));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1116_3_lut (.I0(n1645), .I1(n6503), .I2(n1667), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1189_3_lut (.I0(n1756), .I1(n6517), .I2(n1778), .I3(GND_net), 
            .O(n1864));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n35168), 
            .O(n6584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_15 (.CI(n35168), .I0(n2171), .I1(n87), .CO(n35169));
    SB_LUT4 add_3133_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n35167), 
            .O(n6585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_14 (.CI(n35167), .I0(n2172), .I1(n88), .CO(n35168));
    SB_LUT4 add_3133_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n35166), 
            .O(n6586)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1260_3_lut (.I0(n1864), .I1(n6532), .I2(n1886), .I3(GND_net), 
            .O(n1969));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4766));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i550_4_lut (.I0(n785), .I1(n2), .I2(n806), .I3(n99), 
            .O(n917));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i550_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_i637_3_lut (.I0(n917), .I1(n6441), .I2(n938), .I3(GND_net), 
            .O(n1046));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i722_3_lut (.I0(n1046), .I1(n6449), .I2(n1067), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i805_3_lut (.I0(n1172), .I1(n6458), .I2(n1193), .I3(GND_net), 
            .O(n1295));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i886_3_lut (.I0(n1295), .I1(n6468), .I2(n1316), .I3(GND_net), 
            .O(n1415));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13387_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18671));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13388_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18672));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13388_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3133_13 (.CI(n35166), .I0(n2173), .I1(n89), .CO(n35167));
    SB_LUT4 add_3133_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n35165), 
            .O(n6587)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_12 (.CI(n35165), .I0(n2174), .I1(n90), .CO(n35166));
    SB_LUT4 i13085_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n41857), .I3(GND_net), .O(n18369));   // verilog/coms.v(126[12] 289[6])
    defparam i13085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13389_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18673));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n35164), 
            .O(n6588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13390_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18674));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13390_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3133_11 (.CI(n35164), .I0(n2175), .I1(n91), .CO(n35165));
    SB_LUT4 add_3133_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n35163), 
            .O(n6589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_10 (.CI(n35163), .I0(n2176), .I1(n92), .CO(n35164));
    SB_LUT4 i13391_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18675));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13392_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18676));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n35162), 
            .O(n6590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i965_3_lut (.I0(n1415), .I1(n6479), .I2(n1436), .I3(GND_net), 
            .O(n1532));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i965_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3133_9 (.CI(n35162), .I0(n2177), .I1(n93), .CO(n35163));
    SB_LUT4 div_15_i1042_3_lut (.I0(n1532), .I1(n6491), .I2(n1553), .I3(GND_net), 
            .O(n1646));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1117_3_lut (.I0(n1646), .I1(n6504), .I2(n1667), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1190_3_lut (.I0(n1757), .I1(n6518), .I2(n1778), .I3(GND_net), 
            .O(n1865));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1261_3_lut (.I0(n1865), .I1(n6533), .I2(n1886), .I3(GND_net), 
            .O(n1970));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4764));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1262_3_lut (.I0(n1866), .I1(n6534), .I2(n1886), .I3(GND_net), 
            .O(n1971));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n35161), 
            .O(n6591)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4763));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3133_8 (.CI(n35161), .I0(n2178), .I1(n94), .CO(n35162));
    SB_LUT4 div_15_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4585), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n514));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i639_3_lut (.I0(n514), .I1(n6443), .I2(n938), .I3(GND_net), 
            .O(n1048));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i724_3_lut (.I0(n1048), .I1(n6451), .I2(n1067), .I3(GND_net), 
            .O(n1174));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i807_3_lut (.I0(n1174), .I1(n6460), .I2(n1193), .I3(GND_net), 
            .O(n1297));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n35160), 
            .O(n6592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_7 (.CI(n35160), .I0(n2179), .I1(n95), .CO(n35161));
    SB_LUT4 add_3133_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n35159), 
            .O(n6593)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13393_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18677));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i888_3_lut (.I0(n1297), .I1(n6470), .I2(n1316), .I3(GND_net), 
            .O(n1417));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13394_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18678));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_2_lut (.I0(n401), .I1(\PID_CONTROLLER.result [19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4620));   // verilog/motorControl.v(32[23:29])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3133_6 (.CI(n35159), .I0(n2180), .I1(n96), .CO(n35160));
    SB_LUT4 add_3133_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n35158), 
            .O(n6594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13395_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18679));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13395_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3133_5 (.CI(n35158), .I0(n2181), .I1(n97), .CO(n35159));
    SB_LUT4 add_3133_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n35157), 
            .O(n6595)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_4 (.CI(n35157), .I0(n2182), .I1(n98), .CO(n35158));
    SB_LUT4 div_15_i967_3_lut (.I0(n1417), .I1(n6481), .I2(n1436), .I3(GND_net), 
            .O(n1534));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1044_3_lut (.I0(n1534), .I1(n6493), .I2(n1553), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1119_3_lut (.I0(n1648), .I1(n6506), .I2(n1667), .I3(GND_net), 
            .O(n1759));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1192_3_lut (.I0(n1759), .I1(n6520), .I2(n1778), .I3(GND_net), 
            .O(n1867));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1263_3_lut (.I0(n1867), .I1(n6535), .I2(n1886), .I3(GND_net), 
            .O(n1972));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4762));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4579), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1125_3_lut (.I0(n520), .I1(n6512), .I2(n1667), .I3(GND_net), 
            .O(n1765));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1198_3_lut (.I0(n1765), .I1(n6526), .I2(n1778), .I3(GND_net), 
            .O(n1873));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1269_3_lut (.I0(n1873), .I1(n6541), .I2(n1886), .I3(GND_net), 
            .O(n1978));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4752));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1264_3_lut (.I0(n1868), .I1(n6536), .I2(n1886), .I3(GND_net), 
            .O(n1973));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13396_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18680));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3133_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n35156), 
            .O(n6596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_3 (.CI(n35156), .I0(n2183), .I1(n99), .CO(n35157));
    SB_LUT4 add_3133_2_lut (.I0(GND_net), .I1(n525), .I2(n558), .I3(VCC_net), 
            .O(n6597)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3133_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3133_2 (.CI(VCC_net), .I0(n525), .I1(n558), .CO(n35156));
    SB_LUT4 add_3132_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n35155), 
            .O(n6563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13397_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18681));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13398_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18682));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_2_lut (.I0(n410), .I1(\PID_CONTROLLER.result [10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4617));   // verilog/motorControl.v(32[23:29])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3132_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n35154), 
            .O(n6564)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_16 (.CI(n35154), .I0(n2070), .I1(n86), .CO(n35155));
    SB_LUT4 add_3132_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n35153), 
            .O(n6565)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_15 (.CI(n35153), .I0(n2071), .I1(n87), .CO(n35154));
    SB_LUT4 i13399_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18683));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13039_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n41851), 
            .I3(GND_net), .O(n18323));   // verilog/coms.v(126[12] 289[6])
    defparam i13039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13400_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18684));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13401_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18685));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4761));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4583), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i809_3_lut (.I0(n516), .I1(n6462), .I2(n1193), .I3(GND_net), 
            .O(n1299));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13402_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18686));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i890_3_lut (.I0(n1299), .I1(n6472), .I2(n1316), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i969_3_lut (.I0(n1419), .I1(n6483), .I2(n1436), .I3(GND_net), 
            .O(n1536));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1046_3_lut (.I0(n1536), .I1(n6495), .I2(n1553), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1121_3_lut (.I0(n1650), .I1(n6508), .I2(n1667), .I3(GND_net), 
            .O(n1761));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3132_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n35152), 
            .O(n6566)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1194_3_lut (.I0(n1761), .I1(n6522), .I2(n1778), .I3(GND_net), 
            .O(n1869));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1265_3_lut (.I0(n1869), .I1(n6537), .I2(n1886), .I3(GND_net), 
            .O(n1974));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4759));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3132_14 (.CI(n35152), .I0(n2072), .I1(n88), .CO(n35153));
    SB_LUT4 div_15_i1271_3_lut (.I0(n522), .I1(n6543), .I2(n1886), .I3(GND_net), 
            .O(n1980));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13403_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18687));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13040_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n41851), 
            .I3(GND_net), .O(n18324));   // verilog/coms.v(126[12] 289[6])
    defparam i13040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13404_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18688));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13405_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18689));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13406_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18690));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13407_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18691));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13408_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18692));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3132_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n35151), 
            .O(n6567)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_13 (.CI(n35151), .I0(n2073), .I1(n89), .CO(n35152));
    SB_LUT4 i13409_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18693));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13410_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18694));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13411_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18695));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13412_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18696));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13413_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18697));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13041_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n41851), 
            .I3(GND_net), .O(n18325));   // verilog/coms.v(126[12] 289[6])
    defparam i13041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13414_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n18698));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3132_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n35150), 
            .O(n6568)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_12 (.CI(n35150), .I0(n2074), .I1(n90), .CO(n35151));
    SB_LUT4 add_3132_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n35149), 
            .O(n6569)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25_2_lut (.I0(n416), .I1(\PID_CONTROLLER.result [4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4615));   // verilog/motorControl.v(32[23:29])
    defparam i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3132_11 (.CI(n35149), .I0(n2075), .I1(n91), .CO(n35150));
    SB_LUT4 add_3132_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n35148), 
            .O(n6570)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_10 (.CI(n35148), .I0(n2076), .I1(n92), .CO(n35149));
    SB_LUT4 add_3132_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n35147), 
            .O(n6571)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_2_lut_adj_1572 (.I0(n403), .I1(\PID_CONTROLLER.result [17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4619));   // verilog/motorControl.v(32[23:29])
    defparam i7_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i17_2_lut (.I0(n414), .I1(\PID_CONTROLLER.result [6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4616));   // verilog/motorControl.v(32[23:29])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13417_4_lut (.I0(n27708), .I1(r_Clock_Count[0]), .I2(n226), 
            .I3(n17657), .O(n18701));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13417_4_lut.LUT_INIT = 16'ha088;
    SB_CARRY add_3132_9 (.CI(n35147), .I0(n2077), .I1(n93), .CO(n35148));
    SB_LUT4 add_3132_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n35146), 
            .O(n6572)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_8 (.CI(n35146), .I0(n2078), .I1(n94), .CO(n35147));
    SB_LUT4 i15_2_lut_adj_1573 (.I0(n407), .I1(\PID_CONTROLLER.result [13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4618));   // verilog/motorControl.v(32[23:29])
    defparam i15_2_lut_adj_1573.LUT_INIT = 16'h6666;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n46632), .I2(n43079), .I3(GND_net), 
            .O(n40132));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3132_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n35145), 
            .O(n6573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4659), .I3(n35588), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_15_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4660), .I3(n35587), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_7 (.CI(n35145), .I0(n2079), .I1(n95), .CO(n35146));
    SB_LUT4 add_3132_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n35144), 
            .O(n6574)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_24 (.CI(n35587), .I0(GND_net), .I1(n3_adj_4660), 
            .CO(n35588));
    SB_CARRY add_3132_6 (.CI(n35144), .I0(n2080), .I1(n96), .CO(n35145));
    SB_LUT4 add_3132_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n35143), 
            .O(n6575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4661), .I3(n35586), .O(n4_adj_4587)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_23 (.CI(n35586), .I0(GND_net), .I1(n4_adj_4661), 
            .CO(n35587));
    SB_DFF color_i17 (.Q(color[16]), .C(clk32MHz), .D(color_23__N_1[16]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_CARRY add_3132_5 (.CI(n35143), .I0(n2081), .I1(n97), .CO(n35144));
    SB_LUT4 i13_3_lut_adj_1574 (.I0(bit_ctr[5]), .I1(n46633), .I2(n43079), 
            .I3(GND_net), .O(n40136));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1574.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1575 (.I0(bit_ctr[6]), .I1(n46634), .I2(n43079), 
            .I3(GND_net), .O(n40140));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1575.LUT_INIT = 16'hacac;
    SB_LUT4 add_3132_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n35142), 
            .O(n6576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF color_i16 (.Q(color[15]), .C(clk32MHz), .D(color_23__N_1[15]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i15 (.Q(color[14]), .C(clk32MHz), .D(color_23__N_1[14]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i14 (.Q(color[13]), .C(clk32MHz), .D(color_23__N_1[13]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i13 (.Q(color[12]), .C(clk32MHz), .D(color_23__N_1[12]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i12 (.Q(color[11]), .C(clk32MHz), .D(color_23__N_1[11]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i11 (.Q(color[10]), .C(clk32MHz), .D(color_23__N_1[10]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i10 (.Q(color[9]), .C(clk32MHz), .D(color_23__N_1[9]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i9 (.Q(color[8]), .C(clk32MHz), .D(color_23__N_1[8]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i8 (.Q(color[7]), .C(clk32MHz), .D(color_23__N_1[7]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i7 (.Q(color[6]), .C(clk32MHz), .D(color_23__N_1[6]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i6 (.Q(color[5]), .C(clk32MHz), .D(color_23__N_1[5]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i5 (.Q(color[4]), .C(clk32MHz), .D(color_23__N_1[4]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i4 (.Q(color[3]), .C(clk32MHz), .D(color_23__N_1[3]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i3 (.Q(color[2]), .C(clk32MHz), .D(color_23__N_1[2]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i2 (.Q(color[1]), .C(clk32MHz), .D(color_23__N_1[1]));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_25[23]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_25[22]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_LUT4 i13_3_lut_adj_1576 (.I0(bit_ctr[7]), .I1(n46635), .I2(n43079), 
            .I3(GND_net), .O(n40144));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1576.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1137_i26_4_lut (.I0(n521), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4662), .I3(n35585), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_22 (.CI(n35585), .I0(GND_net), .I1(n5_adj_4662), 
            .CO(n35586));
    SB_LUT4 div_15_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4750));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_25[21]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_25[20]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_25[19]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_25[18]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_25[17]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_25[16]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_25[15]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_25[14]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_25[13]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_25[12]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_25[11]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_25[10]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_25[9]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_25[8]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_25[7]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_25[6]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_25[5]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_25[4]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_25[3]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_25[2]));   // verilog/TinyFPGA_B.v(179[10] 181[6])
    SB_LUT4 div_15_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4663), .I3(n35584), .O(n6_adj_4586)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_21 (.CI(n35584), .I0(GND_net), .I1(n6_adj_4663), 
            .CO(n35585));
    SB_LUT4 div_15_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4664), .I3(n35583), .O(n7_adj_4585)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38904_4_lut (.I0(n29_adj_4756), .I1(n27_adj_4754), .I2(n25_adj_4752), 
            .I3(n23_adj_4750), .O(n46806));
    defparam i38904_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY div_15_unary_minus_2_add_3_20 (.CI(n35583), .I0(GND_net), .I1(n7_adj_4664), 
            .CO(n35584));
    SB_LUT4 i38900_4_lut (.I0(n35_adj_4761), .I1(n33_adj_4759), .I2(n31_adj_4758), 
            .I3(n46806), .O(n46802));
    defparam i38900_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4665), .I3(n35582), .O(n8_adj_4584)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1281_i22_4_lut (.I0(n523), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4749));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_1281_i30_3_lut (.I0(n28_adj_4755), .I1(n93), 
            .I2(n33_adj_4759), .I3(GND_net), .O(n30_adj_4757));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3132_4 (.CI(n35142), .I0(n2082), .I1(n98), .CO(n35143));
    SB_CARRY div_15_unary_minus_2_add_3_19 (.CI(n35582), .I0(GND_net), .I1(n8_adj_4665), 
            .CO(n35583));
    SB_LUT4 div_15_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4666), .I3(n35581), .O(n9_adj_4583)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1281_i34_3_lut (.I0(n26_adj_4753), .I1(n91), 
            .I2(n37_adj_4762), .I3(GND_net), .O(n34_adj_4760));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13_3_lut_adj_1577 (.I0(bit_ctr[8]), .I1(n46636), .I2(n43079), 
            .I3(GND_net), .O(n40148));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1577.LUT_INIT = 16'hacac;
    SB_LUT4 i41031_4_lut (.I0(n34_adj_4760), .I1(n24_adj_4751), .I2(n37_adj_4762), 
            .I3(n46800), .O(n48934));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41031_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41032_3_lut (.I0(n48934), .I1(n90), .I2(n39_adj_4763), .I3(GND_net), 
            .O(n48935));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41032_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_15_unary_minus_2_add_3_18 (.CI(n35581), .I0(GND_net), .I1(n9_adj_4666), 
            .CO(n35582));
    SB_LUT4 i40933_3_lut (.I0(n48935), .I1(n89), .I2(n41_adj_4764), .I3(GND_net), 
            .O(n48836));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40933_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4667), .I3(n35580), .O(n10_adj_4582)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40530_4_lut (.I0(n41_adj_4764), .I1(n39_adj_4763), .I2(n37_adj_4762), 
            .I3(n46802), .O(n48433));
    defparam i40530_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i40739_4_lut (.I0(n30_adj_4757), .I1(n22_adj_4749), .I2(n33_adj_4759), 
            .I3(n46804), .O(n48642));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40739_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40852_3_lut (.I0(n48836), .I1(n88), .I2(n43_adj_4766), .I3(GND_net), 
            .O(n42_adj_4765));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40852_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40958_4_lut (.I0(n42_adj_4765), .I1(n48642), .I2(n43_adj_4766), 
            .I3(n48433), .O(n48861));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40958_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40959_3_lut (.I0(n48861), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n48862));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40959_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY div_15_unary_minus_2_add_3_17 (.CI(n35580), .I0(GND_net), .I1(n10_adj_4667), 
            .CO(n35581));
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n48862), .I1(n16651), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'hceef;
    SB_LUT4 add_3132_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n35141), 
            .O(n6577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4668), .I3(n35579), .O(n11_adj_4581)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_16 (.CI(n35579), .I0(GND_net), .I1(n11_adj_4668), 
            .CO(n35580));
    SB_CARRY add_3132_3 (.CI(n35141), .I0(n2083), .I1(n99), .CO(n35142));
    SB_LUT4 div_15_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4669), .I3(n35578), .O(n12_adj_4580)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3132_2_lut (.I0(GND_net), .I1(n524), .I2(n558), .I3(VCC_net), 
            .O(n6578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3132_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_15 (.CI(n35578), .I0(GND_net), .I1(n12_adj_4669), 
            .CO(n35579));
    SB_LUT4 div_15_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4670), .I3(n35577), .O(n13_adj_4579)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_adj_1579 (.I0(bit_ctr[9]), .I1(n46637), .I2(n43079), 
            .I3(GND_net), .O(n40152));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1579.LUT_INIT = 16'hacac;
    SB_LUT4 i13042_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n41851), 
            .I3(GND_net), .O(n18326));   // verilog/coms.v(126[12] 289[6])
    defparam i13042_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_2_add_3_14 (.CI(n35577), .I0(GND_net), .I1(n13_adj_4670), 
            .CO(n35578));
    SB_LUT4 div_15_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4671), .I3(n35576), .O(n14_adj_4578)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_13 (.CI(n35576), .I0(GND_net), .I1(n14_adj_4671), 
            .CO(n35577));
    SB_LUT4 div_15_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4672), .I3(n35575), .O(n15_adj_4577)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3132_2 (.CI(VCC_net), .I0(n524), .I1(n558), .CO(n35141));
    SB_CARRY div_15_unary_minus_2_add_3_12 (.CI(n35575), .I0(GND_net), .I1(n15_adj_4672), 
            .CO(n35576));
    SB_LUT4 div_15_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4673), .I3(n35574), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_11 (.CI(n35574), .I0(GND_net), .I1(n16_adj_4673), 
            .CO(n35575));
    SB_LUT4 div_15_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4674), .I3(n35573), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_10 (.CI(n35573), .I0(GND_net), .I1(n17_adj_4674), 
            .CO(n35574));
    SB_LUT4 div_15_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4675), .I3(n35572), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1187_3_lut (.I0(n1754), .I1(n6515), .I2(n1778), .I3(GND_net), 
            .O(n1862));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1187_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_2_add_3_9 (.CI(n35572), .I0(GND_net), .I1(n18_adj_4675), 
            .CO(n35573));
    SB_LUT4 div_15_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1580 (.I0(n97), .I1(n16617), .I2(GND_net), .I3(GND_net), 
            .O(n16688));
    defparam i1_2_lut_adj_1580.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n224), .I1(n99), .I2(n16614), .I3(n558), 
            .O(n5_adj_4603));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'h555d;
    SB_LUT4 i13_3_lut_adj_1582 (.I0(bit_ctr[10]), .I1(n46638), .I2(n43079), 
            .I3(GND_net), .O(n40156));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1582.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4676), .I3(n35571), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_8 (.CI(n35571), .I0(GND_net), .I1(n19_adj_4676), 
            .CO(n35572));
    SB_LUT4 div_15_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4677), .I3(n35570), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_7 (.CI(n35570), .I0(GND_net), .I1(n20_adj_4677), 
            .CO(n35571));
    SB_LUT4 i13_3_lut_adj_1583 (.I0(bit_ctr[11]), .I1(n46639), .I2(n43079), 
            .I3(GND_net), .O(n40160));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1583.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4678), .I3(n35569), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_6 (.CI(n35569), .I0(GND_net), .I1(n21_adj_4678), 
            .CO(n35570));
    SB_LUT4 div_15_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4679), .I3(n35568), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_adj_1584 (.I0(bit_ctr[12]), .I1(n46640), .I2(n43079), 
            .I3(GND_net), .O(n40164));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1584.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_2_add_3_5 (.CI(n35568), .I0(GND_net), .I1(n22_adj_4679), 
            .CO(n35569));
    SB_LUT4 div_15_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4680), .I3(n35567), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_4 (.CI(n35567), .I0(GND_net), .I1(n23_adj_4680), 
            .CO(n35568));
    SB_LUT4 div_15_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4681), .I3(n35566), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_3 (.CI(n35566), .I0(GND_net), .I1(n24_adj_4681), 
            .CO(n35567));
    SB_LUT4 i1_2_lut_adj_1585 (.I0(n17980), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41224));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'h8888;
    SB_LUT4 div_15_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4682), .I3(VCC_net), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4682), 
            .CO(n35566));
    SB_LUT4 div_15_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4635), .I3(n35565), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_15_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4636), .I3(n35564), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_24 (.CI(n35564), .I0(GND_net), .I1(n3_adj_4636), 
            .CO(n35565));
    SB_LUT4 div_15_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4637), .I3(n35563), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_23 (.CI(n35563), .I0(GND_net), .I1(n4_adj_4637), 
            .CO(n35564));
    SB_LUT4 i39059_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n46549));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39059_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_15_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4638), .I3(n35562), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n46549), .I1(n16614), .I2(n99), .I3(n5_adj_4603), 
            .O(n392));
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'hefce;
    SB_LUT4 div_15_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28734_2_lut (.I0(n511), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4562));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28734_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i39468_3_lut (.I0(n369), .I1(n558), .I2(n392), .I3(GND_net), 
            .O(n510));
    defparam i39468_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY div_15_unary_minus_4_add_3_22 (.CI(n35562), .I0(GND_net), .I1(n5_adj_4638), 
            .CO(n35563));
    SB_LUT4 div_15_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n512));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28831_2_lut (.I0(n513), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28831_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i39425_3_lut (.I0(n512), .I1(n558), .I2(n671), .I3(GND_net), 
            .O(n785));
    defparam i39425_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_15_i460_4_lut (.I0(n649), .I1(n2_adj_4972), .I2(n671), 
            .I3(n99), .O(n784));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i460_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4639), .I3(n35561), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_297_i46_4_lut (.I0(n511), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(n17977), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41130));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(n17955), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41074));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h8888;
    SB_LUT4 i13_3_lut_adj_1589 (.I0(bit_ctr[13]), .I1(n46641), .I2(n43079), 
            .I3(GND_net), .O(n40168));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1589.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_21 (.CI(n35561), .I0(GND_net), .I1(n6_adj_4639), 
            .CO(n35562));
    SB_LUT4 div_15_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4640), .I3(n35560), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_adj_1590 (.I0(bit_ctr[14]), .I1(n46642), .I2(n43079), 
            .I3(GND_net), .O(n40172));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1590.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1591 (.I0(bit_ctr[15]), .I1(n46643), .I2(n43079), 
            .I3(GND_net), .O(n40176));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1591.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_20 (.CI(n35560), .I0(GND_net), .I1(n7_adj_4640), 
            .CO(n35561));
    SB_LUT4 div_15_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4641), .I3(n35559), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n46), .I1(n16688), .I2(n98), .I3(n42499), 
            .O(n533));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'hefce;
    SB_LUT4 div_15_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4587), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28799_2_lut (.I0(n512), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4972));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28799_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_15_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i39467_3_lut (.I0(n511), .I1(n558), .I2(n533), .I3(GND_net), 
            .O(n649));
    defparam i39467_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_15_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_390_i44_4_lut (.I0(n512), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40575_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n48478));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40575_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13_3_lut_adj_1593 (.I0(bit_ctr[16]), .I1(n46644), .I2(n43079), 
            .I3(GND_net), .O(n40180));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1593.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1594 (.I0(n48478), .I1(n16617), .I2(n97), .I3(n42501), 
            .O(n671));
    defparam i1_4_lut_adj_1594.LUT_INIT = 16'hefce;
    SB_LUT4 div_15_i368_4_lut (.I0(n510), .I1(n2_adj_4562), .I2(n533), 
            .I3(n99), .O(n648));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i368_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i28847_3_lut (.I0(n784), .I1(n98), .I2(n4), .I3(GND_net), 
            .O(n6_adj_4559));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28847_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_15_i459_4_lut (.I0(n648), .I1(n4_adj_4965), .I2(n671), 
            .I3(n98), .O(n783));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i459_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_i548_4_lut (.I0(n783), .I1(n6_adj_4559), .I2(n806), 
            .I3(n97), .O(n915));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i548_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_15_i635_3_lut (.I0(n915), .I1(n6439), .I2(n938), .I3(GND_net), 
            .O(n1044));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i720_3_lut (.I0(n1044), .I1(n6447), .I2(n1067), .I3(GND_net), 
            .O(n1170));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i720_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_19 (.CI(n35559), .I0(GND_net), .I1(n8_adj_4641), 
            .CO(n35560));
    SB_LUT4 div_15_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4642), .I3(n35558), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i803_3_lut (.I0(n1170), .I1(n6456), .I2(n1193), .I3(GND_net), 
            .O(n1293));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i884_3_lut (.I0(n1293), .I1(n6466), .I2(n1316), .I3(GND_net), 
            .O(n1413));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i963_3_lut (.I0(n1413), .I1(n6477), .I2(n1436), .I3(GND_net), 
            .O(n1530));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1040_3_lut (.I0(n1530), .I1(n6489), .I2(n1553), .I3(GND_net), 
            .O(n1644));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1115_3_lut (.I0(n1644), .I1(n6502), .I2(n1667), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1188_3_lut (.I0(n1755), .I1(n6516), .I2(n1778), .I3(GND_net), 
            .O(n1863));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4748));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4584), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i725_3_lut (.I0(n515), .I1(n6452), .I2(n1067), .I3(GND_net), 
            .O(n1175));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i808_3_lut (.I0(n1175), .I1(n6461), .I2(n1193), .I3(GND_net), 
            .O(n1298));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1595 (.I0(bit_ctr[17]), .I1(n46645), .I2(n43079), 
            .I3(GND_net), .O(n40184));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1595.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_18 (.CI(n35558), .I0(GND_net), .I1(n9_adj_4642), 
            .CO(n35559));
    SB_LUT4 div_15_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4643), .I3(n35557), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_17 (.CI(n35557), .I0(GND_net), .I1(n10_adj_4643), 
            .CO(n35558));
    SB_LUT4 div_15_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4644), .I3(n35556), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_16 (.CI(n35556), .I0(GND_net), .I1(n11_adj_4644), 
            .CO(n35557));
    SB_LUT4 div_15_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4645), .I3(n35555), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_15 (.CI(n35555), .I0(GND_net), .I1(n12_adj_4645), 
            .CO(n35556));
    SB_LUT4 div_15_i889_3_lut (.I0(n1298), .I1(n6471), .I2(n1316), .I3(GND_net), 
            .O(n1418));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i968_3_lut (.I0(n1418), .I1(n6482), .I2(n1436), .I3(GND_net), 
            .O(n1535));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1045_3_lut (.I0(n1535), .I1(n6494), .I2(n1553), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1120_3_lut (.I0(n1649), .I1(n6507), .I2(n1667), .I3(GND_net), 
            .O(n1760));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_i1193_3_lut (.I0(n1760), .I1(n6521), .I2(n1778), .I3(GND_net), 
            .O(n1868));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4741));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_481_i42_4_lut (.I0(n513), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40492_3_lut (.I0(n42), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n48395));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40492_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13_3_lut_adj_1596 (.I0(bit_ctr[18]), .I1(n46646), .I2(n43079), 
            .I3(GND_net), .O(n40188));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1596.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1597 (.I0(bit_ctr[19]), .I1(n46647), .I2(n43079), 
            .I3(GND_net), .O(n40192));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1597.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4646), .I3(n35554), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_14 (.CI(n35554), .I0(GND_net), .I1(n13_adj_4646), 
            .CO(n35555));
    SB_LUT4 div_15_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4647), .I3(n35553), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_13 (.CI(n35553), .I0(GND_net), .I1(n14_adj_4647), 
            .CO(n35554));
    SB_LUT4 i40493_3_lut (.I0(n48395), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n48396));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40493_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1598 (.I0(n48396), .I1(n16621), .I2(n96), .I3(n42503), 
            .O(n806));
    defparam i1_4_lut_adj_1598.LUT_INIT = 16'hefce;
    SB_LUT4 div_15_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4586), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4648), .I3(n35552), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_570_i40_4_lut (.I0(n514), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_570_i44_3_lut (.I0(n42_adj_4683), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4684));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_15_unary_minus_4_add_3_12 (.CI(n35552), .I0(GND_net), .I1(n15_adj_4648), 
            .CO(n35553));
    SB_LUT4 i40579_4_lut (.I0(n44_adj_4684), .I1(n40), .I2(n45), .I3(n47061), 
            .O(n48482));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40579_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1599 (.I0(n48482), .I1(n16624), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1599.LUT_INIT = 16'hceef;
    SB_LUT4 i39420_3_lut (.I0(n513), .I1(n558), .I2(n806), .I3(GND_net), 
            .O(n918));
    defparam i39420_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_15_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4649), .I3(n35551), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_11 (.CI(n35551), .I0(GND_net), .I1(n16_adj_4649), 
            .CO(n35552));
    SB_LUT4 div_15_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4650), .I3(n35550), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_10 (.CI(n35550), .I0(GND_net), .I1(n17_adj_4650), 
            .CO(n35551));
    SB_LUT4 div_15_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4651), .I3(n35549), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_657_i38_4_lut (.I0(n515), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_657_i42_3_lut (.I0(n40_adj_4685), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4686));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40938_4_lut (.I0(n42_adj_4686), .I1(n38), .I2(n43), .I3(n47055), 
            .O(n48841));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40938_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40939_3_lut (.I0(n48841), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n48842));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40939_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1600 (.I0(n48842), .I1(n16627), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1600.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i638_3_lut (.I0(n918), .I1(n6442), .I2(n938), .I3(GND_net), 
            .O(n1047));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13043_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n41851), 
            .I3(GND_net), .O(n18327));   // verilog/coms.v(126[12] 289[6])
    defparam i13043_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_9 (.CI(n35549), .I0(GND_net), .I1(n18_adj_4651), 
            .CO(n35550));
    SB_LUT4 div_15_LessThan_742_i36_4_lut (.I0(n516), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_742_i40_3_lut (.I0(n38_adj_4687), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4688));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40976_4_lut (.I0(n40_adj_4688), .I1(n36), .I2(n41), .I3(n47041), 
            .O(n48879));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40976_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_15_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4652), .I3(n35548), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_8 (.CI(n35548), .I0(GND_net), .I1(n19_adj_4652), 
            .CO(n35549));
    SB_LUT4 div_15_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4653), .I3(n35547), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_7 (.CI(n35547), .I0(GND_net), .I1(n20_adj_4653), 
            .CO(n35548));
    SB_LUT4 div_15_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4654), .I3(n35546), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_6_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b011001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_24_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b000001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13_3_lut_adj_1601 (.I0(bit_ctr[20]), .I1(n46648), .I2(n43079), 
            .I3(GND_net), .O(n40196));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1601.LUT_INIT = 16'hacac;
    SB_CARRY div_15_unary_minus_4_add_3_6 (.CI(n35546), .I0(GND_net), .I1(n21_adj_4654), 
            .CO(n35547));
    SB_LUT4 div_15_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4655), .I3(n35545), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_5 (.CI(n35545), .I0(GND_net), .I1(n22_adj_4655), 
            .CO(n35546));
    SB_LUT4 div_15_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4656), .I3(n35544), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_4 (.CI(n35544), .I0(GND_net), .I1(n23_adj_4656), 
            .CO(n35545));
    SB_LUT4 div_15_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4657), .I3(n35543), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40977_3_lut (.I0(n48879), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n48880));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40977_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i40792_3_lut (.I0(n48880), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n48695));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40792_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(n48695), .I1(n16630), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i723_3_lut (.I0(n1047), .I1(n6450), .I2(n1067), .I3(GND_net), 
            .O(n1173));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_825_i34_4_lut (.I0(n517), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40841_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4692), .I3(GND_net), 
            .O(n48744));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40841_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40842_3_lut (.I0(n48744), .I1(n94), .I2(n43_adj_4693), .I3(GND_net), 
            .O(n48745));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40842_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_15_unary_minus_4_add_3_3 (.CI(n35543), .I0(GND_net), .I1(n24_adj_4657), 
            .CO(n35544));
    SB_LUT4 i39893_4_lut (.I0(n43_adj_4693), .I1(n41_adj_4692), .I2(n39_adj_4691), 
            .I3(n47021), .O(n47796));
    defparam i39893_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_15_LessThan_825_i38_3_lut (.I0(n36_adj_4689), .I1(n96), 
            .I2(n39_adj_4691), .I3(GND_net), .O(n38_adj_4690));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13_3_lut_adj_1603 (.I0(bit_ctr[21]), .I1(n46649), .I2(n43079), 
            .I3(GND_net), .O(n40200));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1603.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4658), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_15_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_15_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4658), 
            .CO(n35543));
    SB_LUT4 i13044_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n41851), 
            .I3(GND_net), .O(n18328));   // verilog/coms.v(126[12] 289[6])
    defparam i13044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40584_3_lut (.I0(n48745), .I1(n93), .I2(n45_adj_4695), .I3(GND_net), 
            .O(n44_adj_4694));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40584_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40327_4_lut (.I0(n44_adj_4694), .I1(n38_adj_4690), .I2(n45_adj_4695), 
            .I3(n47796), .O(n48230));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40327_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n48230), .I1(n16633), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i806_3_lut (.I0(n1173), .I1(n6459), .I2(n1193), .I3(GND_net), 
            .O(n1296));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_906_i32_4_lut (.I0(n518), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40757_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4697), .I3(GND_net), 
            .O(n48660));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40757_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40758_3_lut (.I0(n48660), .I1(n94), .I2(n41_adj_4698), .I3(GND_net), 
            .O(n48661));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40758_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39876_4_lut (.I0(n41_adj_4698), .I1(n39_adj_4697), .I2(n37), 
            .I3(n46992), .O(n47779));
    defparam i39876_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40329_3_lut (.I0(n34_adj_4696), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n48232));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40329_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13045_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n41851), 
            .I3(GND_net), .O(n18329));   // verilog/coms.v(126[12] 289[6])
    defparam i13045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40586_3_lut (.I0(n48661), .I1(n93), .I2(n43_adj_4699), .I3(GND_net), 
            .O(n48489));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40586_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40755_4_lut (.I0(n48489), .I1(n48232), .I2(n43_adj_4699), 
            .I3(n47779), .O(n48658));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40755_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40756_3_lut (.I0(n48658), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n48659));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40756_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1605 (.I0(n48659), .I1(n16636), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1605.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i887_3_lut (.I0(n1296), .I1(n6469), .I2(n1316), .I3(GND_net), 
            .O(n1416));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i39063_4_lut (.I0(n37_adj_4703), .I1(n35_adj_4702), .I2(n33), 
            .I3(n31), .O(n46965));
    defparam i39063_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13158_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18442));   // verilog/coms.v(126[12] 289[6])
    defparam i13158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1606 (.I0(bit_ctr[22]), .I1(n46650), .I2(n43079), 
            .I3(GND_net), .O(n40204));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1606.LUT_INIT = 16'hacac;
    SB_LUT4 add_3131_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n35118), 
            .O(n6546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n35117), 
            .O(n6547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_15 (.CI(n35117), .I0(n1968), .I1(n87), .CO(n35118));
    SB_LUT4 div_15_LessThan_985_i42_3_lut (.I0(n34_adj_4701), .I1(n91), 
            .I2(n45_adj_4708), .I3(GND_net), .O(n42_adj_4706));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_985_i30_4_lut (.I0(n519), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40753_3_lut (.I0(n30), .I1(n95), .I2(n37_adj_4703), .I3(GND_net), 
            .O(n48656));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40753_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40754_3_lut (.I0(n48656), .I1(n94), .I2(n39_adj_4704), .I3(GND_net), 
            .O(n48657));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40754_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39049_4_lut (.I0(n43_adj_4707), .I1(n41_adj_4705), .I2(n39_adj_4704), 
            .I3(n46965), .O(n46951));
    defparam i39049_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40331_4_lut (.I0(n42_adj_4706), .I1(n32_adj_4700), .I2(n45_adj_4708), 
            .I3(n46947), .O(n48234));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40331_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40592_3_lut (.I0(n48657), .I1(n93), .I2(n41_adj_4705), .I3(GND_net), 
            .O(n48495));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40592_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40845_4_lut (.I0(n48495), .I1(n48234), .I2(n45_adj_4708), 
            .I3(n46951), .O(n48748));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40845_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13_3_lut_adj_1607 (.I0(bit_ctr[23]), .I1(n46651), .I2(n43079), 
            .I3(GND_net), .O(n40208));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1607.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1608 (.I0(bit_ctr[24]), .I1(n46652), .I2(n43079), 
            .I3(GND_net), .O(n40212));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1608.LUT_INIT = 16'hacac;
    SB_LUT4 add_3131_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n35116), 
            .O(n6548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_14 (.CI(n35116), .I0(n1969), .I1(n88), .CO(n35117));
    SB_LUT4 add_3131_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n35115), 
            .O(n6549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(n48748), .I1(n16639), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i966_3_lut (.I0(n1416), .I1(n6480), .I2(n1436), .I3(GND_net), 
            .O(n1533));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4709));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i39006_4_lut (.I0(n35_adj_4714), .I1(n33_adj_4713), .I2(n31_adj_4711), 
            .I3(n29_adj_4709), .O(n46908));
    defparam i39006_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3131_13 (.CI(n35115), .I0(n1970), .I1(n89), .CO(n35116));
    SB_LUT4 i13_3_lut_adj_1610 (.I0(bit_ctr[25]), .I1(n46653), .I2(n43079), 
            .I3(GND_net), .O(n40216));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1610.LUT_INIT = 16'hacac;
    SB_LUT4 i34815_4_lut (.I0(n20911), .I1(state[1]), .I2(state[0]), .I3(n16572), 
            .O(n41781));
    defparam i34815_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i13_3_lut_adj_1611 (.I0(bit_ctr[26]), .I1(n46654), .I2(n43079), 
            .I3(GND_net), .O(n40220));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1611.LUT_INIT = 16'hacac;
    SB_LUT4 add_3131_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n35114), 
            .O(n6550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_12 (.CI(n35114), .I0(n1971), .I1(n90), .CO(n35115));
    SB_LUT4 div_15_LessThan_1062_i40_3_lut (.I0(n32_adj_4712), .I1(n91), 
            .I2(n43_adj_4719), .I3(GND_net), .O(n40_adj_4717));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_1062_i28_4_lut (.I0(n520), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40751_3_lut (.I0(n28), .I1(n95), .I2(n35_adj_4714), .I3(GND_net), 
            .O(n48654));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40751_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40752_3_lut (.I0(n48654), .I1(n94), .I2(n37_adj_4715), .I3(GND_net), 
            .O(n48655));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40752_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i38990_4_lut (.I0(n41_adj_4718), .I1(n39_adj_4716), .I2(n37_adj_4715), 
            .I3(n46908), .O(n46892));
    defparam i38990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40749_4_lut (.I0(n40_adj_4717), .I1(n30_adj_4710), .I2(n43_adj_4719), 
            .I3(n46889), .O(n48652));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40749_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40594_3_lut (.I0(n48655), .I1(n93), .I2(n39_adj_4716), .I3(GND_net), 
            .O(n48497));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40594_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13_3_lut_adj_1612 (.I0(bit_ctr[27]), .I1(n46655), .I2(n43079), 
            .I3(GND_net), .O(n40224));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1612.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1613 (.I0(bit_ctr[28]), .I1(n46656), .I2(n43079), 
            .I3(GND_net), .O(n40228));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1613.LUT_INIT = 16'hacac;
    SB_LUT4 add_3131_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n35113), 
            .O(n6551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_11 (.CI(n35113), .I0(n1972), .I1(n91), .CO(n35114));
    SB_LUT4 add_3131_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n35112), 
            .O(n6552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_adj_1614 (.I0(bit_ctr[29]), .I1(n46657), .I2(n43079), 
            .I3(GND_net), .O(n40232));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1614.LUT_INIT = 16'hacac;
    SB_LUT4 i28686_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4976));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28686_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_15_i274_4_lut (.I0(n5_adj_4603), .I1(n2_adj_4976), .I2(n392), 
            .I3(n99), .O(n42499));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i274_4_lut.LUT_INIT = 16'ha9a6;
    SB_CARRY add_3131_10 (.CI(n35112), .I0(n1973), .I1(n92), .CO(n35113));
    SB_LUT4 div_15_i367_4_lut (.I0(n42499), .I1(n4_adj_4561), .I2(n533), 
            .I3(n98), .O(n42501));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i367_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i28815_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_4965), .I3(GND_net), 
            .O(n6_adj_4964));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28815_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_15_i458_4_lut (.I0(n42501), .I1(n6_adj_4964), .I2(n671), 
            .I3(n97), .O(n42503));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i458_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 add_3131_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n35111), 
            .O(n6553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_9 (.CI(n35111), .I0(n1974), .I1(n93), .CO(n35112));
    SB_LUT4 i28855_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4559), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28855_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_15_i547_4_lut (.I0(n42503), .I1(n8), .I2(n806), .I3(n96), 
            .O(n914));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i547_4_lut.LUT_INIT = 16'h5659;
    SB_LUT4 div_15_i634_3_lut (.I0(n914), .I1(n6438), .I2(n938), .I3(GND_net), 
            .O(n1043));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1615 (.I0(bit_ctr[30]), .I1(n46658), .I2(n43079), 
            .I3(GND_net), .O(n40236));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1615.LUT_INIT = 16'hacac;
    SB_LUT4 add_3131_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n35110), 
            .O(n6554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_118[23]), 
            .I2(n3_adj_4598), .I3(n34867), .O(displacement_23__N_25[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_8 (.CI(n35110), .I0(n1975), .I1(n94), .CO(n35111));
    SB_LUT4 add_3131_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n35109), 
            .O(n6555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_7 (.CI(n35109), .I0(n1976), .I1(n95), .CO(n35110));
    SB_LUT4 add_3131_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n35108), 
            .O(n6556)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_118[22]), 
            .I2(n3_adj_4598), .I3(n34866), .O(displacement_23__N_25[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n34866), .I0(displacement_23__N_118[22]), 
            .I1(n3_adj_4598), .CO(n34867));
    SB_LUT4 i13_3_lut_adj_1616 (.I0(bit_ctr[31]), .I1(n46659), .I2(n43079), 
            .I3(GND_net), .O(n40240));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1616.LUT_INIT = 16'hacac;
    SB_CARRY add_3131_6 (.CI(n35108), .I0(n1977), .I1(n96), .CO(n35109));
    SB_LUT4 add_3131_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n35107), 
            .O(n6557)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13159_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18443));   // verilog/coms.v(126[12] 289[6])
    defparam i13159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12606_4_lut (.I0(n17849), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n17707), .O(n17890));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12606_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i41074_4_lut (.I0(n48497), .I1(n48652), .I2(n43_adj_4719), 
            .I3(n46892), .O(n48977));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41074_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3131_5 (.CI(n35107), .I0(n1978), .I1(n97), .CO(n35108));
    SB_LUT4 add_3131_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n35106), 
            .O(n6558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_4 (.CI(n35106), .I0(n1979), .I1(n98), .CO(n35107));
    SB_LUT4 i12603_4_lut (.I0(n17849), .I1(r_Bit_Index[2]), .I2(n4694), 
            .I3(n17707), .O(n17887));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12603_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i1_2_lut_adj_1617 (.I0(n17872), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41442));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1617.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1618 (.I0(n17869), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41444));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1618.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1619 (.I0(n17866), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41446));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1619.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(r_SM_Main_adj_5024[2]), .I1(n44294), 
            .I2(n44245), .I3(n118), .O(n5_adj_4982));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'haaae;
    SB_LUT4 i1_2_lut_adj_1621 (.I0(n17863), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41336));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1621.LUT_INIT = 16'h8888;
    SB_LUT4 add_3131_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n35105), 
            .O(n6559)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_3 (.CI(n35105), .I0(n1980), .I1(n99), .CO(n35106));
    SB_LUT4 add_3131_2_lut (.I0(GND_net), .I1(n523), .I2(n558), .I3(VCC_net), 
            .O(n6560)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_118[21]), 
            .I2(n3_adj_4598), .I3(n34865), .O(displacement_23__N_25[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n34865), .I0(displacement_23__N_118[21]), 
            .I1(n3_adj_4598), .CO(n34866));
    SB_LUT4 i40747_3_lut (.I0(n26), .I1(n95), .I2(n33_adj_4725), .I3(GND_net), 
            .O(n48650));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40747_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_118[20]), 
            .I2(n3_adj_4598), .I3(n34864), .O(displacement_23__N_25[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_2 (.CI(VCC_net), .I0(n523), .I1(n558), .CO(n35105));
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n34864), .I0(displacement_23__N_118[20]), 
            .I1(n3_adj_4598), .CO(n34865));
    SB_LUT4 add_3130_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n35104), 
            .O(n6530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_15_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_19_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b000001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3130_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n35103), 
            .O(n6531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_14 (.CI(n35103), .I0(n1863), .I1(n88), .CO(n35104));
    SB_LUT4 add_3130_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n35102), 
            .O(n6532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i629_1_lut (.I0(pwm[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(GATES_5__N_3405));   // verilog/TinyFPGA_B.v(44[8:13])
    defparam i629_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3130_13 (.CI(n35102), .I0(n1864), .I1(n89), .CO(n35103));
    SB_LUT4 add_3130_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n35101), 
            .O(n6533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41075_3_lut (.I0(n48977), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n48978));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41075_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY add_3130_12 (.CI(n35101), .I0(n1865), .I1(n90), .CO(n35102));
    SB_LUT4 i1_4_lut_adj_1622 (.I0(n48978), .I1(n16642), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1622.LUT_INIT = 16'hceef;
    SB_LUT4 i40748_3_lut (.I0(n48650), .I1(n94), .I2(n35_adj_4726), .I3(GND_net), 
            .O(n48651));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40748_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i38969_4_lut (.I0(n39_adj_4729), .I1(n37_adj_4727), .I2(n35_adj_4726), 
            .I3(n46877), .O(n46871));
    defparam i38969_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3130_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n35100), 
            .O(n6534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41027_4_lut (.I0(n38_adj_4728), .I1(n28_adj_4721), .I2(n41_adj_4730), 
            .I3(n46865), .O(n48930));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41027_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40598_3_lut (.I0(n48651), .I1(n93), .I2(n37_adj_4727), .I3(GND_net), 
            .O(n48501));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40598_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41141_4_lut (.I0(n48501), .I1(n48930), .I2(n41_adj_4730), 
            .I3(n46871), .O(n49044));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41141_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41142_3_lut (.I0(n49044), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n49045));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41142_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i41102_3_lut (.I0(n49045), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n49005));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41102_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(n49005), .I1(n16645), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i1118_3_lut (.I0(n1647), .I1(n6505), .I2(n1667), .I3(GND_net), 
            .O(n1758));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_i1191_3_lut (.I0(n1758), .I1(n6519), .I2(n1778), .I3(GND_net), 
            .O(n1866));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4744));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4746));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4745));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13160_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18444));   // verilog/coms.v(126[12] 289[6])
    defparam i13160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1043_3_lut (.I0(n1533), .I1(n6492), .I2(n1553), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13163_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18447));   // verilog/coms.v(126[12] 289[6])
    defparam i13163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_50));   // verilog/TinyFPGA_B.v(91[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13161_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18445));   // verilog/coms.v(126[12] 289[6])
    defparam i13161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13162_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18446));   // verilog/coms.v(126[12] 289[6])
    defparam i13162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4732));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6713), 
            .I3(n2724), .O(n41_adj_4960));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6714), 
            .I3(n2724), .O(n39_adj_4959));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n532));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6711), 
            .I3(n2724), .O(n45_adj_4962));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6712), 
            .I3(n2724), .O(n43_adj_4961));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6715), 
            .I3(n2724), .O(n37_adj_4958));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6719), 
            .I3(n2724), .O(n29_adj_4953));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6718), 
            .I3(n2724), .O(n31_adj_4955));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6723), 
            .I3(n2724), .O(n21_adj_4948));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_118[19]), 
            .I2(n6_adj_4576), .I3(n34863), .O(displacement_23__N_25[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6722), 
            .I3(n2724), .O(n23_adj_4949));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY add_3130_11 (.CI(n35100), .I0(n1866), .I1(n91), .CO(n35101));
    SB_LUT4 div_15_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6721), 
            .I3(n2724), .O(n25_adj_4951));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6729), 
            .I3(n2724), .O(n9_adj_4939));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6730), 
            .I3(n2724), .O(n7_adj_4937));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_i1114_3_lut (.I0(n1643), .I1(n6501), .I2(n1667), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1624 (.I0(n87), .I1(n16648), .I2(GND_net), .I3(GND_net), 
            .O(n16645));
    defparam i1_2_lut_adj_1624.LUT_INIT = 16'hdddd;
    SB_LUT4 div_15_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4720));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6716), 
            .I3(n2724), .O(n35_adj_4957));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n34863), .I0(displacement_23__N_118[19]), 
            .I1(n6_adj_4576), .CO(n34864));
    SB_LUT4 i38975_4_lut (.I0(n33_adj_4725), .I1(n31_adj_4724), .I2(n29_adj_4722), 
            .I3(n27_adj_4720), .O(n46877));
    defparam i38975_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6725), 
            .I3(n2724), .O(n17_adj_4946));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6724), 
            .I3(n2724), .O(n19_adj_4947));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_118[18]), 
            .I2(n7), .I3(n34862), .O(displacement_23__N_25[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3130_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n35099), 
            .O(n6535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_631_i15_2_lut (.I0(pwm_count[7]), .I1(pwm[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4627));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6717), 
            .I3(n2724), .O(n33_adj_4956));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 LessThan_631_i9_2_lut (.I0(pwm_count[4]), .I1(pwm[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4624));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6728), 
            .I3(n2724), .O(n11_adj_4941));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6727), 
            .I3(n2724), .O(n13_adj_4943));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_15_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6726), 
            .I3(n2724), .O(n15_adj_4944));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY add_3130_10 (.CI(n35099), .I0(n1867), .I1(n92), .CO(n35100));
    SB_LUT4 add_3130_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n35098), 
            .O(n6536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_9 (.CI(n35098), .I0(n1868), .I1(n93), .CO(n35099));
    SB_LUT4 add_3130_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n35097), 
            .O(n6537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_8 (.CI(n35097), .I0(n1869), .I1(n94), .CO(n35098));
    SB_LUT4 add_3130_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n35096), 
            .O(n6538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_7 (.CI(n35096), .I0(n1870), .I1(n95), .CO(n35097));
    SB_LUT4 add_3130_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n35095), 
            .O(n6539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_6 (.CI(n35095), .I0(n1871), .I1(n96), .CO(n35096));
    SB_LUT4 add_3130_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n35094), 
            .O(n6540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_5 (.CI(n35094), .I0(n1872), .I1(n97), .CO(n35095));
    SB_LUT4 add_3130_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n35093), 
            .O(n6541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_4 (.CI(n35093), .I0(n1873), .I1(n98), .CO(n35094));
    SB_LUT4 add_3130_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n35092), 
            .O(n6542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_3 (.CI(n35092), .I0(n1874), .I1(n99), .CO(n35093));
    SB_LUT4 add_3130_2_lut (.I0(GND_net), .I1(n522), .I2(n558), .I3(VCC_net), 
            .O(n6543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3130_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3130_2 (.CI(VCC_net), .I0(n522), .I1(n558), .CO(n35092));
    SB_LUT4 add_3129_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n35091), 
            .O(n6515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3129_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n35090), 
            .O(n6516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_13 (.CI(n35090), .I0(n1755), .I1(n89), .CO(n35091));
    SB_LUT4 add_3129_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n35089), 
            .O(n6517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_12 (.CI(n35089), .I0(n1756), .I1(n90), .CO(n35090));
    SB_LUT4 add_3129_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n35088), 
            .O(n6518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_11 (.CI(n35088), .I0(n1757), .I1(n91), .CO(n35089));
    SB_LUT4 add_3129_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n35087), 
            .O(n6519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_10 (.CI(n35087), .I0(n1758), .I1(n92), .CO(n35088));
    SB_LUT4 add_3129_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n35086), 
            .O(n6520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_9 (.CI(n35086), .I0(n1759), .I1(n93), .CO(n35087));
    SB_LUT4 add_3129_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n35085), 
            .O(n6521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_8 (.CI(n35085), .I0(n1760), .I1(n94), .CO(n35086));
    SB_LUT4 add_3129_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n35084), 
            .O(n6522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_7 (.CI(n35084), .I0(n1761), .I1(n95), .CO(n35085));
    SB_LUT4 add_3129_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n35083), 
            .O(n6523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_6 (.CI(n35083), .I0(n1762), .I1(n96), .CO(n35084));
    SB_LUT4 add_3129_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n35082), 
            .O(n6524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_5 (.CI(n35082), .I0(n1763), .I1(n97), .CO(n35083));
    SB_LUT4 add_3129_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n35081), 
            .O(n6525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_4 (.CI(n35081), .I0(n1764), .I1(n98), .CO(n35082));
    SB_LUT4 add_3129_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n35080), 
            .O(n6526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_3 (.CI(n35080), .I0(n1765), .I1(n99), .CO(n35081));
    SB_LUT4 add_3129_2_lut (.I0(GND_net), .I1(n521), .I2(n558), .I3(VCC_net), 
            .O(n6527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3129_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3129_2 (.CI(VCC_net), .I0(n521), .I1(n558), .CO(n35080));
    SB_LUT4 div_15_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6720), 
            .I3(n2724), .O(n27_adj_4952));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n34862), .I0(displacement_23__N_118[18]), 
            .I1(n7), .CO(n34863));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_118[17]), 
            .I2(n8_adj_4575), .I3(n34861), .O(displacement_23__N_25[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n34861), .I0(displacement_23__N_118[17]), 
            .I1(n8_adj_4575), .CO(n34862));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_118[16]), 
            .I2(n9), .I3(n34860), .O(displacement_23__N_25[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n34860), .I0(displacement_23__N_118[16]), 
            .I1(n9), .CO(n34861));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_118[15]), 
            .I2(n10), .I3(n34859), .O(displacement_23__N_25[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39531_4_lut (.I0(n27_adj_4952), .I1(n15_adj_4944), .I2(n13_adj_4943), 
            .I3(n11_adj_4941), .O(n47434));
    defparam i39531_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n34859), .I0(displacement_23__N_118[15]), 
            .I1(n10), .CO(n34860));
    SB_LUT4 LessThan_631_i13_2_lut (.I0(pwm_count[6]), .I1(pwm[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4626));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_631_i11_2_lut (.I0(pwm_count[5]), .I1(pwm[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4625));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4956), 
            .I3(GND_net), .O(n12_adj_4942));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_118[14]), 
            .I2(n11), .I3(n34858), .O(displacement_23__N_25[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39525_2_lut (.I0(n33_adj_4956), .I1(n15_adj_4944), .I2(GND_net), 
            .I3(GND_net), .O(n47428));
    defparam i39525_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_15_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4943), 
            .I3(GND_net), .O(n10_adj_4940));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n34858), .I0(displacement_23__N_118[14]), 
            .I1(n11), .CO(n34859));
    SB_LUT4 div_15_LessThan_1830_i30_3_lut (.I0(n12_adj_4942), .I1(n83), 
            .I2(n35_adj_4957), .I3(GND_net), .O(n30_adj_4954));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_118[13]), 
            .I2(n12), .I3(n34857), .O(displacement_23__N_25[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n34857), .I0(displacement_23__N_118[13]), 
            .I1(n12), .CO(n34858));
    SB_LUT4 div_15_i1828_3_lut (.I0(n2720), .I1(n6731), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_118[12]), 
            .I2(n13), .I3(n34856), .O(displacement_23__N_25[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39548_3_lut (.I0(n7_adj_4937), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n47451));
    defparam i39548_3_lut.LUT_INIT = 16'hebeb;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n34856), .I0(displacement_23__N_118[12]), 
            .I1(n13), .CO(n34857));
    SB_LUT4 i40193_4_lut (.I0(n13_adj_4943), .I1(n11_adj_4941), .I2(n9_adj_4939), 
            .I3(n47451), .O(n48096));
    defparam i40193_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40189_4_lut (.I0(n19_adj_4947), .I1(n17_adj_4946), .I2(n15_adj_4944), 
            .I3(n48096), .O(n48092));
    defparam i40189_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_118[11]), 
            .I2(n14), .I3(n34855), .O(displacement_23__N_25[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_631_i4_4_lut (.I0(pwm_count[0]), .I1(pwm[1]), .I2(pwm_count[1]), 
            .I3(pwm[0]), .O(n4_adj_4621));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i40500_3_lut (.I0(n4_adj_4621), .I1(pwm[5]), .I2(n11_adj_4625), 
            .I3(GND_net), .O(n48403));   // verilog/motorControl.v(65[19:32])
    defparam i40500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40966_4_lut (.I0(n25_adj_4951), .I1(n23_adj_4949), .I2(n21_adj_4948), 
            .I3(n48092), .O(n48869));
    defparam i40966_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n34855), .I0(displacement_23__N_118[11]), 
            .I1(n14), .CO(n34856));
    SB_LUT4 i40458_4_lut (.I0(n31_adj_4955), .I1(n29_adj_4953), .I2(n27_adj_4952), 
            .I3(n48869), .O(n48361));
    defparam i40458_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40501_3_lut (.I0(n48403), .I1(pwm[6]), .I2(n13_adj_4626), 
            .I3(GND_net), .O(n48404));   // verilog/motorControl.v(65[19:32])
    defparam i40501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41053_4_lut (.I0(n37_adj_4958), .I1(n35_adj_4957), .I2(n33_adj_4956), 
            .I3(n48361), .O(n48956));
    defparam i41053_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_15_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4961), 
            .I3(GND_net), .O(n16_adj_4945));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i39963_4_lut (.I0(n13_adj_4626), .I1(n11_adj_4625), .I2(n9_adj_4624), 
            .I3(n47079), .O(n47866));
    defparam i39963_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_631_i8_3_lut (.I0(n6_adj_4622), .I1(pwm[4]), .I2(n9_adj_4624), 
            .I3(GND_net), .O(n8_adj_4623));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39835_3_lut (.I0(n48404), .I1(pwm[7]), .I2(n15_adj_4627), 
            .I3(GND_net), .O(n47738));   // verilog/motorControl.v(65[19:32])
    defparam i39835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4937), 
            .I3(GND_net), .O(n6_adj_4936));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i40765_3_lut (.I0(n6_adj_4936), .I1(n90), .I2(n21_adj_4948), 
            .I3(GND_net), .O(n48668));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40765_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40766_3_lut (.I0(n48668), .I1(n89), .I2(n23_adj_4949), .I3(GND_net), 
            .O(n48669));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40766_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40571_4_lut (.I0(n47738), .I1(n8_adj_4623), .I2(n15_adj_4627), 
            .I3(n47866), .O(n48474));   // verilog/motorControl.v(65[19:32])
    defparam i40571_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3128_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n35056), 
            .O(n6501)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39537_4_lut (.I0(n21_adj_4948), .I1(n19_adj_4947), .I2(n17_adj_4946), 
            .I3(n9_adj_4939), .O(n47440));
    defparam i39537_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39489_2_lut (.I0(n43_adj_4961), .I1(n19_adj_4947), .I2(GND_net), 
            .I3(GND_net), .O(n47392));
    defparam i39489_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_15_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4946), 
            .I3(GND_net), .O(n8_adj_4938));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_15_LessThan_1830_i24_3_lut (.I0(n16_adj_4945), .I1(n78), 
            .I2(n45_adj_4962), .I3(GND_net), .O(n24_adj_4950));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39491_4_lut (.I0(n43_adj_4961), .I1(n25_adj_4951), .I2(n23_adj_4949), 
            .I3(n47440), .O(n47394));
    defparam i39491_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40657_4_lut (.I0(n24_adj_4950), .I1(n8_adj_4938), .I2(n45_adj_4962), 
            .I3(n47392), .O(n48560));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40657_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39930_3_lut (.I0(n48669), .I1(n88), .I2(n25_adj_4951), .I3(GND_net), 
            .O(n47833));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39930_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1829_3_lut (.I0(n531), .I1(n6732), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1830_i4_4_lut (.I0(n532), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4935));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3128_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n35055), 
            .O(n6502)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40763_3_lut (.I0(n4_adj_4935), .I1(n87), .I2(n27_adj_4952), 
            .I3(GND_net), .O(n48666));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40763_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_118[10]), 
            .I2(n15_adj_4574), .I3(n34854), .O(displacement_23__N_25[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3128_12 (.CI(n35055), .I0(n1644), .I1(n90), .CO(n35056));
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n34854), .I0(displacement_23__N_118[10]), 
            .I1(n15_adj_4574), .CO(n34855));
    SB_LUT4 add_3128_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n35054), 
            .O(n6503)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40764_3_lut (.I0(n48666), .I1(n86), .I2(n29_adj_4953), .I3(GND_net), 
            .O(n48667));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40764_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_634_i9_2_lut (.I0(pwm_count[4]), .I1(n872), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4633));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_634_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_118[9]), 
            .I2(n16_adj_4573), .I3(n34853), .O(displacement_23__N_25[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39527_4_lut (.I0(n33_adj_4956), .I1(n31_adj_4955), .I2(n29_adj_4953), 
            .I3(n47434), .O(n47430));
    defparam i39527_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n34853), .I0(displacement_23__N_118[9]), 
            .I1(n16_adj_4573), .CO(n34854));
    SB_CARRY add_3128_11 (.CI(n35054), .I0(n1645), .I1(n91), .CO(n35055));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_118[8]), 
            .I2(n17_adj_4572), .I3(n34852), .O(displacement_23__N_25[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41023_4_lut (.I0(n30_adj_4954), .I1(n10_adj_4940), .I2(n35_adj_4957), 
            .I3(n47428), .O(n48926));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41023_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3128_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n35053), 
            .O(n6504)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_634_i4_3_lut (.I0(n46548), .I1(n875), .I2(pwm_count[1]), 
            .I3(GND_net), .O(n4_adj_4630));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_634_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39932_3_lut (.I0(n48667), .I1(n85), .I2(n31_adj_4955), .I3(GND_net), 
            .O(n47835));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39932_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41139_4_lut (.I0(n47835), .I1(n48926), .I2(n35_adj_4957), 
            .I3(n47430), .O(n49042));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41139_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_634_i8_3_lut (.I0(n6_adj_4631), .I1(n872), .I2(n9_adj_4633), 
            .I3(GND_net), .O(n8_adj_4632));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_634_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41140_3_lut (.I0(n49042), .I1(n82), .I2(n37_adj_4958), .I3(GND_net), 
            .O(n49043));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41140_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41117_3_lut (.I0(n49043), .I1(n81), .I2(n39_adj_4959), .I3(GND_net), 
            .O(n49020));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41117_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39493_4_lut (.I0(n43_adj_4961), .I1(n41_adj_4960), .I2(n39_adj_4959), 
            .I3(n48956), .O(n47396));
    defparam i39493_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i41005_4_lut (.I0(n47833), .I1(n48560), .I2(n45_adj_4962), 
            .I3(n47394), .O(n48908));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41005_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40954_4_lut (.I0(n8_adj_4632), .I1(n4_adj_4630), .I2(n9_adj_4633), 
            .I3(n47071), .O(n48857));   // verilog/motorControl.v(86[28:44])
    defparam i40954_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39938_3_lut (.I0(n49020), .I1(n80), .I2(n41_adj_4960), .I3(GND_net), 
            .O(n47841));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39938_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40955_3_lut (.I0(n48857), .I1(n871), .I2(pwm_count[5]), .I3(GND_net), 
            .O(n48858));   // verilog/motorControl.v(86[28:44])
    defparam i40955_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_15_i1807_3_lut (.I0(n2699), .I1(n6710), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3128_10 (.CI(n35053), .I0(n1646), .I1(n92), .CO(n35054));
    SB_LUT4 add_3128_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n35052), 
            .O(n6505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n34852), .I0(displacement_23__N_118[8]), 
            .I1(n17_adj_4572), .CO(n34853));
    SB_CARRY add_3128_9 (.CI(n35052), .I0(n1647), .I1(n93), .CO(n35053));
    SB_LUT4 add_3128_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n35051), 
            .O(n6506)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41007_4_lut (.I0(n47841), .I1(n48908), .I2(n45_adj_4962), 
            .I3(n47396), .O(n48910));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41007_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40798_3_lut (.I0(n48858), .I1(n870), .I2(pwm_count[6]), .I3(GND_net), 
            .O(n48701));   // verilog/motorControl.v(86[28:44])
    defparam i40798_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i41008_3_lut (.I0(n48910), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41008_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39861_3_lut (.I0(n48701), .I1(n869), .I2(pwm_count[7]), .I3(GND_net), 
            .O(n16_adj_4634));   // verilog/motorControl.v(86[28:44])
    defparam i39861_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i12_4_lut (.I0(n857), .I1(n855), .I2(n865), .I3(n866), .O(n28_adj_4968));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_118[7]), 
            .I2(n18_adj_4571), .I3(n34851), .O(displacement_23__N_25[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3128_8 (.CI(n35051), .I0(n1648), .I1(n94), .CO(n35052));
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n34851), .I0(displacement_23__N_118[7]), 
            .I1(n18_adj_4571), .CO(n34852));
    SB_LUT4 add_3128_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n35050), 
            .O(n6507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_634_i18_3_lut (.I0(n16_adj_4634), .I1(n868), .I2(pwm_count[8]), 
            .I3(GND_net), .O(n2677));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_634_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i10_4_lut (.I0(n861), .I1(n856), .I2(n859), .I3(n860), .O(n26_adj_4969));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n44276), .I1(n28_adj_4968), .I2(n862), .I3(n853), 
            .O(n30_adj_4967));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3128_7 (.CI(n35050), .I0(n1649), .I1(n95), .CO(n35051));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_118[6]), 
            .I2(n19_adj_4570), .I3(n34850), .O(displacement_23__N_25[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut (.I0(n2677), .I1(n864), .I2(n863), .I3(n867), .O(n25_adj_4970));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_15_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4934));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i38945_4_lut (.I0(n31_adj_4738), .I1(n29_adj_4736), .I2(n27_adj_4734), 
            .I3(n25_adj_4732), .O(n46847));
    defparam i38945_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38939_4_lut (.I0(n37_adj_4743), .I1(n35_adj_4741), .I2(n33_adj_4740), 
            .I3(n46847), .O(n46841));
    defparam i38939_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1210_i24_4_lut (.I0(n522), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4731));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_15_LessThan_1210_i32_3_lut (.I0(n30_adj_4737), .I1(n93), 
            .I2(n35_adj_4741), .I3(GND_net), .O(n32_adj_4739));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3128_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n35049), 
            .O(n6508)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3128_6 (.CI(n35049), .I0(n1650), .I1(n96), .CO(n35050));
    SB_LUT4 add_3128_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n35048), 
            .O(n6509)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n34850), .I0(displacement_23__N_118[6]), 
            .I1(n19_adj_4570), .CO(n34851));
    SB_LUT4 div_15_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4930));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3128_5 (.CI(n35048), .I0(n1651), .I1(n97), .CO(n35049));
    SB_LUT4 add_3128_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n35047), 
            .O(n6510)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3128_4 (.CI(n35047), .I0(n1652), .I1(n98), .CO(n35048));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_118[5]), 
            .I2(n20_adj_4569), .I3(n34849), .O(displacement_23__N_25[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4932));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4933));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n531));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n34849), .I0(displacement_23__N_118[5]), 
            .I1(n20_adj_4569), .CO(n34850));
    SB_LUT4 add_3128_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n35046), 
            .O(n6511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4927));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4928));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_118[4]), 
            .I2(n21_adj_4568), .I3(n34848), .O(displacement_23__N_25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4925));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4926));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13014_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n41848), 
            .I3(GND_net), .O(n18298));   // verilog/coms.v(126[12] 289[6])
    defparam i13014_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4916));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4918));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4924));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12748_2_lut_2_lut (.I0(pwm[23]), .I1(pwm[22]), .I2(GND_net), 
            .I3(GND_net), .O(n18032));   // verilog/TinyFPGA_B.v(44[8:13])
    defparam i12748_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_15_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4920));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4922));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4923));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12749_2_lut_2_lut (.I0(pwm[23]), .I1(pwm[21]), .I2(GND_net), 
            .I3(GND_net), .O(n18033));   // verilog/TinyFPGA_B.v(44[8:13])
    defparam i12749_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_15_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4929));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12750_2_lut_2_lut (.I0(pwm[23]), .I1(pwm[20]), .I2(GND_net), 
            .I3(GND_net), .O(n18034));   // verilog/TinyFPGA_B.v(44[8:13])
    defparam i12750_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_15_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39571_4_lut (.I0(n29_adj_4929), .I1(n17_adj_4923), .I2(n15_adj_4922), 
            .I3(n13_adj_4920), .O(n47474));
    defparam i39571_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39608_4_lut (.I0(n11_adj_4918), .I1(n9_adj_4916), .I2(n2719), 
            .I3(n98), .O(n47511));
    defparam i39608_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i40223_4_lut (.I0(n17_adj_4923), .I1(n15_adj_4922), .I2(n13_adj_4920), 
            .I3(n47511), .O(n48126));
    defparam i40223_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40219_4_lut (.I0(n23_adj_4926), .I1(n21_adj_4925), .I2(n19_adj_4924), 
            .I3(n48126), .O(n48122));
    defparam i40219_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_3128_3 (.CI(n35046), .I0(n1653), .I1(n99), .CO(n35047));
    SB_LUT4 i39575_4_lut (.I0(n29_adj_4929), .I1(n27_adj_4928), .I2(n25_adj_4927), 
            .I3(n48122), .O(n47478));
    defparam i39575_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3128_2_lut (.I0(GND_net), .I1(n520), .I2(n558), .I3(VCC_net), 
            .O(n6512)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3128_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3128_2 (.CI(VCC_net), .I0(n520), .I1(n558), .CO(n35046));
    SB_LUT4 add_3127_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n35045), 
            .O(n6488)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3127_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n35044), 
            .O(n6489)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1777_i6_4_lut (.I0(n531), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4914));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3127_11 (.CI(n35044), .I0(n1530), .I1(n91), .CO(n35045));
    SB_LUT4 i40482_3_lut (.I0(n6_adj_4914), .I1(n87), .I2(n29_adj_4929), 
            .I3(GND_net), .O(n48385));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40482_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3127_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n35043), 
            .O(n6490)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(pwm[23]), .I1(hall1), .I2(hall2), .I3(GATES_5__N_3398[5]), 
            .O(n5_adj_4984));   // verilog/TinyFPGA_B.v(44[8:13])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h55fd;
    SB_LUT4 div_15_LessThan_1777_i32_3_lut (.I0(n14_adj_4921), .I1(n83), 
            .I2(n37_adj_4934), .I3(GND_net), .O(n32_adj_4931));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13015_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n41848), 
            .I3(GND_net), .O(n18299));   // verilog/coms.v(126[12] 289[6])
    defparam i13015_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n34848), .I0(displacement_23__N_118[4]), 
            .I1(n21_adj_4568), .CO(n34849));
    SB_LUT4 i13016_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n41848), 
            .I3(GND_net), .O(n18300));   // verilog/coms.v(126[12] 289[6])
    defparam i13016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40483_3_lut (.I0(n48385), .I1(n86), .I2(n31_adj_4930), .I3(GND_net), 
            .O(n48386));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40483_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39562_4_lut (.I0(n35_adj_4933), .I1(n33_adj_4932), .I2(n31_adj_4930), 
            .I3(n47474), .O(n47465));
    defparam i39562_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40956_4_lut (.I0(n32_adj_4931), .I1(n12_adj_4919), .I2(n37_adj_4934), 
            .I3(n47461), .O(n48859));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40956_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39918_3_lut (.I0(n48386), .I1(n85), .I2(n33_adj_4932), .I3(GND_net), 
            .O(n47821));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39918_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13017_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n41848), 
            .I3(GND_net), .O(n18301));   // verilog/coms.v(126[12] 289[6])
    defparam i13017_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3127_10 (.CI(n35043), .I0(n1531), .I1(n92), .CO(n35044));
    SB_LUT4 add_3127_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n35042), 
            .O(n6491)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_118[3]), 
            .I2(n22_adj_4567), .I3(n34847), .O(displacement_23__N_25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3127_9 (.CI(n35042), .I0(n1532), .I1(n93), .CO(n35043));
    SB_LUT4 add_3127_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n35041), 
            .O(n6492)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3127_8 (.CI(n35041), .I0(n1533), .I1(n94), .CO(n35042));
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n34847), .I0(displacement_23__N_118[3]), 
            .I1(n22_adj_4567), .CO(n34848));
    SB_LUT4 add_3127_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n35040), 
            .O(n6493)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40484_3_lut (.I0(n8_adj_4915), .I1(n90), .I2(n23_adj_4926), 
            .I3(GND_net), .O(n48387));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40484_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3127_7 (.CI(n35040), .I0(n1534), .I1(n95), .CO(n35041));
    SB_LUT4 i13018_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n41848), 
            .I3(GND_net), .O(n18302));   // verilog/coms.v(126[12] 289[6])
    defparam i13018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3127_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n35039), 
            .O(n6494)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3127_6 (.CI(n35039), .I0(n1535), .I1(n96), .CO(n35040));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_118[2]), 
            .I2(n23_adj_4566), .I3(n34846), .O(displacement_23__N_25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40485_3_lut (.I0(n48387), .I1(n89), .I2(n25_adj_4927), .I3(GND_net), 
            .O(n48388));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40485_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n34846), .I0(displacement_23__N_118[2]), 
            .I1(n23_adj_4566), .CO(n34847));
    SB_LUT4 i40215_4_lut (.I0(n25_adj_4927), .I1(n23_adj_4926), .I2(n21_adj_4925), 
            .I3(n47492), .O(n48118));
    defparam i40215_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3127_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n35038), 
            .O(n6495)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3127_5 (.CI(n35038), .I0(n1536), .I1(n97), .CO(n35039));
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_118[1]), 
            .I2(n24_adj_4565), .I3(n34845), .O(displacement_23__N_25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n34845), .I0(displacement_23__N_118[1]), 
            .I1(n24_adj_4565), .CO(n34846));
    SB_LUT4 add_3127_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n35037), 
            .O(n6496)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3127_4 (.CI(n35037), .I0(n1537), .I1(n98), .CO(n35038));
    SB_LUT4 add_3127_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n35036), 
            .O(n6497)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13019_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n41848), 
            .I3(GND_net), .O(n18303));   // verilog/coms.v(126[12] 289[6])
    defparam i13019_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3127_3 (.CI(n35036), .I0(n1538), .I1(n99), .CO(n35037));
    SB_LUT4 add_3127_2_lut (.I0(GND_net), .I1(n519), .I2(n558), .I3(VCC_net), 
            .O(n6498)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3127_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40655_3_lut (.I0(n10_adj_4917), .I1(n91), .I2(n21_adj_4925), 
            .I3(GND_net), .O(n48558));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40655_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3127_2 (.CI(VCC_net), .I0(n519), .I1(n558), .CO(n35036));
    SB_LUT4 add_3126_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n35035), 
            .O(n6476)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_118[0]), 
            .I2(n25_adj_4564), .I3(VCC_net), .O(displacement_23__N_25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3126_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n35034), 
            .O(n6477)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_10 (.CI(n35034), .I0(n1413), .I1(n92), .CO(n35035));
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_118[0]), 
            .I1(n25_adj_4564), .CO(n34845));
    SB_LUT4 add_3126_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n35033), 
            .O(n6478)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_9 (.CI(n35033), .I0(n1414), .I1(n93), .CO(n35034));
    SB_LUT4 div_15_LessThan_1210_i36_3_lut (.I0(n28_adj_4735), .I1(n91), 
            .I2(n39_adj_4744), .I3(GND_net), .O(n36_adj_4742));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39916_3_lut (.I0(n48388), .I1(n88), .I2(n27_adj_4928), .I3(GND_net), 
            .O(n47819));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39916_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3126_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n35032), 
            .O(n6479)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_8 (.CI(n35032), .I0(n1415), .I1(n94), .CO(n35033));
    SB_LUT4 add_3126_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n35031), 
            .O(n6480)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_7 (.CI(n35031), .I0(n1416), .I1(n95), .CO(n35032));
    SB_LUT4 add_3126_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n35030), 
            .O(n6481)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_6 (.CI(n35030), .I0(n1417), .I1(n96), .CO(n35031));
    SB_LUT4 add_3126_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n35029), 
            .O(n6482)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40777_4_lut (.I0(n35_adj_4933), .I1(n33_adj_4932), .I2(n31_adj_4930), 
            .I3(n47478), .O(n48680));
    defparam i40777_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3126_5 (.CI(n35029), .I0(n1418), .I1(n97), .CO(n35030));
    SB_LUT4 add_3126_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n35028), 
            .O(n6483)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_4 (.CI(n35028), .I0(n1419), .I1(n98), .CO(n35029));
    SB_LUT4 i41111_4_lut (.I0(n47821), .I1(n48859), .I2(n37_adj_4934), 
            .I3(n47465), .O(n49014));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41111_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13020_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n41848), 
            .I3(GND_net), .O(n18304));   // verilog/coms.v(126[12] 289[6])
    defparam i13020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40781_4_lut (.I0(n47819), .I1(n48558), .I2(n27_adj_4928), 
            .I3(n48118), .O(n48684));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40781_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3126_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n35027), 
            .O(n6484)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3126_3 (.CI(n35027), .I0(n1420), .I1(n99), .CO(n35028));
    SB_LUT4 add_3126_2_lut (.I0(GND_net), .I1(n518), .I2(n558), .I3(VCC_net), 
            .O(n6485)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3126_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41159_4_lut (.I0(n48684), .I1(n49014), .I2(n37_adj_4934), 
            .I3(n48680), .O(n49062));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41159_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41160_3_lut (.I0(n49062), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n49063));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41160_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY add_3126_2 (.CI(VCC_net), .I0(n518), .I1(n558), .CO(n35027));
    SB_LUT4 i41057_3_lut (.I0(n49063), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n48960));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41057_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i40972_3_lut (.I0(n48960), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n48875));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40972_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i41029_4_lut (.I0(n36_adj_4742), .I1(n26_adj_4733), .I2(n39_adj_4744), 
            .I3(n46839), .O(n48932));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41029_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41030_3_lut (.I0(n48932), .I1(n90), .I2(n41_adj_4745), .I3(GND_net), 
            .O(n48933));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41030_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40973_3_lut (.I0(n48875), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n48876));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40973_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1971_4_lut (.I0(n48876), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1971_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i13021_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n41848), 
            .I3(GND_net), .O(n18305));   // verilog/coms.v(126[12] 289[6])
    defparam i13021_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4911));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4913));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4909));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3125_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n35002), 
            .O(n6465)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3125_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n35001), 
            .O(n6466)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_9 (.CI(n35001), .I0(n1293), .I1(n93), .CO(n35002));
    SB_LUT4 add_3125_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n35000), 
            .O(n6467)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_8 (.CI(n35000), .I0(n1294), .I1(n94), .CO(n35001));
    SB_LUT4 div_15_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n530));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3125_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n34999), 
            .O(n6468)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_7 (.CI(n34999), .I0(n1295), .I1(n95), .CO(n35000));
    SB_LUT4 add_3125_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n34998), 
            .O(n6469)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4912));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3125_6 (.CI(n34998), .I0(n1296), .I1(n96), .CO(n34999));
    SB_LUT4 div_15_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4906));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4907));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3125_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n34997), 
            .O(n6470)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_5 (.CI(n34997), .I0(n1297), .I1(n97), .CO(n34998));
    SB_LUT4 div_15_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4904));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3125_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n34996), 
            .O(n6471)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_4 (.CI(n34996), .I0(n1298), .I1(n98), .CO(n34997));
    SB_LUT4 div_15_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4905));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3125_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n34995), 
            .O(n6472)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3125_3 (.CI(n34995), .I0(n1299), .I1(n99), .CO(n34996));
    SB_LUT4 add_3125_2_lut (.I0(GND_net), .I1(n517), .I2(n558), .I3(VCC_net), 
            .O(n6473)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3125_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4903));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3125_2 (.CI(VCC_net), .I0(n517), .I1(n558), .CO(n34995));
    SB_LUT4 add_3124_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n34994), 
            .O(n6455)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3124_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n34993), 
            .O(n6456)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3124_8 (.CI(n34993), .I0(n1170), .I1(n94), .CO(n34994));
    SB_LUT4 div_15_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4894));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4896));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3124_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n34992), 
            .O(n6457)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF color_i18 (.Q(color[17]), .C(clk32MHz), .D(n18034));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i19 (.Q(color[18]), .C(clk32MHz), .D(n18033));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_DFF color_i20 (.Q(color[19]), .C(clk32MHz), .D(n18032));   // verilog/TinyFPGA_B.v(43[10] 50[6])
    SB_LUT4 i40935_3_lut (.I0(n48933), .I1(n89), .I2(n43_adj_4746), .I3(GND_net), 
            .O(n48838));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40935_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3124_7 (.CI(n34992), .I0(n1171), .I1(n95), .CO(n34993));
    SB_LUT4 div_15_i1470_3_lut_3_lut (.I0(n2192), .I1(n6592), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4898));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4900));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1459_3_lut_3_lut (.I0(n2192), .I1(n6581), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1471_3_lut_3_lut (.I0(n2192), .I1(n6593), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1467_3_lut_3_lut (.I0(n2192), .I1(n6589), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4901));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4908));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3124_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n34991), 
            .O(n6458)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3124_6 (.CI(n34991), .I0(n1172), .I1(n96), .CO(n34992));
    SB_LUT4 div_15_i1465_3_lut_3_lut (.I0(n2192), .I1(n6587), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643_adj_4602));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38831_4_lut (.I0(n31_adj_4908), .I1(n19_adj_4901), .I2(n17_adj_4900), 
            .I3(n15_adj_4898), .O(n46733));
    defparam i38831_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39678_4_lut (.I0(n13_adj_4896), .I1(n11_adj_4894), .I2(n2637), 
            .I3(n98), .O(n47581));
    defparam i39678_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 add_3124_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n34990), 
            .O(n6459)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40257_4_lut (.I0(n19_adj_4901), .I1(n17_adj_4900), .I2(n15_adj_4898), 
            .I3(n47581), .O(n48160));
    defparam i40257_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40255_4_lut (.I0(n25_adj_4905), .I1(n23_adj_4904), .I2(n21_adj_4903), 
            .I3(n48160), .O(n48158));
    defparam i40255_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40546_4_lut (.I0(n43_adj_4746), .I1(n41_adj_4745), .I2(n39_adj_4744), 
            .I3(n46841), .O(n48449));
    defparam i40546_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3124_5 (.CI(n34990), .I0(n1173), .I1(n97), .CO(n34991));
    SB_LUT4 add_3124_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n34989), 
            .O(n6460)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3124_4 (.CI(n34989), .I0(n1174), .I1(n98), .CO(n34990));
    SB_LUT4 add_3124_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n34988), 
            .O(n6461)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1475_3_lut_3_lut (.I0(n2192), .I1(n6597), .I2(n525), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38833_4_lut (.I0(n31_adj_4908), .I1(n29_adj_4907), .I2(n27_adj_4906), 
            .I3(n48158), .O(n46735));
    defparam i38833_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3124_3 (.CI(n34988), .I0(n1175), .I1(n99), .CO(n34989));
    SB_LUT4 add_3124_2_lut (.I0(GND_net), .I1(n516), .I2(n558), .I3(VCC_net), 
            .O(n6462)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3124_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_15_i1463_3_lut_3_lut (.I0(n2192), .I1(n6585), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3124_2 (.CI(VCC_net), .I0(n516), .I1(n558), .CO(n34988));
    SB_LUT4 add_3140_25_lut (.I0(n249), .I1(n49780), .I2(n248), .I3(n35333), 
            .O(displacement_23__N_118[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_15_LessThan_1722_i8_4_lut (.I0(n530), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4892));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3140_24_lut (.I0(n393), .I1(n49780), .I2(n392), .I3(n35332), 
            .O(displacement_23__N_118[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_15_i1462_3_lut_3_lut (.I0(n2192), .I1(n6584), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i40709_3_lut (.I0(n8_adj_4892), .I1(n87), .I2(n31_adj_4908), 
            .I3(GND_net), .O(n48612));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40709_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3140_24 (.CI(n35332), .I0(n49780), .I1(n392), .CO(n35333));
    SB_LUT4 div_15_i1461_3_lut_3_lut (.I0(n2192), .I1(n6583), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i40710_3_lut (.I0(n48612), .I1(n86), .I2(n33_adj_4909), .I3(GND_net), 
            .O(n48613));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40710_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1464_3_lut_3_lut (.I0(n2192), .I1(n6586), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3140_23_lut (.I0(n534), .I1(n49780), .I2(n533), .I3(n35331), 
            .O(displacement_23__N_118[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_15_i1460_3_lut_3_lut (.I0(n2192), .I1(n6582), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1474_3_lut_3_lut (.I0(n2192), .I1(n6596), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1472_3_lut_3_lut (.I0(n2192), .I1(n6594), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3140_23 (.CI(n35331), .I0(n49780), .I1(n533), .CO(n35332));
    SB_LUT4 add_3140_22_lut (.I0(n672), .I1(n49780), .I2(n671), .I3(n35330), 
            .O(displacement_23__N_118[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_15_i1473_3_lut_3_lut (.I0(n2192), .I1(n6595), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i34_3_lut (.I0(n16_adj_4899), .I1(n83), 
            .I2(n39_adj_4913), .I3(GND_net), .O(n34_adj_4910));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1469_3_lut_3_lut (.I0(n2192), .I1(n6591), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3140_22 (.CI(n35330), .I0(n49780), .I1(n671), .CO(n35331));
    SB_LUT4 add_3140_21_lut (.I0(n807), .I1(n49780), .I2(n806), .I3(n35329), 
            .O(displacement_23__N_118[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_21 (.CI(n35329), .I0(n49780), .I1(n806), .CO(n35330));
    SB_LUT4 i38821_4_lut (.I0(n37_adj_4912), .I1(n35_adj_4911), .I2(n33_adj_4909), 
            .I3(n46733), .O(n46723));
    defparam i38821_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3140_20_lut (.I0(n939), .I1(n49780), .I2(n938), .I3(n35328), 
            .O(displacement_23__N_118[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_20 (.CI(n35328), .I0(n49780), .I1(n938), .CO(n35329));
    SB_LUT4 add_3140_19_lut (.I0(n1068), .I1(n49780), .I2(n1067), .I3(n35327), 
            .O(displacement_23__N_118[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i41049_4_lut (.I0(n34_adj_4910), .I1(n14_adj_4897), .I2(n39_adj_4913), 
            .I3(n46719), .O(n48952));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41049_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_15_i1468_3_lut_3_lut (.I0(n2192), .I1(n6590), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i40648_3_lut (.I0(n48613), .I1(n85), .I2(n35_adj_4911), .I3(GND_net), 
            .O(n48551));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40648_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1466_3_lut_3_lut (.I0(n2192), .I1(n6588), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3140_19 (.CI(n35327), .I0(n49780), .I1(n1067), .CO(n35328));
    SB_LUT4 add_3140_18_lut (.I0(n1194), .I1(n49780), .I2(n1193), .I3(n35326), 
            .O(displacement_23__N_118[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_18 (.CI(n35326), .I0(n49780), .I1(n1193), .CO(n35327));
    SB_LUT4 add_3140_17_lut (.I0(n1317), .I1(n49780), .I2(n1316), .I3(n35325), 
            .O(displacement_23__N_118[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_17 (.CI(n35325), .I0(n49780), .I1(n1316), .CO(n35326));
    SB_LUT4 i40711_3_lut (.I0(n10_adj_4893), .I1(n90), .I2(n25_adj_4905), 
            .I3(GND_net), .O(n48614));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40711_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40712_3_lut (.I0(n48614), .I1(n89), .I2(n27_adj_4906), .I3(GND_net), 
            .O(n48615));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40712_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3140_16_lut (.I0(n1437), .I1(n49780), .I2(n1436), .I3(n35324), 
            .O(displacement_23__N_118[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i39658_4_lut (.I0(n27_adj_4906), .I1(n25_adj_4905), .I2(n23_adj_4904), 
            .I3(n46759), .O(n47561));
    defparam i39658_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_15_LessThan_1722_i20_3_lut (.I0(n12_adj_4895), .I1(n91), 
            .I2(n23_adj_4904), .I3(GND_net), .O(n20_adj_4902));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40646_3_lut (.I0(n48615), .I1(n88), .I2(n29_adj_4907), .I3(GND_net), 
            .O(n48549));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40646_3_lut.LUT_INIT = 16'h3a3a;
    GND i1 (.Y(GND_net));
    SB_LUT4 i40494_4_lut (.I0(n37_adj_4912), .I1(n35_adj_4911), .I2(n33_adj_4909), 
            .I3(n46735), .O(n48397));
    defparam i40494_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3140_16 (.CI(n35324), .I0(n49780), .I1(n1436), .CO(n35325));
    SB_LUT4 i41145_4_lut (.I0(n48551), .I1(n48952), .I2(n39_adj_4913), 
            .I3(n46723), .O(n49048));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41145_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40603_4_lut (.I0(n32_adj_4739), .I1(n24_adj_4731), .I2(n35_adj_4741), 
            .I3(n46845), .O(n48506));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40603_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40651_4_lut (.I0(n48549), .I1(n20_adj_4902), .I2(n29_adj_4907), 
            .I3(n47561), .O(n48554));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40651_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3140_15_lut (.I0(n1554), .I1(n49780), .I2(n1553), .I3(n35323), 
            .O(displacement_23__N_118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i41167_4_lut (.I0(n48554), .I1(n49048), .I2(n39_adj_4913), 
            .I3(n48397), .O(n49070));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13038_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n41851), 
            .I3(GND_net), .O(n18322));   // verilog/coms.v(126[12] 289[6])
    defparam i13038_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3140_15 (.CI(n35323), .I0(n49780), .I1(n1553), .CO(n35324));
    SB_LUT4 add_3140_14_lut (.I0(n1668), .I1(n49780), .I2(n1667), .I3(n35322), 
            .O(displacement_23__N_118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_14 (.CI(n35322), .I0(n49780), .I1(n1667), .CO(n35323));
    SB_LUT4 add_3140_13_lut (.I0(n1779), .I1(n49780), .I2(n1778), .I3(n35321), 
            .O(displacement_23__N_118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3140_13 (.CI(n35321), .I0(n49780), .I1(n1778), .CO(n35322));
    SB_LUT4 add_3140_12_lut (.I0(n1887), .I1(n49780), .I2(n1886), .I3(n35320), 
            .O(displacement_23__N_118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i41168_3_lut (.I0(n49070), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n49071));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41168_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13178_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[6] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18462));   // verilog/coms.v(126[12] 289[6])
    defparam i13178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i41162_3_lut (.I0(n49071), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n49065));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41162_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i40653_3_lut (.I0(n49065), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n48556));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40653_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13179_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[6] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18463));   // verilog/coms.v(126[12] 289[6])
    defparam i13179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(n48556), .I1(n16672), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'hceef;
    SB_LUT4 i13180_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[5] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18464));   // verilog/coms.v(126[12] 289[6])
    defparam i13180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18426_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[5] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n23694));
    defparam i18426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13182_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[5] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18466));   // verilog/coms.v(126[12] 289[6])
    defparam i13182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4889));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13183_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[5] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18467));   // verilog/coms.v(126[12] 289[6])
    defparam i13183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4891));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13184_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[5] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18468));   // verilog/coms.v(126[12] 289[6])
    defparam i13184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4887));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13185_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[5] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18469));   // verilog/coms.v(126[12] 289[6])
    defparam i13185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n529));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13186_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[5] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18470));   // verilog/coms.v(126[12] 289[6])
    defparam i13186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4884));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4885));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13187_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[5] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18471));   // verilog/coms.v(126[12] 289[6])
    defparam i13187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13188_3_lut (.I0(\PID_CONTROLLER.err_prev [1]), .I1(\PID_CONTROLLER.err [1]), 
            .I2(n43362), .I3(GND_net), .O(n18472));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13189_3_lut (.I0(\PID_CONTROLLER.err_prev [2]), .I1(\PID_CONTROLLER.err [2]), 
            .I2(n43362), .I3(GND_net), .O(n18473));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4890));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13190_3_lut (.I0(\PID_CONTROLLER.err_prev [3]), .I1(\PID_CONTROLLER.err [3]), 
            .I2(n43362), .I3(GND_net), .O(n18474));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13191_3_lut (.I0(\PID_CONTROLLER.err_prev [4]), .I1(\PID_CONTROLLER.err [4]), 
            .I2(n43362), .I3(GND_net), .O(n18475));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4881));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13192_3_lut (.I0(\PID_CONTROLLER.err_prev [5]), .I1(\PID_CONTROLLER.err [5]), 
            .I2(n43362), .I3(GND_net), .O(n18476));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4882));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4883));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13193_3_lut (.I0(\PID_CONTROLLER.err_prev [6]), .I1(\PID_CONTROLLER.err [6]), 
            .I2(n43362), .I3(GND_net), .O(n18477));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13194_3_lut (.I0(\PID_CONTROLLER.err_prev [7]), .I1(\PID_CONTROLLER.err [7]), 
            .I2(n43362), .I3(GND_net), .O(n18478));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13195_3_lut (.I0(\PID_CONTROLLER.err_prev [8]), .I1(\PID_CONTROLLER.err [8]), 
            .I2(n43362), .I3(GND_net), .O(n18479));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4872));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13196_3_lut (.I0(\PID_CONTROLLER.err_prev [9]), .I1(\PID_CONTROLLER.err [9]), 
            .I2(n43362), .I3(GND_net), .O(n18480));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4874));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13197_3_lut (.I0(\PID_CONTROLLER.err_prev [10]), .I1(\PID_CONTROLLER.err [10]), 
            .I2(n43362), .I3(GND_net), .O(n18481));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4876));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4878));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13198_3_lut (.I0(\PID_CONTROLLER.err_prev [11]), .I1(\PID_CONTROLLER.err [11]), 
            .I2(n43362), .I3(GND_net), .O(n18482));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4879));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4886));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13199_3_lut (.I0(\PID_CONTROLLER.err_prev [12]), .I1(\PID_CONTROLLER.err [12]), 
            .I2(n43362), .I3(GND_net), .O(n18483));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13200_3_lut (.I0(\PID_CONTROLLER.err_prev [13]), .I1(\PID_CONTROLLER.err [13]), 
            .I2(n43362), .I3(GND_net), .O(n18484));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38926_4_lut (.I0(n33_adj_4886), .I1(n21_adj_4879), .I2(n19_adj_4878), 
            .I3(n17_adj_4876), .O(n46828));
    defparam i38926_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13201_3_lut (.I0(\PID_CONTROLLER.err_prev [14]), .I1(\PID_CONTROLLER.err [14]), 
            .I2(n43362), .I3(GND_net), .O(n18485));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13201_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39746_4_lut (.I0(n15_adj_4874), .I1(n13_adj_4872), .I2(n2552), 
            .I3(n98), .O(n47649));
    defparam i39746_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i40287_4_lut (.I0(n21_adj_4879), .I1(n19_adj_4878), .I2(n17_adj_4876), 
            .I3(n47649), .O(n48190));
    defparam i40287_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40285_4_lut (.I0(n27_adj_4883), .I1(n25_adj_4882), .I2(n23_adj_4881), 
            .I3(n48190), .O(n48188));
    defparam i40285_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i38928_4_lut (.I0(n33_adj_4886), .I1(n31_adj_4885), .I2(n29_adj_4884), 
            .I3(n48188), .O(n46830));
    defparam i38928_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13202_3_lut (.I0(\PID_CONTROLLER.err_prev [15]), .I1(\PID_CONTROLLER.err [15]), 
            .I2(n43362), .I3(GND_net), .O(n18486));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13203_3_lut (.I0(\PID_CONTROLLER.err_prev [16]), .I1(\PID_CONTROLLER.err [16]), 
            .I2(n43362), .I3(GND_net), .O(n18487));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i10_4_lut (.I0(n529), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4870));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i13204_3_lut (.I0(\PID_CONTROLLER.err_prev [17]), .I1(\PID_CONTROLLER.err [17]), 
            .I2(n43362), .I3(GND_net), .O(n18488));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40715_3_lut (.I0(n10_adj_4870), .I1(n87), .I2(n33_adj_4886), 
            .I3(GND_net), .O(n48618));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40715_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40716_3_lut (.I0(n48618), .I1(n86), .I2(n35_adj_4887), .I3(GND_net), 
            .O(n48619));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40716_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13205_3_lut (.I0(\PID_CONTROLLER.err_prev [18]), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n43362), .I3(GND_net), .O(n18489));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13206_3_lut (.I0(\PID_CONTROLLER.err_prev [19]), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n43362), .I3(GND_net), .O(n18490));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13207_3_lut (.I0(\PID_CONTROLLER.err_prev [20]), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n43362), .I3(GND_net), .O(n18491));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i36_3_lut (.I0(n18_adj_4877), .I1(n83), 
            .I2(n41_adj_4891), .I3(GND_net), .O(n36_adj_4888));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i38910_4_lut (.I0(n39_adj_4890), .I1(n37_adj_4889), .I2(n35_adj_4887), 
            .I3(n46828), .O(n46812));
    defparam i38910_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13208_3_lut (.I0(\PID_CONTROLLER.err_prev [21]), .I1(\PID_CONTROLLER.err [21]), 
            .I2(n43362), .I3(GND_net), .O(n18492));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i41047_4_lut (.I0(n36_adj_4888), .I1(n16_adj_4875), .I2(n41_adj_4891), 
            .I3(n46808), .O(n48950));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41047_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13209_3_lut (.I0(\PID_CONTROLLER.err_prev [22]), .I1(\PID_CONTROLLER.err [22]), 
            .I2(n43362), .I3(GND_net), .O(n18493));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40642_3_lut (.I0(n48619), .I1(n85), .I2(n37_adj_4889), .I3(GND_net), 
            .O(n48545));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40642_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13210_3_lut (.I0(\PID_CONTROLLER.err_prev [23]), .I1(\PID_CONTROLLER.err [23]), 
            .I2(n43362), .I3(GND_net), .O(n18494));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13211_3_lut (.I0(\PID_CONTROLLER.err_prev [31]), .I1(\PID_CONTROLLER.err [31]), 
            .I2(n43362), .I3(GND_net), .O(n18495));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1665_i22_3_lut (.I0(n14_adj_4873), .I1(n91), 
            .I2(n25_adj_4882), .I3(GND_net), .O(n22_adj_4880));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41045_4_lut (.I0(n22_adj_4880), .I1(n12_adj_4871), .I2(n25_adj_4882), 
            .I3(n46849), .O(n48948));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41045_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41046_3_lut (.I0(n48948), .I1(n90), .I2(n27_adj_4883), .I3(GND_net), 
            .O(n48949));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41046_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40919_3_lut (.I0(n48949), .I1(n89), .I2(n29_adj_4884), .I3(GND_net), 
            .O(n48822));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40919_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40542_4_lut (.I0(n39_adj_4890), .I1(n37_adj_4889), .I2(n35_adj_4887), 
            .I3(n46830), .O(n48445));
    defparam i40542_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i41143_4_lut (.I0(n48545), .I1(n48950), .I2(n41_adj_4891), 
            .I3(n46812), .O(n49046));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41143_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40873_3_lut (.I0(n48822), .I1(n88), .I2(n31_adj_4885), .I3(GND_net), 
            .O(n48776));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40873_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41171_4_lut (.I0(n48776), .I1(n49046), .I2(n41_adj_4891), 
            .I3(n48445), .O(n49074));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41172_3_lut (.I0(n49074), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n49075));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41172_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i41164_3_lut (.I0(n49075), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n49067));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41164_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n49067), .I1(n16669), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_i1533_3_lut_3_lut (.I0(n2288), .I1(n6611), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4867));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4865));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1522_3_lut_3_lut (.I0(n2288), .I1(n6600), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4869));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4868));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n528));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4862));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4863));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4859));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1523_3_lut_3_lut (.I0(n2288), .I1(n6601), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4860));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4861));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4850));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4852));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1525_3_lut_3_lut (.I0(n2288), .I1(n6603), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4854));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4856));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4857));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut (.I0(n7_adj_4629), .I1(n5_adj_4628), .I2(n123), .I3(n5_adj_4981), 
            .O(n8_adj_4600));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 div_15_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4864));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1526_3_lut_3_lut (.I0(n2288), .I1(n6604), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1535_3_lut_3_lut (.I0(n2288), .I1(n6613), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i4_4_lut (.I0(n50704), .I1(n8_adj_4600), .I2(n16678), .I3(n2484), 
            .O(n50009));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 div_15_i1532_3_lut_3_lut (.I0(n2288), .I1(n6610), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38994_4_lut (.I0(n35_adj_4864), .I1(n23_adj_4857), .I2(n21_adj_4856), 
            .I3(n19_adj_4854), .O(n46896));
    defparam i38994_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39862_4_lut (.I0(n17_adj_4852), .I1(n15_adj_4850), .I2(n2464), 
            .I3(n98), .O(n47765));
    defparam i39862_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i40313_4_lut (.I0(n23_adj_4857), .I1(n21_adj_4856), .I2(n19_adj_4854), 
            .I3(n47765), .O(n48216));
    defparam i40313_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_15_i1340_3_lut_3_lut (.I0(n1991), .I1(n6559), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i40309_4_lut (.I0(n29_adj_4861), .I1(n27_adj_4860), .I2(n25_adj_4859), 
            .I3(n48216), .O(n48212));
    defparam i40309_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_15_i1331_3_lut_3_lut (.I0(n1991), .I1(n6550), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i39011_4_lut (.I0(n35_adj_4864), .I1(n33_adj_4863), .I2(n31_adj_4862), 
            .I3(n48212), .O(n46913));
    defparam i39011_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1606_i12_4_lut (.I0(n528), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4848));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40721_3_lut (.I0(n12_adj_4848), .I1(n87), .I2(n35_adj_4864), 
            .I3(GND_net), .O(n48624));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40721_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1531_3_lut_3_lut (.I0(n2288), .I1(n6609), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1530_3_lut_3_lut (.I0(n2288), .I1(n6608), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13213_3_lut (.I0(encoder0_position[1]), .I1(n2665), .I2(count_enable), 
            .I3(GND_net), .O(n18497));   // quad.v(35[10] 41[6])
    defparam i13213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_3_lut_adj_1627 (.I0(bit_ctr[3]), .I1(n46631), .I2(n43079), 
            .I3(GND_net), .O(n40128));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1627.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_adj_1628 (.I0(bit_ctr[2]), .I1(n46630), .I2(n43079), 
            .I3(GND_net), .O(n40124));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1628.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1606_i38_3_lut (.I0(n20_adj_4855), .I1(n83), 
            .I2(n43_adj_4869), .I3(GND_net), .O(n38_adj_4866));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1529_3_lut_3_lut (.I0(n2288), .I1(n6607), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_3_lut_adj_1629 (.I0(bit_ctr[1]), .I1(n46629), .I2(n43079), 
            .I3(GND_net), .O(n40120));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1629.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1528_3_lut_3_lut (.I0(n2288), .I1(n6606), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13225_2_lut (.I0(n25520), .I1(n18507), .I2(GND_net), .I3(GND_net), 
            .O(n18509));   // verilog/coms.v(126[12] 289[6])
    defparam i13225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40722_3_lut (.I0(n48624), .I1(n86), .I2(n37_adj_4865), .I3(GND_net), 
            .O(n48625));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40722_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13226_3_lut (.I0(encoder0_position[2]), .I1(n2664), .I2(count_enable), 
            .I3(GND_net), .O(n18510));   // quad.v(35[10] 41[6])
    defparam i13226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38985_4_lut (.I0(n41_adj_4868), .I1(n39_adj_4867), .I2(n37_adj_4865), 
            .I3(n46896), .O(n46887));
    defparam i38985_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4756));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13227_3_lut (.I0(encoder0_position[3]), .I1(n2663), .I2(count_enable), 
            .I3(GND_net), .O(n18511));   // quad.v(35[10] 41[6])
    defparam i13227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4758));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i40719_4_lut (.I0(n38_adj_4866), .I1(n18_adj_4853), .I2(n43_adj_4869), 
            .I3(n46881), .O(n48622));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40719_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13228_3_lut (.I0(encoder0_position[4]), .I1(n2662), .I2(count_enable), 
            .I3(GND_net), .O(n18512));   // quad.v(35[10] 41[6])
    defparam i13228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13229_3_lut (.I0(encoder0_position[5]), .I1(n2661), .I2(count_enable), 
            .I3(GND_net), .O(n18513));   // quad.v(35[10] 41[6])
    defparam i13229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40636_3_lut (.I0(n48625), .I1(n85), .I2(n39_adj_4867), .I3(GND_net), 
            .O(n48539));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40636_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13230_3_lut (.I0(encoder0_position[6]), .I1(n2660), .I2(count_enable), 
            .I3(GND_net), .O(n18514));   // quad.v(35[10] 41[6])
    defparam i13230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13231_3_lut (.I0(encoder0_position[7]), .I1(n2659), .I2(count_enable), 
            .I3(GND_net), .O(n18515));   // quad.v(35[10] 41[6])
    defparam i13231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1524_3_lut_3_lut (.I0(n2288), .I1(n6602), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13232_3_lut (.I0(encoder0_position[8]), .I1(n2658), .I2(count_enable), 
            .I3(GND_net), .O(n18516));   // quad.v(35[10] 41[6])
    defparam i13232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1539_3_lut_3_lut (.I0(n2288), .I1(n6617), .I2(n526), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4692));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4693));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13233_3_lut (.I0(encoder0_position[9]), .I1(n2657), .I2(count_enable), 
            .I3(GND_net), .O(n18517));   // quad.v(35[10] 41[6])
    defparam i13233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4691));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4695));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1606_i24_3_lut (.I0(n16_adj_4851), .I1(n91), 
            .I2(n27_adj_4860), .I3(GND_net), .O(n24_adj_4858));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13234_3_lut (.I0(encoder0_position[10]), .I1(n2656), .I2(count_enable), 
            .I3(GND_net), .O(n18518));   // quad.v(35[10] 41[6])
    defparam i13234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4697));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13235_3_lut (.I0(encoder0_position[11]), .I1(n2655), .I2(count_enable), 
            .I3(GND_net), .O(n18519));   // quad.v(35[10] 41[6])
    defparam i13235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4698));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13236_3_lut (.I0(encoder0_position[12]), .I1(n2654), .I2(count_enable), 
            .I3(GND_net), .O(n18520));   // quad.v(35[10] 41[6])
    defparam i13236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4699));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i41043_4_lut (.I0(n24_adj_4858), .I1(n14_adj_4849), .I2(n27_adj_4860), 
            .I3(n46949), .O(n48946));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41043_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_15_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4702));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13237_3_lut (.I0(encoder0_position[13]), .I1(n2653), .I2(count_enable), 
            .I3(GND_net), .O(n18521));   // quad.v(35[10] 41[6])
    defparam i13237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41044_3_lut (.I0(n48946), .I1(n90), .I2(n29_adj_4861), .I3(GND_net), 
            .O(n48947));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41044_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4703));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13238_3_lut (.I0(encoder0_position[14]), .I1(n2652), .I2(count_enable), 
            .I3(GND_net), .O(n18522));   // quad.v(35[10] 41[6])
    defparam i13238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4704));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4707));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13239_3_lut (.I0(encoder0_position[15]), .I1(n2651), .I2(count_enable), 
            .I3(GND_net), .O(n18523));   // quad.v(35[10] 41[6])
    defparam i13239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4705));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4708));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i40921_3_lut (.I0(n48947), .I1(n89), .I2(n31_adj_4862), .I3(GND_net), 
            .O(n48824));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40921_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4713));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13240_3_lut (.I0(encoder0_position[16]), .I1(n2650), .I2(count_enable), 
            .I3(GND_net), .O(n18524));   // quad.v(35[10] 41[6])
    defparam i13240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40558_4_lut (.I0(n41_adj_4868), .I1(n39_adj_4867), .I2(n37_adj_4865), 
            .I3(n46913), .O(n48461));
    defparam i40558_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_15_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4711));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13241_3_lut (.I0(encoder0_position[17]), .I1(n2649), .I2(count_enable), 
            .I3(GND_net), .O(n18525));   // quad.v(35[10] 41[6])
    defparam i13241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41021_4_lut (.I0(n48539), .I1(n48622), .I2(n43_adj_4869), 
            .I3(n46887), .O(n48924));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41021_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_15_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4714));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4715));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13242_3_lut (.I0(encoder0_position[18]), .I1(n2648), .I2(count_enable), 
            .I3(GND_net), .O(n18526));   // quad.v(35[10] 41[6])
    defparam i13242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4718));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4716));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1534_3_lut_3_lut (.I0(n2288), .I1(n6612), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4719));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1527_3_lut_3_lut (.I0(n2288), .I1(n6605), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13243_3_lut (.I0(encoder0_position[19]), .I1(n2647), .I2(count_enable), 
            .I3(GND_net), .O(n18527));   // quad.v(35[10] 41[6])
    defparam i13243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40871_3_lut (.I0(n48824), .I1(n88), .I2(n33_adj_4863), .I3(GND_net), 
            .O(n48774));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40871_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4724));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13244_3_lut (.I0(encoder0_position[20]), .I1(n2646), .I2(count_enable), 
            .I3(GND_net), .O(n18528));   // quad.v(35[10] 41[6])
    defparam i13244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4722));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4725));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13245_3_lut (.I0(encoder0_position[21]), .I1(n2645), .I2(count_enable), 
            .I3(GND_net), .O(n18529));   // quad.v(35[10] 41[6])
    defparam i13245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4726));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4729));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i41149_4_lut (.I0(n48774), .I1(n48924), .I2(n43_adj_4869), 
            .I3(n48461), .O(n49052));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41149_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_15_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4727));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4730));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13246_3_lut (.I0(encoder0_position[22]), .I1(n2644), .I2(count_enable), 
            .I3(GND_net), .O(n18530));   // quad.v(35[10] 41[6])
    defparam i13246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41150_3_lut (.I0(n49052), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n49053));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41150_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(n49053), .I1(n16666), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4738));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4740));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4736));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13247_3_lut (.I0(encoder0_position[23]), .I1(n2643), .I2(count_enable), 
            .I3(GND_net), .O(n18531));   // quad.v(35[10] 41[6])
    defparam i13247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4743));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4734));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1538_3_lut_3_lut (.I0(n2288), .I1(n6616), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13248_3_lut (.I0(encoder1_position[1]), .I1(n2615), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18532));   // quad.v(35[10] 41[6])
    defparam i13248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13251_2_lut (.I0(n25520), .I1(n18533), .I2(GND_net), .I3(GND_net), 
            .O(n18535));   // verilog/coms.v(126[12] 289[6])
    defparam i13251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_15_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4847));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4845));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1329_3_lut_3_lut (.I0(n1991), .I1(n6548), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13254_2_lut (.I0(n25520), .I1(n18536), .I2(GND_net), .I3(GND_net), 
            .O(n18538));   // verilog/coms.v(126[12] 289[6])
    defparam i13254_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13257_2_lut (.I0(n25520), .I1(n18539), .I2(GND_net), .I3(GND_net), 
            .O(n18541));   // verilog/coms.v(126[12] 289[6])
    defparam i13257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_15_i1537_3_lut_3_lut (.I0(n2288), .I1(n6615), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13260_2_lut (.I0(n25520), .I1(n18542), .I2(GND_net), .I3(GND_net), 
            .O(n18544));   // verilog/coms.v(126[12] 289[6])
    defparam i13260_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13263_2_lut (.I0(n25520), .I1(n18545), .I2(GND_net), .I3(GND_net), 
            .O(n18547));   // verilog/coms.v(126[12] 289[6])
    defparam i13263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13266_2_lut (.I0(n25520), .I1(n18548), .I2(GND_net), .I3(GND_net), 
            .O(n18550));   // verilog/coms.v(126[12] 289[6])
    defparam i13266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_15_i1536_3_lut_3_lut (.I0(n2288), .I1(n6614), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1330_3_lut_3_lut (.I0(n1991), .I1(n6549), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1327_3_lut_3_lut (.I0(n1991), .I1(n6546), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1328_3_lut_3_lut (.I0(n1991), .I1(n6547), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13268_4_lut (.I0(n17802), .I1(state[1]), .I2(state_3__N_248[1]), 
            .I3(n17665), .O(n18552));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13268_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut_adj_1631 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4973));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1631.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_i1339_3_lut_3_lut (.I0(n1991), .I1(n6558), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i4_4_lut_adj_1632 (.I0(n17503), .I1(\data_in_frame[8] [0]), 
            .I2(n41916), .I3(n6), .O(n37561));
    defparam i4_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 i13271_4_lut (.I0(n27708), .I1(r_Clock_Count[1]), .I2(n225), 
            .I3(n17657), .O(n18555));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13271_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i3_4_lut_adj_1633 (.I0(n42432), .I1(n42357), .I2(\data_in_frame[13] [7]), 
            .I3(n42125), .O(n42079));
    defparam i3_4_lut_adj_1633.LUT_INIT = 16'h6996;
    SB_LUT4 div_15_i1337_3_lut_3_lut (.I0(n1991), .I1(n6556), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1338_3_lut_3_lut (.I0(n1991), .I1(n6557), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1634 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42219));
    defparam i1_2_lut_adj_1634.LUT_INIT = 16'h6666;
    SB_LUT4 div_15_i1335_3_lut_3_lut (.I0(n1991), .I1(n6554), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1635 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28_adj_4975));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1635.LUT_INIT = 16'h6666;
    SB_LUT4 i13283_4_lut (.I0(n27708), .I1(r_Clock_Count[5]), .I2(n221), 
            .I3(n17657), .O(n18567));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13283_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_15_i1336_3_lut_3_lut (.I0(n1991), .I1(n6555), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13078_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n41857), .I3(GND_net), .O(n18362));   // verilog/coms.v(126[12] 289[6])
    defparam i13078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13079_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n41857), .I3(GND_net), .O(n18363));   // verilog/coms.v(126[12] 289[6])
    defparam i13079_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40850_3_lut (.I0(n48838), .I1(n88), .I2(n45_adj_4748), .I3(GND_net), 
            .O(n44_adj_4747));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40850_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13080_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n41857), .I3(GND_net), .O(n18364));   // verilog/coms.v(126[12] 289[6])
    defparam i13080_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13290_4_lut (.I0(pwm_23__N_3307), .I1(n471), .I2(PWMLimit[0]), 
            .I3(n387), .O(n18574));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13290_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1636 (.I0(n18575), .I1(n5_adj_4982), .I2(GND_net), 
            .I3(GND_net), .O(n41348));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_1636.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1637 (.I0(n37512), .I1(n42459), .I2(\data_in_frame[14] [1]), 
            .I3(Kp_23__N_679), .O(n42330));
    defparam i3_4_lut_adj_1637.LUT_INIT = 16'h6996;
    SB_LUT4 i13299_3_lut (.I0(n17849), .I1(r_Bit_Index[0]), .I2(n17707), 
            .I3(GND_net), .O(n18583));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13299_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_15_i1334_3_lut_3_lut (.I0(n1991), .I1(n6553), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1638 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42429));
    defparam i1_2_lut_adj_1638.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(\data_in_frame[13] [6]), .I1(n43056), 
            .I2(GND_net), .I3(GND_net), .O(n42125));
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'h9999;
    SB_LUT4 i5_3_lut (.I0(n38230), .I1(\data_in_frame[12] [0]), .I2(n42125), 
            .I3(GND_net), .O(n14_adj_4979));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(n42429), .I1(\data_in_frame[14] [0]), .I2(n17283), 
            .I3(n42330), .O(n15_adj_4978));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13303_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4588), 
            .I3(n16566), .O(n18587));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13303_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13_3_lut_adj_1640 (.I0(bit_ctr[0]), .I1(n46628), .I2(n43079), 
            .I3(GND_net), .O(n40116));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13_3_lut_adj_1640.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1341_3_lut_3_lut (.I0(n1991), .I1(n6560), .I2(n523), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1333_3_lut_3_lut (.I0(n1991), .I1(n6552), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1332_3_lut_3_lut (.I0(n1991), .I1(n6551), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13309_4_lut (.I0(n25520), .I1(byte_transmit_counter[0]), .I2(n2244), 
            .I3(n4497), .O(n18593));   // verilog/coms.v(126[12] 289[6])
    defparam i13309_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i13310_3_lut (.I0(encoder1_position[2]), .I1(n2614), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18594));   // quad.v(35[10] 41[6])
    defparam i13310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13311_3_lut (.I0(encoder1_position[3]), .I1(n2613), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18595));   // quad.v(35[10] 41[6])
    defparam i13311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13312_3_lut (.I0(encoder1_position[4]), .I1(n2612), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18596));   // quad.v(35[10] 41[6])
    defparam i13312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13313_3_lut (.I0(encoder1_position[5]), .I1(n2611), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18597));   // quad.v(35[10] 41[6])
    defparam i13313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13314_3_lut (.I0(encoder1_position[6]), .I1(n2610), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18598));   // quad.v(35[10] 41[6])
    defparam i13314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13315_3_lut (.I0(encoder1_position[7]), .I1(n2609), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18599));   // quad.v(35[10] 41[6])
    defparam i13315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13316_3_lut (.I0(encoder1_position[8]), .I1(n2608), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18600));   // quad.v(35[10] 41[6])
    defparam i13316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13317_3_lut (.I0(encoder1_position[9]), .I1(n2607), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18601));   // quad.v(35[10] 41[6])
    defparam i13317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13318_3_lut (.I0(encoder1_position[10]), .I1(n2606), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18602));   // quad.v(35[10] 41[6])
    defparam i13318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13081_3_lut (.I0(\data_in_frame[12] [3]), .I1(rx_data[3]), 
            .I2(n41857), .I3(GND_net), .O(n18365));   // verilog/coms.v(126[12] 289[6])
    defparam i13081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13319_3_lut (.I0(encoder1_position[11]), .I1(n2605), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18603));   // quad.v(35[10] 41[6])
    defparam i13319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13320_3_lut (.I0(encoder1_position[12]), .I1(n2604), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18604));   // quad.v(35[10] 41[6])
    defparam i13320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13321_3_lut (.I0(encoder1_position[13]), .I1(n2603), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18605));   // quad.v(35[10] 41[6])
    defparam i13321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13322_3_lut (.I0(encoder1_position[14]), .I1(n2602), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18606));   // quad.v(35[10] 41[6])
    defparam i13322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13082_3_lut (.I0(\data_in_frame[12] [4]), .I1(rx_data[4]), 
            .I2(n41857), .I3(GND_net), .O(n18366));   // verilog/coms.v(126[12] 289[6])
    defparam i13082_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13323_3_lut (.I0(encoder1_position[15]), .I1(n2601), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18607));   // quad.v(35[10] 41[6])
    defparam i13323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13324_3_lut (.I0(encoder1_position[16]), .I1(n2600), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18608));   // quad.v(35[10] 41[6])
    defparam i13324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13083_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n41857), .I3(GND_net), .O(n18367));   // verilog/coms.v(126[12] 289[6])
    defparam i13083_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13325_3_lut (.I0(encoder1_position[17]), .I1(n2599), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18609));   // quad.v(35[10] 41[6])
    defparam i13325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13326_3_lut (.I0(encoder1_position[18]), .I1(n2598), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18610));   // quad.v(35[10] 41[6])
    defparam i13326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13327_3_lut (.I0(encoder1_position[19]), .I1(n2597), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18611));   // quad.v(35[10] 41[6])
    defparam i13327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13328_3_lut (.I0(encoder1_position[20]), .I1(n2596), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18612));   // quad.v(35[10] 41[6])
    defparam i13328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13329_3_lut (.I0(encoder1_position[21]), .I1(n2595), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18613));   // quad.v(35[10] 41[6])
    defparam i13329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13330_3_lut (.I0(encoder1_position[22]), .I1(n2594), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18614));   // quad.v(35[10] 41[6])
    defparam i13330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13331_3_lut (.I0(encoder1_position[23]), .I1(n2593), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n18615));   // quad.v(35[10] 41[6])
    defparam i13331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13332_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n44088), 
            .I3(GND_net), .O(n18616));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13084_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n41857), .I3(GND_net), .O(n18368));   // verilog/coms.v(126[12] 289[6])
    defparam i13084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13334_3_lut (.I0(quadA_debounced_adj_4589), .I1(reg_B_adj_5037[1]), 
            .I2(n43352), .I3(GND_net), .O(n18618));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13334_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39515_4_lut (.I0(n17574), .I1(n4_adj_4983), .I2(n29), .I3(state[0]), 
            .O(n46660));   // verilog/neopixel.v(35[12] 117[6])
    defparam i39515_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n16614), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 i18_4_lut (.I0(n46660), .I1(n43650), .I2(state[1]), .I3(start), 
            .O(n40242));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i12607_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n16432), 
            .I3(n25329), .O(n17891));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12607_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 i12608_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n25329), 
            .I3(n16566), .O(n17892));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12608_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13338_4_lut (.I0(pwm_23__N_3307), .I1(n470), .I2(PWMLimit[1]), 
            .I3(n387), .O(n18622));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13338_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12609_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n16432), 
            .I3(n4_adj_4596), .O(n17893));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13339_4_lut (.I0(pwm_23__N_3307), .I1(n469), .I2(PWMLimit[2]), 
            .I3(n387), .O(n18623));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13339_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13340_4_lut (.I0(pwm_23__N_3307), .I1(n468), .I2(PWMLimit[3]), 
            .I3(n387), .O(n18624));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13340_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13342_4_lut (.I0(pwm_23__N_3307), .I1(n466), .I2(PWMLimit[5]), 
            .I3(n387), .O(n18626));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13342_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12610_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4596), 
            .I3(n16566), .O(n17894));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12610_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12611_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n16432), 
            .I3(n4_adj_4592), .O(n17895));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13344_4_lut (.I0(pwm_23__N_3307), .I1(n464), .I2(PWMLimit[7]), 
            .I3(n387), .O(n18628));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13344_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13345_4_lut (.I0(pwm_23__N_3307), .I1(n463), .I2(PWMLimit[8]), 
            .I3(n387), .O(n18629));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13345_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13346_4_lut (.I0(pwm_23__N_3307), .I1(n462), .I2(PWMLimit[9]), 
            .I3(n387), .O(n18630));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13346_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12612_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4592), 
            .I3(n16566), .O(n17896));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12612_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13348_4_lut (.I0(pwm_23__N_3307), .I1(n460), .I2(PWMLimit[11]), 
            .I3(n387), .O(n18632));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13348_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13349_4_lut (.I0(pwm_23__N_3307), .I1(n459), .I2(PWMLimit[12]), 
            .I3(n387), .O(n18633));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13349_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13351_4_lut (.I0(pwm_23__N_3307), .I1(n457), .I2(PWMLimit[14]), 
            .I3(n387), .O(n18635));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13351_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13352_4_lut (.I0(pwm_23__N_3307), .I1(n456), .I2(PWMLimit[15]), 
            .I3(n387), .O(n18636));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13352_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13353_4_lut (.I0(pwm_23__N_3307), .I1(n455), .I2(PWMLimit[16]), 
            .I3(n387), .O(n18637));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13353_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12613_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n16432), 
            .I3(n4_adj_4588), .O(n17897));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12613_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12674_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17958));   // verilog/coms.v(126[12] 289[6])
    defparam i12674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12675_3_lut (.I0(Kp[0]), .I1(\data_in_frame[2] [0]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n17959));   // verilog/coms.v(126[12] 289[6])
    defparam i12675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12676_3_lut (.I0(Ki[0]), .I1(\data_in_frame[3] [0]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n17960));   // verilog/coms.v(126[12] 289[6])
    defparam i12676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13355_4_lut (.I0(pwm_23__N_3307), .I1(n453), .I2(PWMLimit[18]), 
            .I3(n387), .O(n18639));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13355_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12677_3_lut (.I0(Kd[0]), .I1(\data_in_frame[4] [0]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n17961));   // verilog/coms.v(126[12] 289[6])
    defparam i12677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13357_4_lut (.I0(pwm_23__N_3307), .I1(n451), .I2(PWMLimit[20]), 
            .I3(n387), .O(n18641));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13357_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12678_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[19] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17962));   // verilog/coms.v(126[12] 289[6])
    defparam i12678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13358_4_lut (.I0(pwm_23__N_3307), .I1(n450), .I2(PWMLimit[21]), 
            .I3(n387), .O(n18642));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13358_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12679_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17963));   // verilog/coms.v(126[12] 289[6])
    defparam i12679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12681_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17965));   // verilog/coms.v(126[12] 289[6])
    defparam i12681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13359_4_lut (.I0(pwm_23__N_3307), .I1(n449), .I2(PWMLimit[22]), 
            .I3(n387), .O(n18643));   // verilog/motorControl.v(38[14] 59[8])
    defparam i13359_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i12682_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[7] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17966));   // verilog/coms.v(126[12] 289[6])
    defparam i12682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12683_3_lut (.I0(\PID_CONTROLLER.err_prev [0]), .I1(\PID_CONTROLLER.err [0]), 
            .I2(n43362), .I3(GND_net), .O(n17967));   // verilog/motorControl.v(38[14] 59[8])
    defparam i12683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34694_2_lut (.I0(n16683), .I1(n740), .I2(GND_net), .I3(GND_net), 
            .O(n42577));
    defparam i34694_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21_2_lut (.I0(pwm_23__N_3310[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4608));   // verilog/motorControl.v(32[23:29])
    defparam i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16_2_lut_adj_1641 (.I0(pwm_23__N_3310[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4609));   // verilog/motorControl.v(32[23:29])
    defparam i16_2_lut_adj_1641.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1642 (.I0(n16680), .I1(n2484), .I2(n2857), .I3(n42577), 
            .O(n8_adj_4985));
    defparam i3_4_lut_adj_1642.LUT_INIT = 16'hcdff;
    SB_LUT4 i2_4_lut_adj_1643 (.I0(n42610), .I1(n16687), .I2(n19921), 
            .I3(n42696), .O(n7_adj_4986));
    defparam i2_4_lut_adj_1643.LUT_INIT = 16'h7577;
    SB_LUT4 i1_4_lut_adj_1644 (.I0(\FRAME_MATCHER.state [0]), .I1(n7_adj_4986), 
            .I2(n14246), .I3(n8_adj_4985), .O(n16_adj_4977));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1644.LUT_INIT = 16'haf8c;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(n16563), .I1(n16_adj_4977), .I2(n16675), 
            .I3(\FRAME_MATCHER.state [3]), .O(n40968));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'hcdcc;
    SB_LUT4 i12685_3_lut (.I0(encoder0_position[0]), .I1(n2666), .I2(count_enable), 
            .I3(GND_net), .O(n17969));   // quad.v(35[10] 41[6])
    defparam i12685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12686_3_lut (.I0(encoder1_position[0]), .I1(n2616), .I2(count_enable_adj_4591), 
            .I3(GND_net), .O(n17970));   // quad.v(35[10] 41[6])
    defparam i12686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12687_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n44088), 
            .I3(GND_net), .O(n17971));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12687_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12689_3_lut (.I0(quadB_debounced_adj_4590), .I1(reg_B_adj_5037[0]), 
            .I2(n43352), .I3(GND_net), .O(n17973));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12689_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12690_3_lut (.I0(tx_o), .I1(n3_adj_4971), .I2(r_SM_Main_adj_5024[2]), 
            .I3(GND_net), .O(n17974));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12690_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4843));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12699_3_lut (.I0(setpoint[0]), .I1(n4446), .I2(n43448), .I3(GND_net), 
            .O(n17983));   // verilog/coms.v(126[12] 289[6])
    defparam i12699_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12700_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n35_adj_4966), .I3(GND_net), .O(n17984));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12700_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12707_3_lut (.I0(deadband[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17991));   // verilog/coms.v(126[12] 289[6])
    defparam i12707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12708_3_lut (.I0(deadband[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17992));   // verilog/coms.v(126[12] 289[6])
    defparam i12708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n527));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12709_3_lut (.I0(deadband[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17993));   // verilog/coms.v(126[12] 289[6])
    defparam i12709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12710_3_lut (.I0(deadband[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17994));   // verilog/coms.v(126[12] 289[6])
    defparam i12710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18666_3_lut (.I0(deadband[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17995));
    defparam i18666_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12712_3_lut (.I0(deadband[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17996));   // verilog/coms.v(126[12] 289[6])
    defparam i12712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18421_3_lut (.I0(deadband[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17997));
    defparam i18421_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12714_3_lut (.I0(deadband[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17998));   // verilog/coms.v(126[12] 289[6])
    defparam i12714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12715_3_lut (.I0(deadband[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17999));   // verilog/coms.v(126[12] 289[6])
    defparam i12715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12716_3_lut (.I0(deadband[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18000));   // verilog/coms.v(126[12] 289[6])
    defparam i12716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17897_3_lut (.I0(deadband[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18001));
    defparam i17897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4846));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12718_3_lut (.I0(deadband[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18002));   // verilog/coms.v(126[12] 289[6])
    defparam i12718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4840));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4841));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4837));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4838));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4839));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12719_3_lut (.I0(deadband[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18003));   // verilog/coms.v(126[12] 289[6])
    defparam i12719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17625_3_lut (.I0(deadband[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18004));
    defparam i17625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4828));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12721_3_lut (.I0(deadband[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18005));   // verilog/coms.v(126[12] 289[6])
    defparam i12721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12722_3_lut (.I0(deadband[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18006));   // verilog/coms.v(126[12] 289[6])
    defparam i12722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12723_3_lut (.I0(deadband[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18007));   // verilog/coms.v(126[12] 289[6])
    defparam i12723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17275_3_lut (.I0(deadband[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18008));
    defparam i17275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12725_3_lut (.I0(deadband[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18009));   // verilog/coms.v(126[12] 289[6])
    defparam i12725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17157_3_lut (.I0(deadband[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18010));
    defparam i17157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12727_3_lut (.I0(deadband[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18011));   // verilog/coms.v(126[12] 289[6])
    defparam i12727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12728_3_lut (.I0(deadband[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18012));   // verilog/coms.v(126[12] 289[6])
    defparam i12728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12729_3_lut (.I0(deadband[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18013));   // verilog/coms.v(126[12] 289[6])
    defparam i12729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12754_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18038));   // verilog/coms.v(126[12] 289[6])
    defparam i12754_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12755_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18039));   // verilog/coms.v(126[12] 289[6])
    defparam i12755_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12756_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18040));   // verilog/coms.v(126[12] 289[6])
    defparam i12756_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12757_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18041));   // verilog/coms.v(126[12] 289[6])
    defparam i12757_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4830));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12758_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18042));   // verilog/coms.v(126[12] 289[6])
    defparam i12758_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12759_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18043));   // verilog/coms.v(126[12] 289[6])
    defparam i12759_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12760_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18044));   // verilog/coms.v(126[12] 289[6])
    defparam i12760_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12761_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18045));   // verilog/coms.v(126[12] 289[6])
    defparam i12761_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12762_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18046));   // verilog/coms.v(126[12] 289[6])
    defparam i12762_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12763_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18047));   // verilog/coms.v(126[12] 289[6])
    defparam i12763_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12764_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18048));   // verilog/coms.v(126[12] 289[6])
    defparam i12764_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12765_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18049));   // verilog/coms.v(126[12] 289[6])
    defparam i12765_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12766_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18050));   // verilog/coms.v(126[12] 289[6])
    defparam i12766_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12767_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18051));   // verilog/coms.v(126[12] 289[6])
    defparam i12767_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12768_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18052));   // verilog/coms.v(126[12] 289[6])
    defparam i12768_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12769_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18053));   // verilog/coms.v(126[12] 289[6])
    defparam i12769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4832));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12770_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18054));   // verilog/coms.v(126[12] 289[6])
    defparam i12770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12771_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18055));   // verilog/coms.v(126[12] 289[6])
    defparam i12771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4834));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12772_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18056));   // verilog/coms.v(126[12] 289[6])
    defparam i12772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4835));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4842));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39093_4_lut (.I0(n37_adj_4842), .I1(n25_adj_4835), .I2(n23_adj_4834), 
            .I3(n21_adj_4832), .O(n46995));
    defparam i39093_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39941_4_lut (.I0(n19_adj_4830), .I1(n17_adj_4828), .I2(n2373), 
            .I3(n98), .O(n47844));
    defparam i39941_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i12773_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18057));   // verilog/coms.v(126[12] 289[6])
    defparam i12773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40342_4_lut (.I0(n25_adj_4835), .I1(n23_adj_4834), .I2(n21_adj_4832), 
            .I3(n47844), .O(n48245));
    defparam i40342_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40333_4_lut (.I0(n31_adj_4839), .I1(n29_adj_4838), .I2(n27_adj_4837), 
            .I3(n48245), .O(n48236));
    defparam i40333_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39098_4_lut (.I0(n37_adj_4842), .I1(n35_adj_4841), .I2(n33_adj_4840), 
            .I3(n48236), .O(n47000));
    defparam i39098_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_LessThan_1545_i14_4_lut (.I0(n527), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4826));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i12774_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18058));   // verilog/coms.v(126[12] 289[6])
    defparam i12774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12775_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18059));   // verilog/coms.v(126[12] 289[6])
    defparam i12775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12776_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18060));   // verilog/coms.v(126[12] 289[6])
    defparam i12776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12777_3_lut (.I0(Kp[1]), .I1(\data_in_frame[2] [1]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18061));   // verilog/coms.v(126[12] 289[6])
    defparam i12777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40725_3_lut (.I0(n14_adj_4826), .I1(n87), .I2(n37_adj_4842), 
            .I3(GND_net), .O(n48628));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40725_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12778_3_lut (.I0(Kp[2]), .I1(\data_in_frame[2] [2]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18062));   // verilog/coms.v(126[12] 289[6])
    defparam i12778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12779_3_lut (.I0(Kp[3]), .I1(\data_in_frame[2] [3]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18063));   // verilog/coms.v(126[12] 289[6])
    defparam i12779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12780_3_lut (.I0(Kp[4]), .I1(\data_in_frame[2] [4]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18064));   // verilog/coms.v(126[12] 289[6])
    defparam i12780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12781_3_lut (.I0(Kp[5]), .I1(\data_in_frame[2] [5]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18065));   // verilog/coms.v(126[12] 289[6])
    defparam i12781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12782_3_lut (.I0(Kp[6]), .I1(\data_in_frame[2] [6]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18066));   // verilog/coms.v(126[12] 289[6])
    defparam i12782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12783_3_lut (.I0(Kp[7]), .I1(\data_in_frame[2] [7]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18067));   // verilog/coms.v(126[12] 289[6])
    defparam i12783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12784_3_lut (.I0(Ki[1]), .I1(\data_in_frame[3] [1]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18068));   // verilog/coms.v(126[12] 289[6])
    defparam i12784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40726_3_lut (.I0(n48628), .I1(n86), .I2(n39_adj_4843), .I3(GND_net), 
            .O(n48629));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40726_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12785_3_lut (.I0(Ki[2]), .I1(\data_in_frame[3] [2]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18069));   // verilog/coms.v(126[12] 289[6])
    defparam i12785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i40_3_lut (.I0(n22_adj_4833), .I1(n83), 
            .I2(n45_adj_4847), .I3(GND_net), .O(n40_adj_4844));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39078_4_lut (.I0(n43_adj_4846), .I1(n41_adj_4845), .I2(n39_adj_4843), 
            .I3(n46995), .O(n46980));
    defparam i39078_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40344_4_lut (.I0(n40_adj_4844), .I1(n20_adj_4831), .I2(n45_adj_4847), 
            .I3(n46971), .O(n48247));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40344_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12786_3_lut (.I0(Ki[3]), .I1(\data_in_frame[3] [3]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18070));   // verilog/coms.v(126[12] 289[6])
    defparam i12786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12787_3_lut (.I0(Ki[4]), .I1(\data_in_frame[3] [4]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18071));   // verilog/coms.v(126[12] 289[6])
    defparam i12787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12788_3_lut (.I0(Ki[5]), .I1(\data_in_frame[3] [5]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18072));   // verilog/coms.v(126[12] 289[6])
    defparam i12788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12789_3_lut (.I0(Ki[6]), .I1(\data_in_frame[3] [6]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18073));   // verilog/coms.v(126[12] 289[6])
    defparam i12789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40632_3_lut (.I0(n48629), .I1(n85), .I2(n41_adj_4845), .I3(GND_net), 
            .O(n48535));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40632_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12790_3_lut (.I0(Ki[7]), .I1(\data_in_frame[3] [7]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18074));   // verilog/coms.v(126[12] 289[6])
    defparam i12790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12791_3_lut (.I0(Kd[1]), .I1(\data_in_frame[4] [1]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18075));   // verilog/coms.v(126[12] 289[6])
    defparam i12791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12792_3_lut (.I0(Kd[2]), .I1(\data_in_frame[4] [2]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18076));   // verilog/coms.v(126[12] 289[6])
    defparam i12792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12793_3_lut (.I0(Kd[3]), .I1(\data_in_frame[4] [3]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18077));   // verilog/coms.v(126[12] 289[6])
    defparam i12793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12794_3_lut (.I0(Kd[4]), .I1(\data_in_frame[4] [4]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18078));   // verilog/coms.v(126[12] 289[6])
    defparam i12794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12795_3_lut (.I0(Kd[5]), .I1(\data_in_frame[4] [5]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18079));   // verilog/coms.v(126[12] 289[6])
    defparam i12795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12796_3_lut (.I0(Kd[6]), .I1(\data_in_frame[4] [6]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18080));   // verilog/coms.v(126[12] 289[6])
    defparam i12796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12797_3_lut (.I0(Kd[7]), .I1(\data_in_frame[4] [7]), .I2(n3_adj_4597), 
            .I3(GND_net), .O(n18081));   // verilog/coms.v(126[12] 289[6])
    defparam i12797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12798_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[19] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18082));   // verilog/coms.v(126[12] 289[6])
    defparam i12798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1545_i26_3_lut (.I0(n18_adj_4829), .I1(n91), 
            .I2(n29_adj_4838), .I3(GND_net), .O(n26_adj_4836));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12799_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[19] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18083));   // verilog/coms.v(126[12] 289[6])
    defparam i12799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12800_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[19] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18084));   // verilog/coms.v(126[12] 289[6])
    defparam i12800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12801_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[19] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18085));   // verilog/coms.v(126[12] 289[6])
    defparam i12801_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12802_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[19] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18086));   // verilog/coms.v(126[12] 289[6])
    defparam i12802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i41041_4_lut (.I0(n26_adj_4836), .I1(n16_adj_4827), .I2(n29_adj_4838), 
            .I3(n47019), .O(n48944));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41041_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12803_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[19] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18087));   // verilog/coms.v(126[12] 289[6])
    defparam i12803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i41042_3_lut (.I0(n48944), .I1(n90), .I2(n31_adj_4839), .I3(GND_net), 
            .O(n48945));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41042_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12804_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[19] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18088));   // verilog/coms.v(126[12] 289[6])
    defparam i12804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12805_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[18] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18089));   // verilog/coms.v(126[12] 289[6])
    defparam i12805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12806_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[18] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18090));   // verilog/coms.v(126[12] 289[6])
    defparam i12806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12807_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[18] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18091));   // verilog/coms.v(126[12] 289[6])
    defparam i12807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12808_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[18] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18092));   // verilog/coms.v(126[12] 289[6])
    defparam i12808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12809_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[18] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18093));   // verilog/coms.v(126[12] 289[6])
    defparam i12809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12810_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[18] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18094));   // verilog/coms.v(126[12] 289[6])
    defparam i12810_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12811_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[18] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18095));   // verilog/coms.v(126[12] 289[6])
    defparam i12811_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40923_3_lut (.I0(n48945), .I1(n89), .I2(n33_adj_4840), .I3(GND_net), 
            .O(n48826));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40923_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12812_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[18] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18096));   // verilog/coms.v(126[12] 289[6])
    defparam i12812_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12813_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[17] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18097));   // verilog/coms.v(126[12] 289[6])
    defparam i12813_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12814_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[17] [1]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18098));   // verilog/coms.v(126[12] 289[6])
    defparam i12814_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12815_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[17] [2]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18099));   // verilog/coms.v(126[12] 289[6])
    defparam i12815_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12816_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[17] [3]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18100));   // verilog/coms.v(126[12] 289[6])
    defparam i12816_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12817_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[17] [4]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18101));   // verilog/coms.v(126[12] 289[6])
    defparam i12817_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12818_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[17] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18102));   // verilog/coms.v(126[12] 289[6])
    defparam i12818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12819_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[17] [6]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18103));   // verilog/coms.v(126[12] 289[6])
    defparam i12819_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40577_4_lut (.I0(n43_adj_4846), .I1(n41_adj_4845), .I2(n39_adj_4843), 
            .I3(n47000), .O(n48480));
    defparam i40577_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i40867_4_lut (.I0(n48535), .I1(n48247), .I2(n45_adj_4847), 
            .I3(n46980), .O(n48770));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40867_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12820_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[17] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18104));   // verilog/coms.v(126[12] 289[6])
    defparam i12820_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12821_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18105));   // verilog/coms.v(126[12] 289[6])
    defparam i12821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12822_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18106));   // verilog/coms.v(126[12] 289[6])
    defparam i12822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[0]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_51[0]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12823_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18107));   // verilog/coms.v(126[12] 289[6])
    defparam i12823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12824_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18108));   // verilog/coms.v(126[12] 289[6])
    defparam i12824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12825_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18109));   // verilog/coms.v(126[12] 289[6])
    defparam i12825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40866_3_lut (.I0(n48826), .I1(n88), .I2(n35_adj_4841), .I3(GND_net), 
            .O(n48769));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40866_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_28_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[1]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_51[1]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12826_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18110));   // verilog/coms.v(126[12] 289[6])
    defparam i12826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12827_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18111));   // verilog/coms.v(126[12] 289[6])
    defparam i12827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12828_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18112));   // verilog/coms.v(126[12] 289[6])
    defparam i12828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12829_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18113));   // verilog/coms.v(126[12] 289[6])
    defparam i12829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12830_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18114));   // verilog/coms.v(126[12] 289[6])
    defparam i12830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12831_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18115));   // verilog/coms.v(126[12] 289[6])
    defparam i12831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12832_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18116));   // verilog/coms.v(126[12] 289[6])
    defparam i12832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12833_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18117));   // verilog/coms.v(126[12] 289[6])
    defparam i12833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12834_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18118));   // verilog/coms.v(126[12] 289[6])
    defparam i12834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12835_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18119));   // verilog/coms.v(126[12] 289[6])
    defparam i12835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12836_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18120));   // verilog/coms.v(126[12] 289[6])
    defparam i12836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12837_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18121));   // verilog/coms.v(126[12] 289[6])
    defparam i12837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40869_4_lut (.I0(n48769), .I1(n48770), .I2(n45_adj_4847), 
            .I3(n48480), .O(n48772));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40869_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12838_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18122));   // verilog/coms.v(126[12] 289[6])
    defparam i12838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12839_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18123));   // verilog/coms.v(126[12] 289[6])
    defparam i12839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12840_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18124));   // verilog/coms.v(126[12] 289[6])
    defparam i12840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12841_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18125));   // verilog/coms.v(126[12] 289[6])
    defparam i12841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[2]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n48772), .I1(n16663), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hceef;
    SB_LUT4 mux_27_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_51[2]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13164_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n18448));   // verilog/coms.v(126[12] 289[6])
    defparam i13164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_28_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[3]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_51[3]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12842_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18126));   // verilog/coms.v(126[12] 289[6])
    defparam i12842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12843_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18127));   // verilog/coms.v(126[12] 289[6])
    defparam i12843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12844_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18128));   // verilog/coms.v(126[12] 289[6])
    defparam i12844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12845_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18129));   // verilog/coms.v(126[12] 289[6])
    defparam i12845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12846_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18130));   // verilog/coms.v(126[12] 289[6])
    defparam i12846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12847_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18131));   // verilog/coms.v(126[12] 289[6])
    defparam i12847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12848_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18132));   // verilog/coms.v(126[12] 289[6])
    defparam i12848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12849_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18133));   // verilog/coms.v(126[12] 289[6])
    defparam i12849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12850_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18134));   // verilog/coms.v(126[12] 289[6])
    defparam i12850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12851_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18135));   // verilog/coms.v(126[12] 289[6])
    defparam i12851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[4]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_51[4]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[5]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_51[5]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n16550), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_4599));   // verilog/TinyFPGA_B.v(155[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12855_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n14276), .I3(GND_net), .O(n18139));   // verilog/coms.v(126[12] 289[6])
    defparam i12855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[6]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_51[6]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1647 (.I0(control_mode[0]), .I1(n16550), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4560));   // verilog/TinyFPGA_B.v(155[5:22])
    defparam i1_2_lut_3_lut_adj_1647.LUT_INIT = 16'hefef;
    SB_LUT4 i12856_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n14276), .I3(GND_net), .O(n18140));   // verilog/coms.v(126[12] 289[6])
    defparam i12856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13102_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n41860), .I3(GND_net), .O(n18386));   // verilog/coms.v(126[12] 289[6])
    defparam i13102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13103_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n41860), .I3(GND_net), .O(n18387));   // verilog/coms.v(126[12] 289[6])
    defparam i13103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_28_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[7]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_51[7]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1595_3_lut_3_lut (.I0(n2381), .I1(n6632), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[8]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_51[8]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1583_3_lut_3_lut (.I0(n2381), .I1(n6620), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13104_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n41860), .I3(GND_net), .O(n18388));   // verilog/coms.v(126[12] 289[6])
    defparam i13104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12857_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n14276), .I3(GND_net), .O(n18141));   // verilog/coms.v(126[12] 289[6])
    defparam i12857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1584_3_lut_3_lut (.I0(n2381), .I1(n6621), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[9]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_51[9]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1587_3_lut_3_lut (.I0(n2381), .I1(n6624), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[10]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_51[10]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1588_3_lut_3_lut (.I0(n2381), .I1(n6625), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[11]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_51[11]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1585_3_lut_3_lut (.I0(n2381), .I1(n6622), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[12]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_51[12]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1586_3_lut_3_lut (.I0(n2381), .I1(n6623), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1601_3_lut_3_lut (.I0(n2381), .I1(n6638), .I2(n527), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[13]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_51[13]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1597_3_lut_3_lut (.I0(n2381), .I1(n6634), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[14]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_51[14]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1598_3_lut_3_lut (.I0(n2381), .I1(n6635), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[15]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_51[15]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1594_3_lut_3_lut (.I0(n2381), .I1(n6631), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[16]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_51[16]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1593_3_lut_3_lut (.I0(n2381), .I1(n6630), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1592_3_lut_3_lut (.I0(n2381), .I1(n6629), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12858_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n14276), .I3(GND_net), .O(n18142));   // verilog/coms.v(126[12] 289[6])
    defparam i12858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[17]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_51[17]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1591_3_lut_3_lut (.I0(n2381), .I1(n6628), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[18]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_51[18]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1590_3_lut_3_lut (.I0(n2381), .I1(n6627), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[19]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_51[19]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1596_3_lut_3_lut (.I0(n2381), .I1(n6633), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[20]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_51[20]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1589_3_lut_3_lut (.I0(n2381), .I1(n6626), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[21]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_51[21]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1600_3_lut_3_lut (.I0(n2381), .I1(n6637), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_28_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[22]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_51[22]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1599_3_lut_3_lut (.I0(n2381), .I1(n6636), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i4_4_lut_adj_1648 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4601));   // verilog/TinyFPGA_B.v(155[5:22])
    defparam i4_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1649 (.I0(control_mode[6]), .I1(n10_adj_4601), 
            .I2(control_mode[2]), .I3(GND_net), .O(n16550));   // verilog/TinyFPGA_B.v(155[5:22])
    defparam i5_3_lut_adj_1649.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n16550), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(156[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_28_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_4560), .O(motor_state_23__N_51[23]));   // verilog/TinyFPGA_B.v(156[5] 159[10])
    defparam mux_28_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_27_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_51[23]), 
            .I2(n15_adj_4599), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(155[5] 159[10])
    defparam mux_27_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4564));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4565));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4566));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4567));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38839_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n46741));
    defparam i38839_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13142_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n41862), .I3(GND_net), .O(n18426));   // verilog/coms.v(126[12] 289[6])
    defparam i13142_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13143_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n41862), .I3(GND_net), .O(n18427));   // verilog/coms.v(126[12] 289[6])
    defparam i13143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13144_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n41862), .I3(GND_net), .O(n18428));   // verilog/coms.v(126[12] 289[6])
    defparam i13144_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13145_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n41862), .I3(GND_net), .O(n18429));   // verilog/coms.v(126[12] 289[6])
    defparam i13145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13146_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n41862), .I3(GND_net), .O(n18430));   // verilog/coms.v(126[12] 289[6])
    defparam i13146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13147_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n41862), .I3(GND_net), .O(n18431));   // verilog/coms.v(126[12] 289[6])
    defparam i13147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13148_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n41862), .I3(GND_net), .O(n18432));   // verilog/coms.v(126[12] 289[6])
    defparam i13148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13149_3_lut (.I0(\data_in_frame[20] [7]), .I1(rx_data[7]), 
            .I2(n41862), .I3(GND_net), .O(n18433));   // verilog/coms.v(126[12] 289[6])
    defparam i13149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12578_3_lut (.I0(deadband[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n17862));   // verilog/coms.v(126[12] 289[6])
    defparam i12578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13105_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n41860), .I3(GND_net), .O(n18389));   // verilog/coms.v(126[12] 289[6])
    defparam i13105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4568));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4807));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38795_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n46697));
    defparam i38795_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4809));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3032[2]), 
            .I3(r_SM_Main[0]), .O(n17632));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n17632), 
            .I3(rx_data_ready), .O(n41150));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 div_15_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4811));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4821));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4825));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4721));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13106_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n41860), .I3(GND_net), .O(n18390));   // verilog/coms.v(126[12] 289[6])
    defparam i13106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4569));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4824));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13107_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n41860), .I3(GND_net), .O(n18391));   // verilog/coms.v(126[12] 289[6])
    defparam i13107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i38801_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n46703));
    defparam i38801_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13108_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n41860), .I3(GND_net), .O(n18392));   // verilog/coms.v(126[12] 289[6])
    defparam i13108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13109_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n41860), .I3(GND_net), .O(n18393));   // verilog/coms.v(126[12] 289[6])
    defparam i13109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4822));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12859_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n14276), .I3(GND_net), .O(n18143));   // verilog/coms.v(126[12] 289[6])
    defparam i12859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12860_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n14276), .I3(GND_net), .O(n18144));   // verilog/coms.v(126[12] 289[6])
    defparam i12860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12861_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n14276), .I3(GND_net), .O(n18145));   // verilog/coms.v(126[12] 289[6])
    defparam i12861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n526));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n89), .I1(n88), .I2(n87), .I3(n16648), 
            .O(n16639));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1650 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[14] [4]), .I3(\data_in_frame[14] [5]), .O(n37_adj_4974));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 div_15_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4817));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4818));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4819));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12862_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n14276), .I3(GND_net), .O(n18146));   // verilog/coms.v(126[12] 289[6])
    defparam i12862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12863_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n14276), .I3(GND_net), .O(n18147));   // verilog/coms.v(126[12] 289[6])
    defparam i12863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12864_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n14276), .I3(GND_net), .O(n18148));   // verilog/coms.v(126[12] 289[6])
    defparam i12864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4570));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12865_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n14276), .I3(GND_net), .O(n18149));   // verilog/coms.v(126[12] 289[6])
    defparam i12865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12866_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n14276), .I3(GND_net), .O(n18150));   // verilog/coms.v(126[12] 289[6])
    defparam i12866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12867_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n14276), .I3(GND_net), .O(n18151));   // verilog/coms.v(126[12] 289[6])
    defparam i12867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12868_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n14276), .I3(GND_net), .O(n18152));   // verilog/coms.v(126[12] 289[6])
    defparam i12868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4814));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12869_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n14276), .I3(GND_net), .O(n18153));   // verilog/coms.v(126[12] 289[6])
    defparam i12869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12870_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n14276), .I3(GND_net), .O(n18154));   // verilog/coms.v(126[12] 289[6])
    defparam i12870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4816));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12871_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n14276), .I3(GND_net), .O(n18155));   // verilog/coms.v(126[12] 289[6])
    defparam i12871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12872_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n14276), .I3(GND_net), .O(n18156));   // verilog/coms.v(126[12] 289[6])
    defparam i12872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12873_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n14276), .I3(GND_net), .O(n18157));   // verilog/coms.v(126[12] 289[6])
    defparam i12873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12874_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n14276), .I3(GND_net), .O(n18158));   // verilog/coms.v(126[12] 289[6])
    defparam i12874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4571));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12875_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n14276), .I3(GND_net), .O(n18159));   // verilog/coms.v(126[12] 289[6])
    defparam i12875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12876_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n14276), .I3(GND_net), .O(n18160));   // verilog/coms.v(126[12] 289[6])
    defparam i12876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12877_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n14276), .I3(GND_net), .O(n18161));   // verilog/coms.v(126[12] 289[6])
    defparam i12877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12878_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n14276), .I3(GND_net), .O(n18162));   // verilog/coms.v(126[12] 289[6])
    defparam i12878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4572));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4573));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4574));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i719_3_lut (.I0(n1043), .I1(n6446), .I2(n1067), .I3(GND_net), 
            .O(n1169));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i802_3_lut (.I0(n1169), .I1(n6455), .I2(n1193), .I3(GND_net), 
            .O(n1292));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i883_3_lut (.I0(n1292), .I1(n6465), .I2(n1316), .I3(GND_net), 
            .O(n1412));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i962_3_lut (.I0(n1412), .I1(n6476), .I2(n1436), .I3(GND_net), 
            .O(n1529));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_i1039_3_lut (.I0(n1529), .I1(n6488), .I2(n1553), .I3(GND_net), 
            .O(n1643));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12879_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n14276), .I3(GND_net), .O(n18163));   // verilog/coms.v(126[12] 289[6])
    defparam i12879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12880_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n14276), .I3(GND_net), .O(n18164));   // verilog/coms.v(126[12] 289[6])
    defparam i12880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12881_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n14276), .I3(GND_net), .O(n18165));   // verilog/coms.v(126[12] 289[6])
    defparam i12881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12882_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n14276), .I3(GND_net), .O(n18166));   // verilog/coms.v(126[12] 289[6])
    defparam i12882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12883_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n14276), .I3(GND_net), .O(n18167));   // verilog/coms.v(126[12] 289[6])
    defparam i12883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12884_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n14276), .I3(GND_net), .O(n18168));   // verilog/coms.v(126[12] 289[6])
    defparam i12884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12885_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n14276), .I3(GND_net), .O(n18169));   // verilog/coms.v(126[12] 289[6])
    defparam i12885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12886_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n14276), .I3(GND_net), .O(n18170));   // verilog/coms.v(126[12] 289[6])
    defparam i12886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12887_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n14276), .I3(GND_net), .O(n18171));   // verilog/coms.v(126[12] 289[6])
    defparam i12887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12888_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n14276), .I3(GND_net), .O(n18172));   // verilog/coms.v(126[12] 289[6])
    defparam i12888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12889_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n14276), .I3(GND_net), .O(n18173));   // verilog/coms.v(126[12] 289[6])
    defparam i12889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12890_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n14276), .I3(GND_net), .O(n18174));   // verilog/coms.v(126[12] 289[6])
    defparam i12890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12891_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n14276), .I3(GND_net), .O(n18175));   // verilog/coms.v(126[12] 289[6])
    defparam i12891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12892_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n14276), .I3(GND_net), .O(n18176));   // verilog/coms.v(126[12] 289[6])
    defparam i12892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12893_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n14276), .I3(GND_net), .O(n18177));   // verilog/coms.v(126[12] 289[6])
    defparam i12893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12894_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n14276), .I3(GND_net), .O(n18178));   // verilog/coms.v(126[12] 289[6])
    defparam i12894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12895_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n14276), .I3(GND_net), .O(n18179));   // verilog/coms.v(126[12] 289[6])
    defparam i12895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12896_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n14276), .I3(GND_net), .O(n18180));   // verilog/coms.v(126[12] 289[6])
    defparam i12896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12897_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n14276), .I3(GND_net), .O(n18181));   // verilog/coms.v(126[12] 289[6])
    defparam i12897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12898_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n14276), .I3(GND_net), .O(n18182));   // verilog/coms.v(126[12] 289[6])
    defparam i12898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12899_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n14276), .I3(GND_net), .O(n18183));   // verilog/coms.v(126[12] 289[6])
    defparam i12899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12900_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n14276), .I3(GND_net), .O(n18184));   // verilog/coms.v(126[12] 289[6])
    defparam i12900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12901_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n14276), .I3(GND_net), .O(n18185));   // verilog/coms.v(126[12] 289[6])
    defparam i12901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12902_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n14276), .I3(GND_net), .O(n18186));   // verilog/coms.v(126[12] 289[6])
    defparam i12902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12903_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n14276), .I3(GND_net), .O(n18187));   // verilog/coms.v(126[12] 289[6])
    defparam i12903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12904_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n14276), .I3(GND_net), .O(n18188));   // verilog/coms.v(126[12] 289[6])
    defparam i12904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12905_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n14276), .I3(GND_net), .O(n18189));   // verilog/coms.v(126[12] 289[6])
    defparam i12905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12906_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n14276), .I3(GND_net), .O(n18190));   // verilog/coms.v(126[12] 289[6])
    defparam i12906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12907_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n14276), .I3(GND_net), .O(n18191));   // verilog/coms.v(126[12] 289[6])
    defparam i12907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12908_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n14276), .I3(GND_net), .O(n18192));   // verilog/coms.v(126[12] 289[6])
    defparam i12908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12909_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n14276), .I3(GND_net), .O(n18193));   // verilog/coms.v(126[12] 289[6])
    defparam i12909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12910_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n14276), .I3(GND_net), .O(n18194));   // verilog/coms.v(126[12] 289[6])
    defparam i12910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12911_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n14276), .I3(GND_net), .O(n18195));   // verilog/coms.v(126[12] 289[6])
    defparam i12911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12912_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n14276), .I3(GND_net), .O(n18196));   // verilog/coms.v(126[12] 289[6])
    defparam i12912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12913_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n14276), .I3(GND_net), .O(n18197));   // verilog/coms.v(126[12] 289[6])
    defparam i12913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12914_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n14276), .I3(GND_net), .O(n18198));   // verilog/coms.v(126[12] 289[6])
    defparam i12914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12915_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n14276), .I3(GND_net), .O(n18199));   // verilog/coms.v(126[12] 289[6])
    defparam i12915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4827));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i39117_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n47019));
    defparam i39117_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12916_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n14276), .I3(GND_net), .O(n18200));   // verilog/coms.v(126[12] 289[6])
    defparam i12916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4575));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4808));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i40605_4_lut (.I0(n44_adj_4747), .I1(n48506), .I2(n45_adj_4748), 
            .I3(n48449), .O(n48508));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40605_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_15_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4810));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12917_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n14276), .I3(GND_net), .O(n18201));   // verilog/coms.v(126[12] 289[6])
    defparam i12917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12918_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n14276), .I3(GND_net), .O(n18202));   // verilog/coms.v(126[12] 289[6])
    defparam i12918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1651 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(n42342), .I3(GND_net), .O(n42216));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_adj_1651.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(n42140), .I3(GND_net), .O(n4_adj_4604));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 i39090_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n46992));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39090_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4696));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4577), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39119_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n47021));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39119_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4689));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4576));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n48508), .I1(n16648), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hceef;
    SB_LUT4 i12919_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n14276), .I3(GND_net), .O(n18203));   // verilog/coms.v(126[12] 289[6])
    defparam i12919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4687));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12920_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n14276), .I3(GND_net), .O(n18204));   // verilog/coms.v(126[12] 289[6])
    defparam i12920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41879_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n49780));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41879_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i39139_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n47041));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39139_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12921_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n14276), .I3(GND_net), .O(n18205));   // verilog/coms.v(126[12] 289[6])
    defparam i12921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12922_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n14276), .I3(GND_net), .O(n18206));   // verilog/coms.v(126[12] 289[6])
    defparam i12922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12923_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n14276), .I3(GND_net), .O(n18207));   // verilog/coms.v(126[12] 289[6])
    defparam i12923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12924_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n14276), .I3(GND_net), .O(n18208));   // verilog/coms.v(126[12] 289[6])
    defparam i12924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12925_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n14276), .I3(GND_net), .O(n18209));   // verilog/coms.v(126[12] 289[6])
    defparam i12925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12926_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n14276), .I3(GND_net), .O(n18210));   // verilog/coms.v(126[12] 289[6])
    defparam i12926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12927_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n14276), .I3(GND_net), .O(n18211));   // verilog/coms.v(126[12] 289[6])
    defparam i12927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12928_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n14276), .I3(GND_net), .O(n18212));   // verilog/coms.v(126[12] 289[6])
    defparam i12928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4685));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12929_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n14276), .I3(GND_net), .O(n18213));   // verilog/coms.v(126[12] 289[6])
    defparam i12929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12930_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n14276), .I3(GND_net), .O(n18214));   // verilog/coms.v(126[12] 289[6])
    defparam i12930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39153_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n47055));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39153_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4829));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4831));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i39069_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n46971));
    defparam i39069_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4833));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n16614), 
            .O(n249));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_15_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4683));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [3]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n13_adj_4980));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1654 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[14] [5]), .I3(GND_net), .O(n42066));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_adj_1654.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(n37696), .I3(\data_in_frame[9] [6]), .O(n41916));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(n88), .I1(n87), .I2(n16648), 
            .I3(GND_net), .O(n16642));
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'hf7f7;
    SB_LUT4 i39159_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n47061));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i39159_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_i1655_3_lut_3_lut (.I0(n2471), .I1(n6654), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1642_3_lut_3_lut (.I0(n2471), .I1(n6641), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1656 (.I0(n90), .I1(n89), .I2(n16642), 
            .I3(GND_net), .O(n16636));
    defparam i1_2_lut_3_lut_adj_1656.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4849));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1657 (.I0(n91), .I1(n90), .I2(n16639), 
            .I3(GND_net), .O(n16633));
    defparam i1_2_lut_3_lut_adj_1657.LUT_INIT = 16'hf7f7;
    SB_LUT4 i39047_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n46949));
    defparam i39047_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_i1643_3_lut_3_lut (.I0(n2471), .I1(n6642), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1658 (.I0(n92), .I1(n91), .I2(n16636), 
            .I3(GND_net), .O(n16630));
    defparam i1_2_lut_3_lut_adj_1658.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4851));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1659 (.I0(n93), .I1(n92), .I2(n16633), 
            .I3(GND_net), .O(n16627));
    defparam i1_2_lut_3_lut_adj_1659.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1660 (.I0(n94), .I1(n93), .I2(n16630), 
            .I3(GND_net), .O(n16624));
    defparam i1_2_lut_3_lut_adj_1660.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_i1644_3_lut_3_lut (.I0(n2471), .I1(n6643), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1647_3_lut_3_lut (.I0(n2471), .I1(n6646), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1645_3_lut_3_lut (.I0(n2471), .I1(n6644), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4853));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38979_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n46881));
    defparam i38979_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4855));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1648_3_lut_3_lut (.I0(n2471), .I1(n6647), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4871));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1661_3_lut_3_lut (.I0(n2471), .I1(n6660), .I2(n528), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1650_3_lut_3_lut (.I0(n2471), .I1(n6649), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1651_3_lut_3_lut (.I0(n2471), .I1(n6650), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38947_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n46849));
    defparam i38947_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i12931_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n14276), .I3(GND_net), .O(n18215));   // verilog/coms.v(126[12] 289[6])
    defparam i12931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1646_3_lut_3_lut (.I0(n2471), .I1(n6645), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1657_3_lut_3_lut (.I0(n2471), .I1(n6656), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12932_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n14276), .I3(GND_net), .O(n18216));   // verilog/coms.v(126[12] 289[6])
    defparam i12932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12933_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n14276), .I3(GND_net), .O(n18217));   // verilog/coms.v(126[12] 289[6])
    defparam i12933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12934_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n14276), .I3(GND_net), .O(n18218));   // verilog/coms.v(126[12] 289[6])
    defparam i12934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12935_3_lut (.I0(\data_out_frame[15] [0]), .I1(pwm[16]), .I2(n14276), 
            .I3(GND_net), .O(n18219));   // verilog/coms.v(126[12] 289[6])
    defparam i12935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12936_3_lut (.I0(\data_out_frame[15] [1]), .I1(pwm[17]), .I2(n14276), 
            .I3(GND_net), .O(n18220));   // verilog/coms.v(126[12] 289[6])
    defparam i12936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12937_3_lut (.I0(\data_out_frame[15] [2]), .I1(pwm[18]), .I2(n14276), 
            .I3(GND_net), .O(n18221));   // verilog/coms.v(126[12] 289[6])
    defparam i12937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12938_3_lut (.I0(\data_out_frame[15] [3]), .I1(pwm[19]), .I2(n14276), 
            .I3(GND_net), .O(n18222));   // verilog/coms.v(126[12] 289[6])
    defparam i12938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12939_3_lut (.I0(\data_out_frame[15] [4]), .I1(pwm[20]), .I2(n14276), 
            .I3(GND_net), .O(n18223));   // verilog/coms.v(126[12] 289[6])
    defparam i12939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12940_3_lut (.I0(\data_out_frame[15] [5]), .I1(pwm[21]), .I2(n14276), 
            .I3(GND_net), .O(n18224));   // verilog/coms.v(126[12] 289[6])
    defparam i12940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12941_3_lut (.I0(\data_out_frame[15] [6]), .I1(pwm[22]), .I2(n14276), 
            .I3(GND_net), .O(n18225));   // verilog/coms.v(126[12] 289[6])
    defparam i12941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12942_3_lut (.I0(\data_out_frame[15] [7]), .I1(pwm[23]), .I2(n14276), 
            .I3(GND_net), .O(n18226));   // verilog/coms.v(126[12] 289[6])
    defparam i12942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12943_3_lut (.I0(\data_out_frame[16] [0]), .I1(pwm[8]), .I2(n14276), 
            .I3(GND_net), .O(n18227));   // verilog/coms.v(126[12] 289[6])
    defparam i12943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4873));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1659_3_lut_3_lut (.I0(n2471), .I1(n6658), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1658_3_lut_3_lut (.I0(n2471), .I1(n6657), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4875));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38906_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n46808));
    defparam i38906_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4877));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1654_3_lut_3_lut (.I0(n2471), .I1(n6653), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1653_3_lut_3_lut (.I0(n2471), .I1(n6652), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4893));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1652_3_lut_3_lut (.I0(n2471), .I1(n6651), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4897));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1656_3_lut_3_lut (.I0(n2471), .I1(n6655), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38817_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n46719));
    defparam i38817_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_i1649_3_lut_3_lut (.I0(n2471), .I1(n6648), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1660_3_lut_3_lut (.I0(n2471), .I1(n6659), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1707_3_lut_3_lut (.I0(n2558), .I1(n6671), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1699_3_lut_3_lut (.I0(n2558), .I1(n6663), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1700_3_lut_3_lut (.I0(n2558), .I1(n6664), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1701_3_lut_3_lut (.I0(n2558), .I1(n6665), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4899));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4895));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1702_3_lut_3_lut (.I0(n2558), .I1(n6666), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1705_3_lut_3_lut (.I0(n2558), .I1(n6669), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1703_3_lut_3_lut (.I0(n2558), .I1(n6667), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1706_3_lut_3_lut (.I0(n2558), .I1(n6670), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1719_3_lut_3_lut (.I0(n2558), .I1(n6683), .I2(n529), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1704_3_lut_3_lut (.I0(n2558), .I1(n6668), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1708_3_lut_3_lut (.I0(n2558), .I1(n6672), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1709_3_lut_3_lut (.I0(n2558), .I1(n6673), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4812));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i38857_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n46759));
    defparam i38857_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4813));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4733));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4915));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4919));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i39558_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n47461));
    defparam i39558_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4806));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1710_3_lut_3_lut (.I0(n2558), .I1(n6674), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4921));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38803_4_lut (.I0(n23_adj_4812), .I1(n21_adj_4810), .I2(n19_adj_4808), 
            .I3(n17_adj_4806), .O(n46705));
    defparam i38803_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_i1711_3_lut_3_lut (.I0(n2558), .I1(n6675), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38799_4_lut (.I0(n29_adj_4816), .I1(n27_adj_4814), .I2(n25_adj_4813), 
            .I3(n46705), .O(n46701));
    defparam i38799_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_15_i1715_3_lut_3_lut (.I0(n2558), .I1(n6679), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i40480_4_lut (.I0(n35_adj_4819), .I1(n33_adj_4818), .I2(n31_adj_4817), 
            .I3(n46701), .O(n48383));
    defparam i40480_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_15_i1718_3_lut_3_lut (.I0(n2558), .I1(n6682), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1717_3_lut_3_lut (.I0(n2558), .I1(n6681), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1482_i16_4_lut (.I0(n526), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4805));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i40729_3_lut (.I0(n16_adj_4805), .I1(n87), .I2(n39_adj_4822), 
            .I3(GND_net), .O(n48632));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40729_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i38937_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n46839));
    defparam i38937_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4917));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i39589_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n47492));
    defparam i39589_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i40730_3_lut (.I0(n48632), .I1(n86), .I2(n41_adj_4824), .I3(GND_net), 
            .O(n48633));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40730_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1404_3_lut_3_lut (.I0(n2093), .I1(n6573), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1716_3_lut_3_lut (.I0(n2558), .I1(n6680), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i39596_4_lut (.I0(n41_adj_4824), .I1(n39_adj_4822), .I2(n27_adj_4814), 
            .I3(n46703), .O(n47499));
    defparam i39596_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40627_3_lut (.I0(n22_adj_4811), .I1(n93), .I2(n27_adj_4814), 
            .I3(GND_net), .O(n48530));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40627_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4735));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1712_3_lut_3_lut (.I0(n2558), .I1(n6676), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38943_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n46845));
    defparam i38943_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4737));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i40626_3_lut (.I0(n48633), .I1(n85), .I2(n43_adj_4825), .I3(GND_net), 
            .O(n40_adj_4823));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40626_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1407_3_lut_3_lut (.I0(n2093), .I1(n6576), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1714_3_lut_3_lut (.I0(n2558), .I1(n6678), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38963_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n46865));
    defparam i38963_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4723));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1406_3_lut_3_lut (.I0(n2093), .I1(n6575), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1482_i28_3_lut (.I0(n20_adj_4809), .I1(n91), 
            .I2(n31_adj_4817), .I3(GND_net), .O(n28_adj_4815));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41039_4_lut (.I0(n28_adj_4815), .I1(n18_adj_4807), .I2(n31_adj_4817), 
            .I3(n46697), .O(n48942));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41039_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41040_3_lut (.I0(n48942), .I1(n90), .I2(n33_adj_4818), .I3(GND_net), 
            .O(n48943));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i41040_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_15_i1713_3_lut_3_lut (.I0(n2558), .I1(n6677), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1397_3_lut_3_lut (.I0(n2093), .I1(n6566), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36354_2_lut_4_lut (.I0(r_Clock_Count_adj_5025[7]), .I1(r_Clock_Count_adj_5025[6]), 
            .I2(r_Clock_Count_adj_5025[8]), .I3(n88_adj_4963), .O(n44245));
    defparam i36354_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i40925_3_lut (.I0(n48943), .I1(n89), .I2(n35_adj_4819), .I3(GND_net), 
            .O(n48828));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40925_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i39600_4_lut (.I0(n41_adj_4824), .I1(n39_adj_4822), .I2(n37_adj_4821), 
            .I3(n48383), .O(n47503));
    defparam i39600_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40787_4_lut (.I0(n40_adj_4823), .I1(n48530), .I2(n43_adj_4825), 
            .I3(n47499), .O(n48690));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40787_4_lut.LUT_INIT = 16'haaac;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n18531(n18531), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n18530(n18530), .n18529(n18529), .n18528(n18528), 
            .n18527(n18527), .n18526(n18526), .n18525(n18525), .n18524(n18524), 
            .n18523(n18523), .n18522(n18522), .n18521(n18521), .n18520(n18520), 
            .n18519(n18519), .n18518(n18518), .n18517(n18517), .n18516(n18516), 
            .n18515(n18515), .n18514(n18514), .n18513(n18513), .n18512(n18512), 
            .n18511(n18511), .n18510(n18510), .n18497(n18497), .data_o({quadA_debounced, 
            quadB_debounced}), .n2642({n2643, n2644, n2645, n2646, 
            n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
            n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
            n2663, n2664, n2665, n2666}), .GND_net(GND_net), .n17969(n17969), 
            .count_enable(count_enable), .n18616(n18616), .reg_B({reg_B}), 
            .PIN_23_c_1(PIN_23_c_1), .PIN_24_c_0(PIN_24_c_0), .n17971(n17971), 
            .n44088(n44088)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(184[15] 189[4])
    SB_LUT4 i28742_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n511), .I3(n558), 
            .O(n4_adj_4561));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28742_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_15_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4710));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38987_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n46889));
    defparam i38987_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4712));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4700));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i39045_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n46947));
    defparam i39045_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4701));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_4_lut_adj_1661 (.I0(n86), .I1(n85), .I2(n84), .I3(n16657), 
            .O(n16648));
    defparam i1_2_lut_4_lut_adj_1661.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1662 (.I0(n85), .I1(n84), .I2(n16657), 
            .I3(GND_net), .O(n16651));
    defparam i1_2_lut_3_lut_adj_1662.LUT_INIT = 16'hf7f7;
    SB_LUT4 i28807_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n512), .I3(n558), 
            .O(n4_adj_4965));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28807_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i28839_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n513), .I3(n558), 
            .O(n4));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i28839_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_3_lut_adj_1663 (.I0(n98), .I1(n97), .I2(n16617), 
            .I3(GND_net), .O(n16614));
    defparam i1_2_lut_3_lut_adj_1663.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1664 (.I0(n96), .I1(n95), .I2(n94), .I3(n16627), 
            .O(n16617));
    defparam i1_2_lut_4_lut_adj_1664.LUT_INIT = 16'hff7f;
    SB_LUT4 div_15_i1396_3_lut_3_lut (.I0(n2093), .I1(n6565), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1665 (.I0(n95), .I1(n94), .I2(n16627), 
            .I3(GND_net), .O(n16621));
    defparam i1_2_lut_3_lut_adj_1665.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4751));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38898_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n46800));
    defparam i38898_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4753));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38902_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n46804));
    defparam i38902_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4755));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i40864_3_lut (.I0(n48828), .I1(n88), .I2(n37_adj_4821), .I3(GND_net), 
            .O(n36_adj_4820));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40864_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i40974_4_lut (.I0(n36_adj_4820), .I1(n48690), .I2(n43_adj_4825), 
            .I3(n47503), .O(n48877));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40974_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i40975_3_lut (.I0(n48877), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n48878));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam i40975_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1666 (.I0(n48878), .I1(n16660), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'hceef;
    SB_LUT4 div_15_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4769));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i38870_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n46772));
    defparam i38870_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4800));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12944_3_lut (.I0(\data_out_frame[16] [1]), .I1(pwm[9]), .I2(n14276), 
            .I3(GND_net), .O(n18228));   // verilog/coms.v(126[12] 289[6])
    defparam i12944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12945_3_lut (.I0(\data_out_frame[16] [2]), .I1(pwm[10]), .I2(n14276), 
            .I3(GND_net), .O(n18229));   // verilog/coms.v(126[12] 289[6])
    defparam i12945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12946_3_lut (.I0(\data_out_frame[16] [3]), .I1(pwm[11]), .I2(n14276), 
            .I3(GND_net), .O(n18230));   // verilog/coms.v(126[12] 289[6])
    defparam i12946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4771));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4598));   // verilog/TinyFPGA_B.v(180[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1395_3_lut_3_lut (.I0(n2093), .I1(n6564), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1398_3_lut_3_lut (.I0(n2093), .I1(n6567), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38877_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n46779));
    defparam i38877_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4773));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12947_3_lut (.I0(\data_out_frame[16] [4]), .I1(pwm[12]), .I2(n14276), 
            .I3(GND_net), .O(n18231));   // verilog/coms.v(126[12] 289[6])
    defparam i12947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12948_3_lut (.I0(\data_out_frame[16] [5]), .I1(pwm[13]), .I2(n14276), 
            .I3(GND_net), .O(n18232));   // verilog/coms.v(126[12] 289[6])
    defparam i12948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12949_3_lut (.I0(\data_out_frame[16] [6]), .I1(pwm[14]), .I2(n14276), 
            .I3(GND_net), .O(n18233));   // verilog/coms.v(126[12] 289[6])
    defparam i12949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12950_3_lut (.I0(\data_out_frame[16] [7]), .I1(pwm[15]), .I2(n14276), 
            .I3(GND_net), .O(n18234));   // verilog/coms.v(126[12] 289[6])
    defparam i12950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12951_3_lut (.I0(\data_out_frame[17] [0]), .I1(pwm[0]), .I2(n14276), 
            .I3(GND_net), .O(n18235));   // verilog/coms.v(126[12] 289[6])
    defparam i12951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12952_3_lut (.I0(\data_out_frame[17] [1]), .I1(pwm[1]), .I2(n14276), 
            .I3(GND_net), .O(n18236));   // verilog/coms.v(126[12] 289[6])
    defparam i12952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12953_3_lut (.I0(\data_out_frame[17] [2]), .I1(pwm[2]), .I2(n14276), 
            .I3(GND_net), .O(n18237));   // verilog/coms.v(126[12] 289[6])
    defparam i12953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12954_3_lut (.I0(\data_out_frame[17] [3]), .I1(pwm[3]), .I2(n14276), 
            .I3(GND_net), .O(n18238));   // verilog/coms.v(126[12] 289[6])
    defparam i12954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4804));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12955_3_lut (.I0(\data_out_frame[17] [4]), .I1(pwm[4]), .I2(n14276), 
            .I3(GND_net), .O(n18239));   // verilog/coms.v(126[12] 289[6])
    defparam i12955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4803));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4801));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1667 (.I0(n83), .I1(n82), .I2(n81), .I3(n16666), 
            .O(n16657));
    defparam i1_2_lut_4_lut_adj_1667.LUT_INIT = 16'hff7f;
    SB_LUT4 div_15_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4658));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4657));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1668 (.I0(n82), .I1(n81), .I2(n16666), 
            .I3(GND_net), .O(n16660));
    defparam i1_2_lut_3_lut_adj_1668.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4656));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12956_3_lut (.I0(\data_out_frame[17] [5]), .I1(pwm[5]), .I2(n14276), 
            .I3(GND_net), .O(n18240));   // verilog/coms.v(126[12] 289[6])
    defparam i12956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4655));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4654));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4787));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4653));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4789));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4652));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12957_3_lut (.I0(\data_out_frame[17] [6]), .I1(pwm[6]), .I2(n14276), 
            .I3(GND_net), .O(n18241));   // verilog/coms.v(126[12] 289[6])
    defparam i12957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4651));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12958_3_lut (.I0(\data_out_frame[17] [7]), .I1(pwm[7]), .I2(n14276), 
            .I3(GND_net), .O(n18242));   // verilog/coms.v(126[12] 289[6])
    defparam i12958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4650));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1669 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n16666));
    defparam i1_2_lut_4_lut_adj_1669.LUT_INIT = 16'hff7f;
    SB_LUT4 div_15_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n525));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4649));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4648));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4647));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12959_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n14276), .I3(GND_net), .O(n18243));   // verilog/coms.v(126[12] 289[6])
    defparam i12959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1670 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n16669));
    defparam i1_2_lut_3_lut_adj_1670.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_15_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4646));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12960_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n14276), .I3(GND_net), .O(n18244));   // verilog/coms.v(126[12] 289[6])
    defparam i12960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12961_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n14276), .I3(GND_net), .O(n18245));   // verilog/coms.v(126[12] 289[6])
    defparam i12961_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    SB_LUT4 i12962_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n14276), .I3(GND_net), .O(n18246));   // verilog/coms.v(126[12] 289[6])
    defparam i12962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1394_3_lut_3_lut (.I0(n2093), .I1(n6563), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    coms setpoint_23__I_0 (.n23171(n23171), .PWMLimit({PWMLimit}), .clk32MHz(clk32MHz), 
         .n18460(n18460), .n18459(n18459), .n18458(n18458), .n18457(n18457), 
         .GND_net(GND_net), .n18456(n18456), .n18455(n18455), .n18454(n18454), 
         .n18453(n18453), .n18452(n18452), .n18451(n18451), .n18450(n18450), 
         .n18449(n18449), .n18448(n18448), .control_mode({control_mode}), 
         .rx_data({rx_data}), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n18447(n18447), .\data_in_frame[19] ({\data_in_frame[19] }), .\data_in_frame[14] ({Open_0, 
         \data_in_frame[14] [6:4], Open_1, Open_2, \data_in_frame[14] [1:0]}), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n18329(n18329), .\data_in_frame[7] ({\data_in_frame[7] }), .n18328(n18328), 
         .n18327(n18327), .n18326(n18326), .n18325(n18325), .n18324(n18324), 
         .n18323(n18323), .n18369(n18369), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n18667(n18667), .setpoint({setpoint}), .n18666(n18666), .n18665(n18665), 
         .n18664(n18664), .n18663(n18663), .n18662(n18662), .n18661(n18661), 
         .n18660(n18660), .n18659(n18659), .n18658(n18658), .n18657(n18657), 
         .n18656(n18656), .n18655(n18655), .n18654(n18654), .n18653(n18653), 
         .n18652(n18652), .n18651(n18651), .n18650(n18650), .n18649(n18649), 
         .n18648(n18648), .n18647(n18647), .n18646(n18646), .n18645(n18645), 
         .n18368(n18368), .n18367(n18367), .n18366(n18366), .n18365(n18365), 
         .n18593(n18593), .VCC_net(VCC_net), .byte_transmit_counter({Open_3, 
         Open_4, Open_5, Open_6, Open_7, Open_8, Open_9, byte_transmit_counter[0]}), 
         .n18364(n18364), .n18363(n18363), .n18362(n18362), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n18550(n18550), .n18547(n18547), .n18544(n18544), .n18541(n18541), 
         .n18538(n18538), .n18535(n18535), .n18509(n18509), .n50009(n50009), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n18471(n18471), .n18470(n18470), 
         .n18469(n18469), .n18468(n18468), .n18467(n18467), .n18466(n18466), 
         .n23694(n23694), .n18464(n18464), .n18463(n18463), .n18462(n18462), 
         .n18322(n18322), .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n18305(n18305), .\data_in_frame[4] ({\data_in_frame[4] }), .n18304(n18304), 
         .n18303(n18303), .n18302(n18302), .n18301(n18301), .n18300(n18300), 
         .n18299(n18299), .n18298(n18298), .rx_data_ready(rx_data_ready), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .n18446(n18446), .n18445(n18445), 
         .n18444(n18444), .n18443(n18443), .n18442(n18442), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .Kp_23__N_679(Kp_23__N_679), 
         .n17503(n17503), .n37696(n37696), .n43448(n43448), .n18266(n18266), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n18265(n18265), 
         .n18264(n18264), .n18263(n18263), .n18262(n18262), .n18261(n18261), 
         .n18260(n18260), .n18259(n18259), .n18258(n18258), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n18257(n18257), .n18256(n18256), .n18255(n18255), .n18254(n18254), 
         .n18253(n18253), .n18252(n18252), .n18251(n18251), .n18250(n18250), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .n18249(n18249), 
         .n18248(n18248), .n18247(n18247), .n18246(n18246), .n18245(n18245), 
         .n18244(n18244), .n18243(n18243), .n18242(n18242), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n18241(n18241), .n18240(n18240), .n18239(n18239), .n18238(n18238), 
         .n18237(n18237), .n18236(n18236), .n18235(n18235), .n18234(n18234), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .n18233(n18233), 
         .n18232(n18232), .n18231(n18231), .n41851(n41851), .n18230(n18230), 
         .n2857(n2857), .n41860(n41860), .n18229(n18229), .n18228(n18228), 
         .n18227(n18227), .n18226(n18226), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n18225(n18225), .n18224(n18224), .n18223(n18223), .n18222(n18222), 
         .n18221(n18221), .n18220(n18220), .n18219(n18219), .n18218(n18218), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n18217(n18217), 
         .n18216(n18216), .n18215(n18215), .n18214(n18214), .n18213(n18213), 
         .n18212(n18212), .n18211(n18211), .n18210(n18210), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n18209(n18209), .n18208(n18208), .n18207(n18207), .n18206(n18206), 
         .n18205(n18205), .n18204(n18204), .n18203(n18203), .n16563(n16563), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .n18202(n18202), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n18201(n18201), .n41862(n41862), .n18507(n18507), .n4497(n4497), 
         .n18200(n18200), .n18199(n18199), .n18198(n18198), .n18197(n18197), 
         .n18196(n18196), .n18195(n18195), .n18194(n18194), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n18193(n18193), .n18192(n18192), .n18191(n18191), .n18190(n18190), 
         .n18189(n18189), .n18188(n18188), .n18187(n18187), .n18186(n18186), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .n18185(n18185), 
         .n18184(n18184), .n18183(n18183), .n18533(n18533), .n18182(n18182), 
         .n18181(n18181), .n18180(n18180), .n18179(n18179), .n18178(n18178), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .n18177(n18177), .n18176(n18176), 
         .n18175(n18175), .n18174(n18174), .n18173(n18173), .n18172(n18172), 
         .n18171(n18171), .n18170(n18170), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .n18169(n18169), .n18168(n18168), .n18167(n18167), .n18536(n18536), 
         .n18166(n18166), .n18165(n18165), .n18164(n18164), .n18163(n18163), 
         .n41848(n41848), .n41857(n41857), .n18162(n18162), .n18161(n18161), 
         .n18160(n18160), .n18159(n18159), .n18158(n18158), .n18157(n18157), 
         .n18156(n18156), .n18155(n18155), .n18154(n18154), .n18153(n18153), 
         .n18152(n18152), .n18151(n18151), .n18150(n18150), .n18149(n18149), 
         .n18148(n18148), .n18147(n18147), .n18146(n18146), .n18145(n18145), 
         .n18144(n18144), .n18143(n18143), .n18393(n18393), .n18392(n18392), 
         .n18391(n18391), .n18390(n18390), .n18539(n18539), .n18389(n18389), 
         .n17862(n17862), .deadband({deadband}), .n37561(n37561), .n18433(n18433), 
         .n18432(n18432), .n18431(n18431), .n18430(n18430), .n18429(n18429), 
         .n18428(n18428), .n18427(n18427), .n18426(n18426), .n38230(n38230), 
         .n42079(n42079), .n37512(n37512), .n18542(n18542), .n18545(n18545), 
         .n18548(n18548), .n2244(n2244), .n18142(n18142), .n18141(n18141), 
         .n18388(n18388), .n18387(n18387), .n18386(n18386), .n18140(n18140), 
         .n18139(n18139), .n18135(n18135), .\data_in[3] ({\data_in[3] }), 
         .n18134(n18134), .n18133(n18133), .n18132(n18132), .n18131(n18131), 
         .n18130(n18130), .n18129(n18129), .n18128(n18128), .n18127(n18127), 
         .\data_in[2] ({\data_in[2] }), .n18126(n18126), .n18125(n18125), 
         .n18124(n18124), .n18123(n18123), .n18122(n18122), .n18121(n18121), 
         .n18120(n18120), .n18119(n18119), .\data_in[1] ({\data_in[1] }), 
         .n18118(n18118), .n18117(n18117), .n18116(n18116), .n18115(n18115), 
         .n18114(n18114), .n18113(n18113), .n18112(n18112), .n18111(n18111), 
         .\data_in[0] ({\data_in[0] }), .n18110(n18110), .n18109(n18109), 
         .n18108(n18108), .n18107(n18107), .n18106(n18106), .n18105(n18105), 
         .n18104(n18104), .gearBoxRatio({gearBoxRatio}), .n18103(n18103), 
         .n18102(n18102), .n18101(n18101), .n18100(n18100), .n18099(n18099), 
         .n18098(n18098), .n18097(n18097), .n18096(n18096), .n18095(n18095), 
         .n18094(n18094), .n18093(n18093), .n18092(n18092), .n18091(n18091), 
         .n18090(n18090), .n18089(n18089), .n18088(n18088), .n18087(n18087), 
         .n18086(n18086), .n18085(n18085), .n18084(n18084), .n18083(n18083), 
         .n18082(n18082), .n18081(n18081), .\Kd[7] (Kd[7]), .n18080(n18080), 
         .\Kd[6] (Kd[6]), .n18079(n18079), .\Kd[5] (Kd[5]), .n18078(n18078), 
         .\Kd[4] (Kd[4]), .n18077(n18077), .\Kd[3] (Kd[3]), .n18076(n18076), 
         .\Kd[2] (Kd[2]), .n18075(n18075), .\Kd[1] (Kd[1]), .n18074(n18074), 
         .\Ki[7] (Ki[7]), .n18073(n18073), .\Ki[6] (Ki[6]), .n18072(n18072), 
         .\Ki[5] (Ki[5]), .n18071(n18071), .\Ki[4] (Ki[4]), .n18070(n18070), 
         .\Ki[3] (Ki[3]), .n18069(n18069), .\Ki[2] (Ki[2]), .n18068(n18068), 
         .\Ki[1] (Ki[1]), .n18067(n18067), .\Kp[7] (Kp[7]), .n18066(n18066), 
         .\Kp[6] (Kp[6]), .n18065(n18065), .\Kp[5] (Kp[5]), .n18064(n18064), 
         .\Kp[4] (Kp[4]), .n18063(n18063), .\Kp[3] (Kp[3]), .n18062(n18062), 
         .\Kp[2] (Kp[2]), .n18061(n18061), .\Kp[1] (Kp[1]), .n18060(n18060), 
         .IntegralLimit({IntegralLimit}), .n18059(n18059), .n18058(n18058), 
         .n18057(n18057), .n18056(n18056), .n18055(n18055), .n18054(n18054), 
         .n18053(n18053), .n18052(n18052), .n18051(n18051), .n18050(n18050), 
         .n18049(n18049), .n18048(n18048), .n18047(n18047), .n18046(n18046), 
         .n18045(n18045), .n18044(n18044), .n18043(n18043), .n18042(n18042), 
         .n18041(n18041), .n18040(n18040), .n18039(n18039), .n18038(n18038), 
         .n18013(n18013), .n18012(n18012), .n18011(n18011), .n18010(n18010), 
         .n18009(n18009), .n18008(n18008), .n18007(n18007), .n18006(n18006), 
         .n18005(n18005), .n18004(n18004), .n18003(n18003), .n18002(n18002), 
         .n18001(n18001), .n18000(n18000), .n17999(n17999), .n17998(n17998), 
         .n17997(n17997), .n17996(n17996), .n17995(n17995), .n17994(n17994), 
         .n17993(n17993), .n17992(n17992), .n17991(n17991), .n17983(n17983), 
         .n40968(n40968), .n17966(n17966), .n17965(n17965), .n17963(n17963), 
         .n17962(n17962), .n17961(n17961), .\Kd[0] (Kd[0]), .n17960(n17960), 
         .\Ki[0] (Ki[0]), .n17959(n17959), .\Kp[0] (Kp[0]), .n17958(n17958), 
         .LED_c(LED_c), .n123(n123), .n740(n740), .n19921(n19921), .n16687(n16687), 
         .n16678(n16678), .n2484(n2484), .n16680(n16680), .n5(n5_adj_4628), 
         .n7(n7_adj_4629), .n50704(n50704), .n41916(n41916), .n28(n28_adj_4975), 
         .n42216(n42216), .n37(n37_adj_4974), .n42140(n42140), .n42342(n42342), 
         .n42357(n42357), .n14246(n14246), .n16683(n16683), .n42066(n42066), 
         .n42219(n42219), .n42330(n42330), .n42459(n42459), .n42429(n42429), 
         .n43056(n43056), .n15(n15_adj_4978), .n13(n13_adj_4980), .n14(n14_adj_4979), 
         .n42432(n42432), .n25520(n25520), .n4446(n4446), .n4447(n4447), 
         .n4448(n4448), .n4449(n4449), .n4450(n4450), .n14276(n14276), 
         .n3(n3_adj_4597), .n16675(n16675), .n6(n6), .n4451(n4451), 
         .n4452(n4452), .n17283(n17283), .n4453(n4453), .n4454(n4454), 
         .n4455(n4455), .n4456(n4456), .n4457(n4457), .n4458(n4458), 
         .n4459(n4459), .n4460(n4460), .n4461(n4461), .n42696(n42696), 
         .n4462(n4462), .n4463(n4463), .n4464(n4464), .n42610(n42610), 
         .n4465(n4465), .n4466(n4466), .n4467(n4467), .n4469(n4469), 
         .n4468(n4468), .n5_adj_15(n5_adj_4981), .n4(n4_adj_4604), .n19(n19_adj_4973), 
         .n41336(n41336), .n41446(n41446), .n41444(n41444), .n41442(n41442), 
         .n41074(n41074), .\r_Clock_Count[8] (r_Clock_Count_adj_5025[8]), 
         .n41130(n41130), .\r_Clock_Count[7] (r_Clock_Count_adj_5025[7]), 
         .n41224(n41224), .\r_Clock_Count[6] (r_Clock_Count_adj_5025[6]), 
         .n41348(n41348), .tx_o(tx_o), .tx_enable(tx_enable), .n88(n88_adj_4963), 
         .n118(n118), .\r_SM_Main[2] (r_SM_Main_adj_5024[2]), .n5_adj_16(n5_adj_4982), 
         .n44294(n44294), .n17955(n17955), .n17977(n17977), .n17980(n17980), 
         .n17863(n17863), .n17866(n17866), .n17869(n17869), .n17872(n17872), 
         .n18575(n18575), .n17974(n17974), .n3_adj_17(n3_adj_4971), .n17887(n17887), 
         .r_Bit_Index({r_Bit_Index}), .n17890(n17890), .n18701(n18701), 
         .\r_Clock_Count[0] (r_Clock_Count[0]), .r_SM_Main({r_SM_Main}), 
         .n18587(n18587), .n41150(n41150), .n18583(n18583), .n18567(n18567), 
         .\r_Clock_Count[5] (r_Clock_Count[5]), .n18555(n18555), .\r_Clock_Count[1] (r_Clock_Count[1]), 
         .\r_SM_Main_2__N_3032[2] (r_SM_Main_2__N_3032[2]), .r_Rx_Data(r_Rx_Data), 
         .PIN_13_N_50(PIN_13_N_50), .n27708(n27708), .n17657(n17657), 
         .n17707(n17707), .n17849(n17849), .n4694(n4694), .n221(n221), 
         .n225(n225), .n226(n226), .n17897(n17897), .n17896(n17896), 
         .n17895(n17895), .n17894(n17894), .n17893(n17893), .n17892(n17892), 
         .n17891(n17891), .n16566(n16566), .n4_adj_19(n4_adj_4588), .n25329(n25329), 
         .n4_adj_20(n4_adj_4596), .n4_adj_21(n4_adj_4592), .n16432(n16432)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(86[8] 106[4])
    SB_LUT4 i12963_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n14276), .I3(GND_net), .O(n18247));   // verilog/coms.v(126[12] 289[6])
    defparam i12963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1402_3_lut_3_lut (.I0(n2093), .I1(n6571), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4797));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4798));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4799));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4791));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4793));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4794));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4796));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_15_i1403_3_lut_3_lut (.I0(n2093), .I1(n6572), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4785));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i38841_4_lut (.I0(n25_adj_4791), .I1(n23_adj_4789), .I2(n21_adj_4787), 
            .I3(n19_adj_4785), .O(n46743));
    defparam i38841_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38837_4_lut (.I0(n31_adj_4796), .I1(n29_adj_4794), .I2(n27_adj_4793), 
            .I3(n46743), .O(n46739));
    defparam i38837_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40496_4_lut (.I0(n37_adj_4799), .I1(n35_adj_4798), .I2(n33_adj_4797), 
            .I3(n46739), .O(n48399));
    defparam i40496_4_lut.LUT_INIT = 16'hfffe;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n2592({n2593, n2594, n2595, 
            n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, 
            n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
            n2612, n2613, n2614, n2615, n2616}), .encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .n18615(n18615), .clk32MHz(clk32MHz), .n18614(n18614), 
            .n18613(n18613), .n18612(n18612), .n18611(n18611), .n18610(n18610), 
            .n18609(n18609), .n18608(n18608), .n18607(n18607), .n18606(n18606), 
            .n18605(n18605), .n18604(n18604), .n18603(n18603), .n18602(n18602), 
            .n18601(n18601), .n18600(n18600), .n18599(n18599), .n18598(n18598), 
            .n18597(n18597), .n18596(n18596), .n18595(n18595), .n18594(n18594), 
            .n18532(n18532), .data_o({quadA_debounced_adj_4589, quadB_debounced_adj_4590}), 
            .n17970(n17970), .count_enable(count_enable_adj_4591), .PIN_18_c_1(PIN_18_c_1), 
            .n18618(n18618), .reg_B({reg_B_adj_5037}), .PIN_19_c_0(PIN_19_c_0), 
            .n17973(n17973), .n43352(n43352)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(192[15] 197[4])
    SB_LUT4 div_15_i1405_3_lut_3_lut (.I0(n2093), .I1(n6574), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1408_3_lut_3_lut (.I0(n2093), .I1(n6577), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12964_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n14276), .I3(GND_net), .O(n18248));   // verilog/coms.v(126[12] 289[6])
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12965_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n14276), .I3(GND_net), .O(n18249));   // verilog/coms.v(126[12] 289[6])
    defparam i12965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12966_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n14276), .I3(GND_net), .O(n18250));   // verilog/coms.v(126[12] 289[6])
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4645));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4644));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4643));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12967_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n14276), .I3(GND_net), .O(n18251));   // verilog/coms.v(126[12] 289[6])
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12968_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n14276), .I3(GND_net), .O(n18252));   // verilog/coms.v(126[12] 289[6])
    defparam i12968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4642));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12969_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n14276), .I3(GND_net), .O(n18253));   // verilog/coms.v(126[12] 289[6])
    defparam i12969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12970_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n14276), .I3(GND_net), .O(n18254));   // verilog/coms.v(126[12] 289[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12971_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n14276), .I3(GND_net), .O(n18255));   // verilog/coms.v(126[12] 289[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12972_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n14276), .I3(GND_net), .O(n18256));   // verilog/coms.v(126[12] 289[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12973_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n14276), .I3(GND_net), .O(n18257));   // verilog/coms.v(126[12] 289[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12974_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n14276), .I3(GND_net), .O(n18258));   // verilog/coms.v(126[12] 289[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1401_3_lut_3_lut (.I0(n2093), .I1(n6570), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1399_3_lut_3_lut (.I0(n2093), .I1(n6568), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1400_3_lut_3_lut (.I0(n2093), .I1(n6569), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12975_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n14276), .I3(GND_net), .O(n18259));   // verilog/coms.v(126[12] 289[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12976_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n14276), .I3(GND_net), .O(n18260));   // verilog/coms.v(126[12] 289[6])
    defparam i12976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12977_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n14276), .I3(GND_net), .O(n18261));   // verilog/coms.v(126[12] 289[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12978_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n14276), .I3(GND_net), .O(n18262));   // verilog/coms.v(126[12] 289[6])
    defparam i12978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12979_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n14276), .I3(GND_net), .O(n18263));   // verilog/coms.v(126[12] 289[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12980_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n14276), .I3(GND_net), .O(n18264));   // verilog/coms.v(126[12] 289[6])
    defparam i12980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12981_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n14276), .I3(GND_net), .O(n18265));   // verilog/coms.v(126[12] 289[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1409_3_lut_3_lut (.I0(n2093), .I1(n6578), .I2(n524), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i17902_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[6] [5]), 
            .I2(n3_adj_4597), .I3(GND_net), .O(n23171));
    defparam i17902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_15_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4790));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_i1769_3_lut_3_lut (.I0(n2642), .I1(n6701), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12982_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n14276), .I3(GND_net), .O(n18266));   // verilog/coms.v(126[12] 289[6])
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_i1754_3_lut_3_lut (.I0(n2642), .I1(n6686), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4641));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4640));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4639));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1755_3_lut_3_lut (.I0(n2642), .I1(n6687), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1757_3_lut_3_lut (.I0(n2642), .I1(n6689), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1756_3_lut_3_lut (.I0(n2642), .I1(n6688), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4638));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4637));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1758_3_lut_3_lut (.I0(n2642), .I1(n6690), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4636));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1759_3_lut_3_lut (.I0(n2642), .I1(n6691), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1760_3_lut_3_lut (.I0(n2642), .I1(n6692), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4786));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_15_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4635));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4682));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4681));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1761_3_lut_3_lut (.I0(n2642), .I1(n6693), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1762_3_lut_3_lut (.I0(n2642), .I1(n6694), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1775_3_lut_3_lut (.I0(n2642), .I1(n6707), .I2(n530), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1764_3_lut_3_lut (.I0(n2642), .I1(n6696), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1765_3_lut_3_lut (.I0(n2642), .I1(n6697), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4680));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_i1767_3_lut_3_lut (.I0(n2642), .I1(n6699), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1766_3_lut_3_lut (.I0(n2642), .I1(n6698), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1773_3_lut_3_lut (.I0(n2642), .I1(n6705), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1774_3_lut_3_lut (.I0(n2642), .I1(n6706), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1771_3_lut_3_lut (.I0(n2642), .I1(n6703), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1763_3_lut_3_lut (.I0(n2642), .I1(n6695), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1772_3_lut_3_lut (.I0(n2642), .I1(n6704), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1768_3_lut_3_lut (.I0(n2642), .I1(n6700), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_i1770_3_lut_3_lut (.I0(n2642), .I1(n6702), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_15_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4679));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4678));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4677));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4676));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_87_i1_3_lut (.I0(pwm[3]), .I1(color[3]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[0]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4675));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4674));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4673));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4672));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39169_3_lut_4_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(pwm_count[2]), .O(n47071));   // verilog/motorControl.v(86[28:44])
    defparam i39169_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_15_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4671));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4670));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4669));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4668));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_634_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(GND_net), .O(n6_adj_4631));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_634_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_15_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4667));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4666));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4665));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39177_3_lut_4_lut (.I0(pwm_count[3]), .I1(pwm[3]), .I2(pwm[2]), 
            .I3(pwm_count[2]), .O(n47079));   // verilog/motorControl.v(65[19:32])
    defparam i39177_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_15_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4664));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4663));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_631_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(pwm[3]), 
            .I2(pwm[2]), .I3(GND_net), .O(n6_adj_4622));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_631_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_15_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4662));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_87_i2_3_lut (.I0(pwm[4]), .I1(color[4]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[1]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i3_3_lut (.I0(pwm[5]), .I1(color[5]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[2]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i4_3_lut (.I0(pwm[6]), .I1(color[6]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[3]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i5_3_lut (.I0(pwm[7]), .I1(color[7]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[4]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i6_3_lut (.I0(pwm[8]), .I1(color[8]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[5]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i7_3_lut (.I0(pwm[9]), .I1(color[9]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[6]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i8_3_lut (.I0(pwm[10]), .I1(color[10]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[7]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i9_3_lut (.I0(pwm[11]), .I1(color[11]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[8]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i10_3_lut (.I0(pwm[12]), .I1(color[12]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[9]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i11_3_lut (.I0(pwm[13]), .I1(color[13]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[10]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i12_3_lut (.I0(pwm[14]), .I1(color[14]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[11]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i13_3_lut (.I0(pwm[15]), .I1(color[15]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[12]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i14_3_lut (.I0(pwm[16]), .I1(color[16]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[13]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i15_3_lut (.I0(pwm[17]), .I1(color[17]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[14]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i16_3_lut (.I0(pwm[18]), .I1(color[18]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[15]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_87_i17_3_lut (.I0(pwm[19]), .I1(color[19]), .I2(pwm[23]), 
            .I3(GND_net), .O(color_23__N_1[16]));   // verilog/TinyFPGA_B.v(47[14] 49[8])
    defparam mux_87_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_15_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4661));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38835_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n46737));
    defparam i38835_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_15_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4660));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_15_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4659));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    motorControl control (.GND_net(GND_net), .deadband({deadband}), .\Kp[4] (Kp[4]), 
            .\PID_CONTROLLER.err[21] (\PID_CONTROLLER.err [21]), .\pwm_23__N_3310[10] (pwm_23__N_3310[10]), 
            .\pwm_23__N_3310[6] (pwm_23__N_3310[6]), .\pwm_23__N_3310[4] (pwm_23__N_3310[4]), 
            .PWMLimit({PWMLimit}), .\PID_CONTROLLER.result[19] (\PID_CONTROLLER.result [19]), 
            .n18644(n18644), .pwm({pwm}), .clk32MHz(clk32MHz), .n18643(n18643), 
            .n18642(n18642), .n18641(n18641), .n18639(n18639), .n18637(n18637), 
            .n18636(n18636), .n18635(n18635), .n18633(n18633), .n18632(n18632), 
            .\PID_CONTROLLER.err[23] (\PID_CONTROLLER.err [23]), .n18630(n18630), 
            .n18629(n18629), .n18628(n18628), .n18626(n18626), .n18624(n18624), 
            .n18623(n18623), .n18622(n18622), .\PID_CONTROLLER.result[17] (\PID_CONTROLLER.result [17]), 
            .\Kp[5] (Kp[5]), .n18574(n18574), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .n21(n21_adj_4613), .n9(n9_adj_4611), .\PID_CONTROLLER.err[31] (\PID_CONTROLLER.err [31]), 
            .n27(n27_adj_4614), .n13(n13_adj_4612), .\Kp[1] (Kp[1]), .\PID_CONTROLLER.err[22] (\PID_CONTROLLER.err [22]), 
            .\Kp[0] (Kp[0]), .n18495(n18495), .\PID_CONTROLLER.err_prev[31] (\PID_CONTROLLER.err_prev [31]), 
            .n18494(n18494), .\PID_CONTROLLER.err_prev[23] (\PID_CONTROLLER.err_prev [23]), 
            .n18493(n18493), .\PID_CONTROLLER.err_prev[22] (\PID_CONTROLLER.err_prev [22]), 
            .n18492(n18492), .\PID_CONTROLLER.err_prev[21] (\PID_CONTROLLER.err_prev [21]), 
            .n18491(n18491), .\PID_CONTROLLER.err_prev[20] (\PID_CONTROLLER.err_prev [20]), 
            .n18490(n18490), .\PID_CONTROLLER.err_prev[19] (\PID_CONTROLLER.err_prev [19]), 
            .n18489(n18489), .\PID_CONTROLLER.err_prev[18] (\PID_CONTROLLER.err_prev [18]), 
            .n18488(n18488), .\PID_CONTROLLER.err_prev[17] (\PID_CONTROLLER.err_prev [17]), 
            .n18487(n18487), .\PID_CONTROLLER.err_prev[16] (\PID_CONTROLLER.err_prev [16]), 
            .n18486(n18486), .\PID_CONTROLLER.err_prev[15] (\PID_CONTROLLER.err_prev [15]), 
            .n18485(n18485), .\PID_CONTROLLER.err_prev[14] (\PID_CONTROLLER.err_prev [14]), 
            .n18484(n18484), .\PID_CONTROLLER.err_prev[13] (\PID_CONTROLLER.err_prev [13]), 
            .n18483(n18483), .\PID_CONTROLLER.err_prev[12] (\PID_CONTROLLER.err_prev [12]), 
            .n18482(n18482), .\PID_CONTROLLER.err_prev[11] (\PID_CONTROLLER.err_prev [11]), 
            .n18481(n18481), .\PID_CONTROLLER.err_prev[10] (\PID_CONTROLLER.err_prev [10]), 
            .n18480(n18480), .\PID_CONTROLLER.err_prev[9] (\PID_CONTROLLER.err_prev [9]), 
            .n18479(n18479), .\PID_CONTROLLER.err_prev[8] (\PID_CONTROLLER.err_prev [8]), 
            .n18478(n18478), .\PID_CONTROLLER.err_prev[7] (\PID_CONTROLLER.err_prev [7]), 
            .n18477(n18477), .\PID_CONTROLLER.err_prev[6] (\PID_CONTROLLER.err_prev [6]), 
            .n18476(n18476), .\PID_CONTROLLER.err_prev[5] (\PID_CONTROLLER.err_prev [5]), 
            .n18475(n18475), .\PID_CONTROLLER.err_prev[4] (\PID_CONTROLLER.err_prev [4]), 
            .n18474(n18474), .\PID_CONTROLLER.err_prev[3] (\PID_CONTROLLER.err_prev [3]), 
            .n18473(n18473), .\PID_CONTROLLER.err_prev[2] (\PID_CONTROLLER.err_prev [2]), 
            .n18472(n18472), .\PID_CONTROLLER.err_prev[1] (\PID_CONTROLLER.err_prev [1]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\PID_CONTROLLER.result[10] (\PID_CONTROLLER.result [10]), 
            .\PID_CONTROLLER.result[13] (\PID_CONTROLLER.result [13]), .n387(n387), 
            .n21_adj_1(n21_adj_4607), .\Kd[1] (Kd[1]), .n9_adj_2(n9_adj_4605), 
            .\Kd[0] (Kd[0]), .\Kd[2] (Kd[2]), .\Ki[0] (Ki[0]), .n27_adj_3(n27), 
            .n13_adj_4(n13_adj_4606), .\Kd[3] (Kd[3]), .\Ki[1] (Ki[1]), 
            .n35(n35), .\Kd[4] (Kd[4]), .n39(n39), .\Kd[5] (Kd[5]), 
            .\Ki[2] (Ki[2]), .\PID_CONTROLLER.err[0] (\PID_CONTROLLER.err [0]), 
            .PIN_7_c_1(PIN_7_c_1), .PIN_6_c_0(PIN_6_c_0), .n22(n22_adj_4610), 
            .\Kd[6] (Kd[6]), .\Ki[3] (Ki[3]), .\Kd[7] (Kd[7]), .VCC_net(VCC_net), 
            .n853(n853), .GATES_5__N_3405(GATES_5__N_3405), .n44276(n44276), 
            .n855(n855), .n856(n856), .\Ki[4] (Ki[4]), .n857(n857), 
            .pwm_23__N_3307(pwm_23__N_3307), .n859(n859), .n860(n860), 
            .n861(n861), .n862(n862), .n863(n863), .n864(n864), .n865(n865), 
            .n866(n866), .n867(n867), .n868(n868), .n869(n869), .n870(n870), 
            .n871(n871), .n872(n872), .n873(n873), .n874(n874), .n875(n875), 
            .n46548(n46548), .\Ki[5] (Ki[5]), .n448(n448), .n449(n449), 
            .n450(n450), .n451(n451), .n453(n453), .n455(n455), .n456(n456), 
            .\PID_CONTROLLER.err[1] (\PID_CONTROLLER.err [1]), .\PID_CONTROLLER.err[2] (\PID_CONTROLLER.err [2]), 
            .\Ki[6] (Ki[6]), .n457(n457), .\PID_CONTROLLER.err[9] (\PID_CONTROLLER.err [9]), 
            .\Ki[7] (Ki[7]), .n459(n459), .n460(n460), .n462(n462), 
            .n463(n463), .n464(n464), .\PID_CONTROLLER.err[5] (\PID_CONTROLLER.err [5]), 
            .\PID_CONTROLLER.result[6] (\PID_CONTROLLER.result [6]), .n466(n466), 
            .\PID_CONTROLLER.result[4] (\PID_CONTROLLER.result [4]), .n468(n468), 
            .n469(n469), .n470(n470), .n471(n471), .n27_adj_5(n27_adj_4618), 
            .n13_adj_6(n13_adj_4616), .n414(n414), .n403(n403), .n35_adj_7(n35_adj_4619), 
            .n9_adj_8(n9_adj_4615), .n21_adj_9(n21_adj_4617), .n410(n410), 
            .n416(n416), .n401(n401), .pwm_count({pwm_count}), .n407(n407), 
            .n39_adj_10(n39_adj_4620), .\PID_CONTROLLER.err[6] (\PID_CONTROLLER.err [6]), 
            .\PID_CONTROLLER.err[7] (\PID_CONTROLLER.err [7]), .\PID_CONTROLLER.err[3] (\PID_CONTROLLER.err [3]), 
            .\PID_CONTROLLER.err[8] (\PID_CONTROLLER.err [8]), .\PID_CONTROLLER.err[4] (\PID_CONTROLLER.err [4]), 
            .hall1(hall1), .hall2(hall2), .\GATES_5__N_3398[5] (GATES_5__N_3398[5]), 
            .hall3(hall3), .n48474(n48474), .\PID_CONTROLLER.err_prev[0] (\PID_CONTROLLER.err_prev [0]), 
            .n25(n25_adj_4970), .n30(n30_adj_4967), .n26(n26_adj_4969), 
            .PIN_8_c_2(PIN_8_c_2), .PIN_9_c_3(PIN_9_c_3), .PIN_10_c_4(PIN_10_c_4), 
            .PIN_11_c_5(PIN_11_c_5), .\PID_CONTROLLER.err[10] (\PID_CONTROLLER.err [10]), 
            .\PID_CONTROLLER.err[11] (\PID_CONTROLLER.err [11]), .\PID_CONTROLLER.err[12] (\PID_CONTROLLER.err [12]), 
            .\PID_CONTROLLER.err[13] (\PID_CONTROLLER.err [13]), .\PID_CONTROLLER.err[14] (\PID_CONTROLLER.err [14]), 
            .\PID_CONTROLLER.err[15] (\PID_CONTROLLER.err [15]), .\PID_CONTROLLER.err[16] (\PID_CONTROLLER.err [16]), 
            .\PID_CONTROLLER.err[17] (\PID_CONTROLLER.err [17]), .\PID_CONTROLLER.err[18] (\PID_CONTROLLER.err [18]), 
            .\PID_CONTROLLER.err[19] (\PID_CONTROLLER.err [19]), .\PID_CONTROLLER.err[20] (\PID_CONTROLLER.err [20]), 
            .\motor_state[23] (motor_state[23]), .\motor_state[22] (motor_state[22]), 
            .\motor_state[21] (motor_state[21]), .\motor_state[20] (motor_state[20]), 
            .\motor_state[19] (motor_state[19]), .\motor_state[18] (motor_state[18]), 
            .\motor_state[17] (motor_state[17]), .\motor_state[16] (motor_state[16]), 
            .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .\motor_state[11] (motor_state[11]), .\motor_state[10] (motor_state[10]), 
            .\motor_state[9] (motor_state[9]), .\motor_state[8] (motor_state[8]), 
            .\motor_state[7] (motor_state[7]), .\motor_state[6] (motor_state[6]), 
            .\motor_state[5] (motor_state[5]), .\motor_state[4] (motor_state[4]), 
            .\motor_state[3] (motor_state[3]), .\motor_state[2] (motor_state[2]), 
            .\motor_state[1] (motor_state[1]), .\motor_state[0] (motor_state[0]), 
            .n17967(n17967), .n43362(n43362), .n13_adj_11(n13_adj_4609), 
            .n9_adj_12(n9_adj_4608), .IntegralLimit({IntegralLimit}), .setpoint({setpoint}), 
            .n16(n16_adj_4634), .n5(n5_adj_4984), .n29(n29_adj_4563)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(161[16] 177[4])
    SB_LUT4 div_15_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4788));   // verilog/TinyFPGA_B.v(180[21:53])
    defparam div_15_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (clk32MHz, timer, bit_ctr, VCC_net, n40240, n40236, 
            n40232, n40228, n40224, n40220, n46646, GND_net, n41781, 
            n40216, n40212, n40208, n40204, n40200, n40196, n46634, 
            n40192, n40188, n40184, n40180, n40176, n40172, n40168, 
            n40164, n40160, n40156, n40152, n40148, n40144, n40140, 
            n40136, n40132, n18698, \neo_pixel_transmitter.t0 , n18697, 
            n18696, n18695, n18694, n18693, n18692, n18691, n18690, 
            n18689, n18688, n18687, n18686, n18685, n18684, n18683, 
            n18682, n18681, n18680, n18679, n18678, n18677, n18676, 
            n18675, n18674, n18673, n18672, n18671, n18670, n18669, 
            n18668, n40242, start, n40116, n18552, \state[1] , n40120, 
            n40124, n40128, n46645, \state[0] , n46644, n46633, 
            n46643, n35, n46642, n29, \state_3__N_248[1] , n16572, 
            n20911, n43079, n46632, n46641, n46631, n46640, n46639, 
            n46630, n17665, n17802, n46629, n46659, n46658, n46638, 
            n46657, n46656, n46655, n46654, n46637, n46653, n17984, 
            n46652, n46651, n46636, n46650, n46628, PIN_14_c, n46649, 
            n46635, n46648, n46647, n17574, \color[2] , \color[3] , 
            n4, n43650, \color[1] , \color[0] , \color[6] , \color[7] , 
            \color[5] , \color[4] , \color[10] , \color[11] , \color[9] , 
            \color[8] , \color[18] , \color[19] , \color[17] , \color[16] , 
            \color[14] , \color[15] , \color[13] , \color[12] ) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    output [31:0]timer;
    output [31:0]bit_ctr;
    input VCC_net;
    input n40240;
    input n40236;
    input n40232;
    input n40228;
    input n40224;
    input n40220;
    output n46646;
    input GND_net;
    input n41781;
    input n40216;
    input n40212;
    input n40208;
    input n40204;
    input n40200;
    input n40196;
    output n46634;
    input n40192;
    input n40188;
    input n40184;
    input n40180;
    input n40176;
    input n40172;
    input n40168;
    input n40164;
    input n40160;
    input n40156;
    input n40152;
    input n40148;
    input n40144;
    input n40140;
    input n40136;
    input n40132;
    input n18698;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n18697;
    input n18696;
    input n18695;
    input n18694;
    input n18693;
    input n18692;
    input n18691;
    input n18690;
    input n18689;
    input n18688;
    input n18687;
    input n18686;
    input n18685;
    input n18684;
    input n18683;
    input n18682;
    input n18681;
    input n18680;
    input n18679;
    input n18678;
    input n18677;
    input n18676;
    input n18675;
    input n18674;
    input n18673;
    input n18672;
    input n18671;
    input n18670;
    input n18669;
    input n18668;
    input n40242;
    output start;
    input n40116;
    input n18552;
    output \state[1] ;
    input n40120;
    input n40124;
    input n40128;
    output n46645;
    output \state[0] ;
    output n46644;
    output n46633;
    output n46643;
    output n35;
    output n46642;
    output n29;
    output \state_3__N_248[1] ;
    output n16572;
    output n20911;
    output n43079;
    output n46632;
    output n46641;
    output n46631;
    output n46640;
    output n46639;
    output n46630;
    output n17665;
    output n17802;
    output n46629;
    output n46659;
    output n46658;
    output n46638;
    output n46657;
    output n46656;
    output n46655;
    output n46654;
    output n46637;
    output n46653;
    input n17984;
    output n46652;
    output n46651;
    output n46636;
    output n46650;
    output n46628;
    output PIN_14_c;
    output n46649;
    output n46635;
    output n46648;
    output n46647;
    output n17574;
    input \color[2] ;
    input \color[3] ;
    output n4;
    output n43650;
    input \color[1] ;
    input \color[0] ;
    input \color[6] ;
    input \color[7] ;
    input \color[5] ;
    input \color[4] ;
    input \color[10] ;
    input \color[11] ;
    input \color[9] ;
    input \color[8] ;
    input \color[18] ;
    input \color[19] ;
    input \color[17] ;
    input \color[16] ;
    input \color[14] ;
    input \color[15] ;
    input \color[13] ;
    input \color[12] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2991, n2892, n2918, n34980, n34981, \neo_pixel_transmitter.done_N_456 , 
        n49991, \neo_pixel_transmitter.done , n2992, n2893, n34979, 
        n2993, n2894, n34978, n2994, n2895, n34977, n2995, n2896, 
        n34976, n2996, n2897, n34975, n2997, n2898, n34974, n2998, 
        n2899, n34973, n2999, n2900, n34972, n3000, n2901, n34971, 
        n3001, n2902, n34970, n3002, n2903, n34969, n22;
    wire [31:0]n51;
    
    wire n34796;
    wire [31:0]one_wire_N_399;
    
    wire n3003, n2904, n34968, n29_c, n34795, n3004, n2905, n34967, 
        n3005, n2906, n34966, n3006, n2907, n34965, n23, n34794, 
        n3007, n2908, n34964, n3008, n2909, n49781, n34963, n30, 
        n34793, n3009, n21, n34792, n34533, n34791, n25, n34790, 
        n26, n34789, n28, n34788, n34787, n34786, n27, n34785, 
        n34784, n34521, n34783, n24, n34782, n34781, n1409, n26058, 
        n1405, n1403, n1406, n16_adj_4424, n1402, n1404, n1400, 
        n1407, n17_adj_4425, n1408, n1401, n1433, n3083, n2984, 
        n3017, n34951, n1334, n49789, n3084, n2985, n34950, n1304, 
        n1305, n10_adj_4426, n1303, n1309, n12_adj_4427, n1306, 
        n1308, n1302, n16_adj_4428, n1307, n1301, n1235, n49788, 
        n1205, n1206, n1204, n1207, n14_adj_4429, n1203, n1209, 
        n9_adj_4430, n1202, n1208, n1136, n49787, n1109, n26064, 
        n1105, n1103, n1108, n12_adj_4431, n1107, n1106, n1104, 
        n1037, n49786, n38183;
    wire [31:0]n971;
    
    wire n1007, n3085, n2986, n34949, n1006, n906, n1005, n905, 
        n42682, n44306, n34780, n17743, n15226, n1009, n1008, 
        n44322, n6_adj_4432, n4_adj_4433, n3086, n2987, n34948, 
        n34779, n3087, n2988, n34947, n3088, n2989, n34946, n3089, 
        n2990, n34945, n838, n3090, n34944, n3091, n34943, n34778, 
        n34777, n3092, n34942, n3093, n34941, n34776, n3094, n34940, 
        n3095, n34939, n34775, n2588, n2489, n2522, n35246, n3096, 
        n34938, n34774, n2589, n2490, n35245, n34773, n2590, n2491, 
        n35244, n3097, n34937, n34772, n2591, n2492, n35243, n34771, 
        n2592, n2493, n35242, n3098, n34936, n34770, n2593, n2494, 
        n35241, n3099, n34935, n34769, n2594, n2495, n35240, n3100, 
        n34934, n34768, n2595, n2496, n35239, n34767, n2596, n2497, 
        n35238, n3101, n34933, n2597, n2498, n35237, n3102, n34932, 
        n120, n34766, n2598, n2499, n35236, n2599, n2500, n35235, 
        n3103, n34931, n3104, n34930, n2600, n2501, n35234, n3105, 
        n34929, n2601, n2502, n35233, n3106, n34928, n34534, n2602, 
        n2503, n35232, n2603, n2504, n35231, n3107, n34927, n2604, 
        n2505, n35230, n2605, n2506, n35229, n2606, n2507, n35228, 
        n3108, n49782, n34926, n3109, n34532, n34522, n807, n60, 
        n2607, n2508, n35227, n3182, n3116, n34925, n2608, n2509, 
        n49783, n35226, n2609, n3183, n34924, n3184, n34923, n3185, 
        n34922, n3186, n34921, n3187, n34920, n608, n3188, n34919, 
        n3189, n34918, n708, n42547, n26074, n739, n3190, n34917, 
        n15228, n3191, n34916, n3192, n34915, n37493, n42530, 
        n3193, n34914, n3194, n34913, n3195, n34912, n3196, n34911, 
        n3197, n34910, n3198, n34909, n3199, n34908, n3200, n34907, 
        n3201, n34906, n3202, n34905, n3203, n34904, n3204, n34903, 
        n3205, n34902, n3206, n34901, n3207, n34900;
    wire [31:0]n133;
    
    wire n3208, n49784, n34899, n3209, n42660, n42605, n36, n37, 
        n16583, n92, n121, n41871, n4_adj_4444, n43103, n14_adj_4445, 
        n7_adj_4446, n34531, n34520, n35633, n35632, n35631, n35630, 
        n35629, n35628, n35627, n35626, n35625, n35624, n35623, 
        n35622, n35621, n35620, n35619, n35618, n34530, n35617, 
        n35616, n35615, n35614, n35613, n35612, n35611, n35610, 
        n35609, n35608, n35607, n35606, n35605, n35604, n35603, 
        n35602, n35601, n35600, n35599, n42, n94, n92_adj_4447, 
        n42563, n6_adj_4448, n1499, n35598, n1500, n35597, n1501, 
        n35596, n1502, n35595, n1503, n35594, n1504, n35593, n1505, 
        n35592, n1506, n35591, n1507, n35590, n1508, n49790, n35589, 
        n1509, n2687, n2621, n35140, n2688, n35139, n2887, n26_adj_4449, 
        n2888, n42_adj_4450, n2886, n40, n2890, n2889, n41, n2891, 
        n39, n36_adj_4451, n44, n48, n2885, n35_adj_4452, n2689, 
        n35138, n2690, n35137, n2691, n35136, n2692, n35135, n2693, 
        n35134, n34529, n2694, n35133, n2695, n35132, n2696, n35131, 
        n2697, n35130, n2698, n35129, n2699, n35128, n2700, n35127, 
        n2701, n35126, n2702, n35125, n2703, n35124, n2704, n35123, 
        n1598, n1532, n35542, n2705, n35122, n2706, n35121, n1599, 
        n35541, n2707, n35120, n1600, n35540, n1601, n35539, n2708, 
        n49791, n35119, n1602, n35538, n2709, n1603, n35537, n1604, 
        n35536, n1605, n35535, n1606, n35534, n1607, n35533, n1608, 
        n49792, n35532, n1609, n1697, n1631, n35531, n1698, n35530, 
        n1699, n35529, n1700, n35528, n1701, n35527, n1702, n35526, 
        n1703, n35525, n1704, n35524, n1705, n35523, n1706, n35522, 
        n6_adj_4453, n1, n128, n1707, n35521, n1708, n49793, n35520, 
        n30_adj_4455, n48_adj_4456, n46, n47, n45, n1709, n44_adj_4457, 
        n43, n54, n49, n4434, n42_adj_4458, n46_adj_4459, n44_adj_4460, 
        n45_adj_4461, n43_adj_4462, n40_adj_4463, n48_adj_4464, n52, 
        n39_adj_4465, n1796, n1730, n35510, n1797, n35509, n1798, 
        n35508, n1799, n35507, n24_adj_4466, n34, n22_adj_4467, 
        n38, n36_adj_4468, n37_adj_4469, n35_adj_4470, n1800, n35506, 
        n34519, n1801, n35505, n1802, n35504, n1803, n35503, n1804, 
        n35502, n1805, n35501, n1806, n35500, n1807, n35499, n1808, 
        n49794, n35498, n1809, n1895, n1829, n35483, n1896, n35482, 
        n1897, n35481, n1898, n35480, n1899, n35479, n1900, n35478, 
        n1901, n35477, n1902, n35476, n1903, n35475, n1904, n35474, 
        n1905, n35473, n1906, n35472, n1907, n35471, n1908, n49795, 
        n35470, n1909, n1994, n1928, n35469, n1995, n35468, n1996, 
        n35467, n1997, n35466, n2786, n2720, n35079, n1998, n35465, 
        n2787, n35078, n1999, n35464, n2000, n35463, n2788, n35077, 
        n2001, n35462, n2002, n35461, n2789, n35076, n2003, n35460, 
        n2004, n35459, n2790, n35075, n2005, n35458, n2006, n35457, 
        n2791, n35074, n2007, n35456, n2008, n49796, n35455, n2792, 
        n35073, n2009, n2093, n2027, n35454, n2094, n35453, n2793, 
        n35072, n2095, n35452, n2096, n35451, n2794, n35071, n2097, 
        n35450, n2098, n35449, n2795, n35070, n2099, n35448, n2796, 
        n35069, n2100, n35447, n2101, n35446, n2797, n35068, n2102, 
        n35445, n2103, n35444, n2798, n35067, n2104, n35443, n2105, 
        n35442, n2799, n35066, n2106, n35441, n2107, n35440, n2800, 
        n35065, n2108, n49798, n35439, n2109, n2801, n35064, n2192, 
        n2126, n35438, n2193, n35437, n2194, n35436, n2802, n35063, 
        n2803, n35062, n2195, n35435, n2196, n35434, n2197, n35433, 
        n2804, n35061, n2805, n35060, n2806, n35059, n2198, n35432, 
        n2199, n35431, n2807, n35058, n2200, n35430, n2808, n49797, 
        n35057, n2201, n35429, n34528, n2202, n35428, n2809, n2203, 
        n35427, n2204, n35426, n34518, n2205, n35425, n2206, n35424, 
        n2207, n35423, n2208, n49799, n35422, n2209, n2291, n2225, 
        n35421, n2292, n35420, n2293, n35419, n2294, n35418, n2295, 
        n35417, n2296, n35416, n2297, n35415, n2298, n35414, n2299, 
        n35413, n34527, n2300, n35412, n2301, n35411, n2302, n35410, 
        n2303, n35409, n2304, n35408, n2305, n35407, n2306, n35406, 
        n2307, n35405, n2308, n49800, n35404, n2309, n2390, n2324, 
        n35403, n2391, n35402, n2392, n35401, n2393, n35400, n2394, 
        n35399, n2819, n35026, n34526, n35025, n2395, n35398, 
        n35024, n34517, n2396, n35397, n35023, n2397, n35396, 
        n35022, n2398, n35395, n35021, n35020, n2399, n35394, 
        n35019, n35018, n2400, n35393, n2401, n35392, n35017, 
        n2402, n35391, n35016, n35015, n2403, n35390, n2404, n35389, 
        n35014, n2405, n35388, n35013, n2406, n35387, n35012, 
        n2407, n35386, n2408, n49801, n35385, n35011, n2409, n35010, 
        n35384, n35383, n35009, n35382, n35008, n35007, n35381;
    wire [3:0]state_3__N_248;
    
    wire n34516, n35380, n35006, n35379, n35378, n35005, n34546, 
        n35004, n35377, n34545, n35376, n35375, n49802, n35003, 
        n35374, n34525, n35373, n35372, n34544, n35371, n35370, 
        n35369, n34543, n35368, n35367, n34542, n35366, n35365, 
        n35364, n35363, n35362, n35361, n34541, n35360, n35359, 
        n35358, n34524, n35357, n35356, n34540, n35355, n35354, 
        n2423, n35353, n35352, n35351, n35350, n35349, n35348, 
        n35347, n35346, n35345, n35344, n35343, n35342, n35341, 
        n35340, n35339, n35338, n35337, n34539, n34538, n35336, 
        n35335, n34523, n49803, n35334, n34987, n34537, \neo_pixel_transmitter.done_N_462 , 
        n17611, n44172, n34536, n34986, n34985, n34535, n34984, 
        n34983, n34982, n26050, n852, n41777, n20959, n11_adj_4471, 
        n40_adj_4472, n44_adj_4473, n42_adj_4474, n43_adj_4475, n41_adj_4476, 
        n38_adj_4477, n46_adj_4478, n49907, n50, n37_adj_4479, n26090;
    wire [4:0]color_bit_N_442;
    
    wire n42557, n41814, n60_adj_4480, n4_adj_4481, n54_adj_4482, 
        n116, n57, n27_adj_4484, n33_adj_4485, n32_adj_4486, n31_adj_4487, 
        n35_adj_4488, n37_adj_4489, n44398, n25994, n48_adj_4490, 
        n46_adj_4491, n47_adj_4492, n45_adj_4493, n44_adj_4494, n43_adj_4495, 
        n54_adj_4496, n49_adj_4497, n49868, n46586, n49808, n40_adj_4498, 
        n38_adj_4499, n39_adj_4500, n37_adj_4501, n34_adj_4502, n42_adj_4503, 
        n46_adj_4504, n33_adj_4505, n25936, n30_adj_4506, n34_adj_4507, 
        n32_adj_4508, n33_adj_4509, n31_adj_4510, n28_adj_4511, n32_adj_4512, 
        n30_adj_4513, n31_adj_4514, n29_adj_4515, n18_adj_4516, n25927, 
        n30_adj_4517, n28_adj_4518, n29_adj_4519, n27_adj_4520, n49901, 
        n44401, n18_adj_4521, n28_adj_4522, n26_adj_4523, n27_adj_4524, 
        n25_adj_4525, n36_adj_4526, n40_adj_4527, n31_adj_4528, n38_adj_4529, 
        n37_adj_4530, n41_adj_4531, n43_adj_4532, n26_adj_4533, n24_adj_4534, 
        n25_adj_4535, n23_adj_4536, n24_adj_4537, n22_adj_4538, n23_adj_4539, 
        n21_adj_4540, n49895, n44404, n49865, n22_adj_4541, n20_adj_4542, 
        n21_adj_4543, n19_adj_4544, n49829, n48564, n20_adj_4545, 
        n13_adj_4546, n18_adj_4547, n22_adj_4548, n18_adj_4549, n20_adj_4550, 
        n15_adj_4551, n49805, n36_adj_4552, n25_adj_4553, n34_adj_4554, 
        n40_adj_4555, n38_adj_4556, n39_adj_4557, n37_adj_4558;
    
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n34980), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n34980), .I0(n2892), .I1(n2918), .CO(n34981));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n49991), .D(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n34979), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n34979), .I0(n2893), .I1(n2918), .CO(n34980));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n34978), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n34978), .I0(n2894), .I1(n2918), .CO(n34979));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n34977), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n34977), .I0(n2895), .I1(n2918), .CO(n34978));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n34976), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n34976), .I0(n2896), .I1(n2918), .CO(n34977));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n34975), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n34975), .I0(n2897), .I1(n2918), .CO(n34976));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n34974), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n34974), .I0(n2898), .I1(n2918), .CO(n34975));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n34973), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n34973), .I0(n2899), .I1(n2918), .CO(n34974));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n34972), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n34972), .I0(n2900), .I1(n2918), .CO(n34973));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n34971), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n34971), .I0(n2901), .I1(n2918), .CO(n34972));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n34970), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n34970), .I0(n2902), .I1(n2918), .CO(n34971));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n34969), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n34969), .I0(n2903), .I1(n2918), .CO(n34970));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_399[22]), .I1(timer[31]), 
            .I2(n51[31]), .I3(n34796), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n34968), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_399[16]), .I1(timer[30]), 
            .I2(n51[30]), .I3(n34795), .O(n29_c)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n34795), .I0(timer[30]), .I1(n51[30]), 
            .CO(n34796));
    SB_CARRY mod_5_add_2009_8 (.CI(n34968), .I0(n2904), .I1(n2918), .CO(n34969));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n34967), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n34967), .I0(n2905), .I1(n2918), .CO(n34968));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n34966), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n34966), .I0(n2906), .I1(n2918), .CO(n34967));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n34965), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_399[19]), .I1(timer[29]), 
            .I2(n51[29]), .I3(n34794), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_5 (.CI(n34965), .I0(n2907), .I1(n2918), .CO(n34966));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n34964), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_31 (.CI(n34794), .I0(timer[29]), .I1(n51[29]), 
            .CO(n34795));
    SB_CARRY mod_5_add_2009_4 (.CI(n34964), .I0(n2908), .I1(n2918), .CO(n34965));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n49781), 
            .I3(n34963), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_399[26]), .I1(timer[28]), 
            .I2(n51[28]), .I3(n34793), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_3 (.CI(n34963), .I0(n2909), .I1(n49781), .CO(n34964));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n49781), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_30 (.CI(n34793), .I0(timer[28]), .I1(n51[28]), 
            .CO(n34794));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n49781), 
            .CO(n34963));
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n40240));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n40236));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n40232));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_399[18]), .I1(timer[27]), 
            .I2(n51[27]), .I3(n34792), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n40228));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n40224));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n40220));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_29 (.CI(n34792), .I0(timer[27]), .I1(n51[27]), 
            .CO(n34793));
    SB_LUT4 add_21_20_lut (.I0(n41781), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n34533), .O(n46646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n40216));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n51[26]), 
            .I3(n34791), .O(one_wire_N_399[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n34791), .I0(timer[26]), .I1(n51[26]), 
            .CO(n34792));
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n40212));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_27_lut (.I0(one_wire_N_399[12]), .I1(timer[25]), 
            .I2(n51[25]), .I3(n34790), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n34790), .I0(timer[25]), .I1(n51[25]), 
            .CO(n34791));
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n40208));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_26_lut (.I0(one_wire_N_399[14]), .I1(timer[24]), 
            .I2(n51[24]), .I3(n34789), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n40204));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_26 (.CI(n34789), .I0(timer[24]), .I1(n51[24]), 
            .CO(n34790));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_399[21]), .I1(timer[23]), 
            .I2(n51[23]), .I3(n34788), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n34788), .I0(timer[23]), .I1(n51[23]), 
            .CO(n34789));
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n40200));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n40196));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n51[22]), 
            .I3(n34787), .O(one_wire_N_399[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_24 (.CI(n34787), .I0(timer[22]), .I1(n51[22]), 
            .CO(n34788));
    SB_LUT4 sub_14_add_2_23_lut (.I0(GND_net), .I1(timer[21]), .I2(n51[21]), 
            .I3(n34786), .O(one_wire_N_399[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_23 (.CI(n34786), .I0(timer[21]), .I1(n51[21]), 
            .CO(n34787));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_399[15]), .I1(timer[20]), 
            .I2(n51[20]), .I3(n34785), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n34785), .I0(timer[20]), .I1(n51[20]), 
            .CO(n34786));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n51[19]), 
            .I3(n34784), .O(one_wire_N_399[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_8_lut (.I0(n41781), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n34521), .O(n46634)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n40192));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n40188));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_21 (.CI(n34784), .I0(timer[19]), .I1(n51[19]), 
            .CO(n34785));
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n40184));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n51[18]), 
            .I3(n34783), .O(one_wire_N_399[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n34783), .I0(timer[18]), .I1(n51[18]), 
            .CO(n34784));
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n40180));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n40176));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n40172));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n40168));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n40164));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n40160));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n40156));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_399[13]), .I1(timer[17]), 
            .I2(n51[17]), .I3(n34782), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n40152));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n40148));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n40144));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n40140));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n40136));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n40132));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_19 (.CI(n34782), .I0(timer[17]), .I1(n51[17]), 
            .CO(n34783));
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n18698));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n18697));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n18696));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n18695));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n18694));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n18693));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n51[16]), 
            .I3(n34781), .O(one_wire_N_399[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20793_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n26058));
    defparam i20793_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n18692));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n18691));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i6_4_lut (.I0(n1405), .I1(n26058), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4424));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n18690));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n18689));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n18688));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n18687));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n18686));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n18685));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n18684));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i7_4_lut (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4425));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n18683));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n18682));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n18681));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i9_4_lut (.I0(n17_adj_4425), .I1(n1408), .I2(n16_adj_4424), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n18680));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n18679));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n18678));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n18677));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n18676));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n18675));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n18674));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n18673));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n18672));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n18671));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n18670));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n18669));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n18668));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n40242));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n40116));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n34951), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i41888_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49789));
    defparam i41888_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n18552));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(VCC_net), 
            .D(n40120));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(VCC_net), 
            .D(n40124));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(VCC_net), 
            .D(n40128));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n34950), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_18 (.CI(n34781), .I0(timer[16]), .I1(n51[16]), 
            .CO(n34782));
    SB_LUT4 i1_2_lut (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4426));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4427));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1428 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4426), 
            .O(n16_adj_4428));
    defparam i7_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16_adj_4428), .I2(n12_adj_4427), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_27 (.CI(n34950), .I0(n2985), .I1(n3017), .CO(n34951));
    SB_LUT4 i41887_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49788));
    defparam i41887_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1429 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4429));
    defparam i6_4_lut_adj_1429.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n9_adj_4430));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1430 (.I0(n9_adj_4430), .I1(n14_adj_4429), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1430.LUT_INIT = 16'hfffe;
    SB_LUT4 i41886_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49787));
    defparam i41886_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20799_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n26064));
    defparam i20799_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n26064), .I3(n1108), 
            .O(n12_adj_4431));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1431 (.I0(n1107), .I1(n12_adj_4431), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 i41885_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49786));
    defparam i41885_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i41867_2_lut (.I0(n38183), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i41867_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n34949), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i41869_2_lut (.I0(n38183), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i41869_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n38183), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36408_3_lut (.I0(n905), .I1(n906), .I2(n42682), .I3(GND_net), 
            .O(n44306));
    defparam i36408_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n51[15]), 
            .I3(n34780), .O(one_wire_N_399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n44306), .I2(n17743), .I3(n15226), 
            .O(n38183));
    defparam i4_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n38183), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n15226), .I1(n971[27]), .I2(n38183), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36422_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n44322));
    defparam i36422_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6_adj_4432));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY sub_14_add_2_17 (.CI(n34780), .I0(timer[15]), .I1(n51[15]), 
            .CO(n34781));
    SB_CARRY mod_5_add_2076_26 (.CI(n34949), .I0(n2986), .I1(n3017), .CO(n34950));
    SB_LUT4 i3_4_lut (.I0(n38183), .I1(n6_adj_4432), .I2(n1005), .I3(n44322), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i41865_2_lut (.I0(n38183), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4433));   // verilog/neopixel.v(22[26:36])
    defparam i41865_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n34948), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n51[14]), 
            .I3(n34779), .O(one_wire_N_399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_25 (.CI(n34948), .I0(n2987), .I1(n3017), .CO(n34949));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n34947), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n34947), .I0(n2988), .I1(n3017), .CO(n34948));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n34946), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n34946), .I0(n2989), .I1(n3017), .CO(n34947));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n34945), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n34945), .I0(n2990), .I1(n3017), .CO(n34946));
    SB_CARRY sub_14_add_2_16 (.CI(n34779), .I0(timer[14]), .I1(n51[14]), 
            .CO(n34780));
    SB_LUT4 i1_2_lut_adj_1432 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n15226));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n34944), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n34944), .I0(n2991), .I1(n3017), .CO(n34945));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n34943), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n51[13]), 
            .I3(n34778), .O(one_wire_N_399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n34778), .I0(timer[13]), .I1(n51[13]), 
            .CO(n34779));
    SB_CARRY mod_5_add_2076_20 (.CI(n34943), .I0(n2992), .I1(n3017), .CO(n34944));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n51[12]), 
            .I3(n34777), .O(one_wire_N_399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n34942), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n34942), .I0(n2993), .I1(n3017), .CO(n34943));
    SB_CARRY sub_14_add_2_14 (.CI(n34777), .I0(timer[12]), .I1(n51[12]), 
            .CO(n34778));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n34941), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n34941), .I0(n2994), .I1(n3017), .CO(n34942));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n51[11]), 
            .I3(n34776), .O(one_wire_N_399[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n34940), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n34940), .I0(n2995), .I1(n3017), .CO(n34941));
    SB_CARRY sub_14_add_2_13 (.CI(n34776), .I0(timer[11]), .I1(n51[11]), 
            .CO(n34777));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n34939), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n34939), .I0(n2996), .I1(n3017), .CO(n34940));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n51[10]), 
            .I3(n34775), .O(one_wire_N_399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n35246), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n34938), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_12 (.CI(n34775), .I0(timer[10]), .I1(n51[10]), 
            .CO(n34776));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n51[9]), 
            .I3(n34774), .O(one_wire_N_399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n35245), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n35245), .I0(n2490), .I1(n2522), .CO(n35246));
    SB_CARRY mod_5_add_2076_15 (.CI(n34938), .I0(n2997), .I1(n3017), .CO(n34939));
    SB_CARRY sub_14_add_2_11 (.CI(n34774), .I0(timer[9]), .I1(n51[9]), 
            .CO(n34775));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n51[8]), 
            .I3(n34773), .O(one_wire_N_399[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n35244), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n35244), .I0(n2491), .I1(n2522), .CO(n35245));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n34937), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n34773), .I0(timer[8]), .I1(n51[8]), 
            .CO(n34774));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n51[7]), 
            .I3(n34772), .O(one_wire_N_399[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n35243), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n35243), .I0(n2492), .I1(n2522), .CO(n35244));
    SB_CARRY mod_5_add_2076_14 (.CI(n34937), .I0(n2998), .I1(n3017), .CO(n34938));
    SB_CARRY sub_14_add_2_9 (.CI(n34772), .I0(timer[7]), .I1(n51[7]), 
            .CO(n34773));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n51[6]), 
            .I3(n34771), .O(one_wire_N_399[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n35242), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n34936), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n35242), .I0(n2493), .I1(n2522), .CO(n35243));
    SB_CARRY mod_5_add_2076_13 (.CI(n34936), .I0(n2999), .I1(n3017), .CO(n34937));
    SB_CARRY sub_14_add_2_8 (.CI(n34771), .I0(timer[6]), .I1(n51[6]), 
            .CO(n34772));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n51[5]), 
            .I3(n34770), .O(one_wire_N_399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n35241), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n35241), .I0(n2494), .I1(n2522), .CO(n35242));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n34935), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_7 (.CI(n34770), .I0(timer[5]), .I1(n51[5]), 
            .CO(n34771));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n51[4]), 
            .I3(n34769), .O(one_wire_N_399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n35240), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n34935), .I0(n3000), .I1(n3017), .CO(n34936));
    SB_CARRY mod_5_add_1741_17 (.CI(n35240), .I0(n2495), .I1(n2522), .CO(n35241));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n34934), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_6 (.CI(n34769), .I0(timer[4]), .I1(n51[4]), 
            .CO(n34770));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n51[3]), 
            .I3(n34768), .O(one_wire_N_399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n35239), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_5 (.CI(n34768), .I0(timer[3]), .I1(n51[3]), 
            .CO(n34769));
    SB_CARRY mod_5_add_1741_16 (.CI(n35239), .I0(n2496), .I1(n2522), .CO(n35240));
    SB_CARRY mod_5_add_2076_11 (.CI(n34934), .I0(n3001), .I1(n3017), .CO(n34935));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n51[2]), 
            .I3(n34767), .O(one_wire_N_399[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n34767), .I0(timer[2]), .I1(n51[2]), 
            .CO(n34768));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n35238), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n34933), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n35238), .I0(n2497), .I1(n2522), .CO(n35239));
    SB_CARRY mod_5_add_2076_10 (.CI(n34933), .I0(n3002), .I1(n3017), .CO(n34934));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n35237), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n35237), .I0(n2498), .I1(n2522), .CO(n35238));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n34932), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_399[0]), .I1(timer[1]), .I2(n51[1]), 
            .I3(n34766), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_3 (.CI(n34766), .I0(timer[1]), .I1(n51[1]), 
            .CO(n34767));
    SB_LUT4 sub_14_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n51[0]), 
            .I3(VCC_net), .O(one_wire_N_399[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n35236), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n34932), .I0(n3003), .I1(n3017), .CO(n34933));
    SB_CARRY mod_5_add_1741_13 (.CI(n35236), .I0(n2499), .I1(n2522), .CO(n35237));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n35235), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n34931), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n51[0]), 
            .CO(n34766));
    SB_CARRY mod_5_add_2076_8 (.CI(n34931), .I0(n3004), .I1(n3017), .CO(n34932));
    SB_CARRY mod_5_add_1741_12 (.CI(n35235), .I0(n2500), .I1(n2522), .CO(n35236));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n34930), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n35234), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n34930), .I0(n3005), .I1(n3017), .CO(n34931));
    SB_CARRY mod_5_add_1741_11 (.CI(n35234), .I0(n2501), .I1(n2522), .CO(n35235));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n34929), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n34929), .I0(n3006), .I1(n3017), .CO(n34930));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n35233), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n34928), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n34533), .I0(bit_ctr[18]), .I1(GND_net), .CO(n34534));
    SB_CARRY mod_5_add_1741_10 (.CI(n35233), .I0(n2502), .I1(n2522), .CO(n35234));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n35232), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n35232), .I0(n2503), .I1(n2522), .CO(n35233));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n35231), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n35231), .I0(n2504), .I1(n2522), .CO(n35232));
    SB_CARRY mod_5_add_2076_5 (.CI(n34928), .I0(n3007), .I1(n3017), .CO(n34929));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n34927), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n34927), .I0(n3008), .I1(n3017), .CO(n34928));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n35230), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n35230), .I0(n2505), .I1(n2522), .CO(n35231));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n35229), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n35229), .I0(n2506), .I1(n2522), .CO(n35230));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n35228), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n49782), 
            .I3(n34926), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n34926), .I0(n3009), .I1(n49782), .CO(n34927));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n49782), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_19_lut (.I0(n41781), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n34532), .O(n46645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_8 (.CI(n34521), .I0(bit_ctr[6]), .I1(GND_net), .CO(n34522));
    SB_CARRY add_21_19 (.CI(n34532), .I0(bit_ctr[17]), .I1(GND_net), .CO(n34533));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n49782), 
            .CO(n34926));
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY mod_5_add_1741_5 (.CI(n35228), .I0(n2507), .I1(n2522), .CO(n35229));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n35227), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n34925), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n35227), .I0(n2508), .I1(n2522), .CO(n35228));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n49783), 
            .I3(n35226), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n35226), .I0(n2509), .I1(n49783), .CO(n35227));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n49783), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n34924), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n34924), .I0(n3084), .I1(n3116), .CO(n34925));
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n49783), 
            .CO(n35226));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n34923), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n34923), .I0(n3085), .I1(n3116), .CO(n34924));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n34922), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n34922), .I0(n3086), .I1(n3116), .CO(n34923));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n34921), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n34921), .I0(n3087), .I1(n3116), .CO(n34922));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n34920), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20753_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i20753_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_2143_24 (.CI(n34920), .I0(n3088), .I1(n3116), .CO(n34921));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n34919), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n34919), .I0(n3089), .I1(n3116), .CO(n34920));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n34918), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n34918), .I0(n3090), .I1(n3116), .CO(n34919));
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n42547), .I3(n26074), 
            .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n34917), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1433 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n15228));
    defparam i1_2_lut_adj_1433.LUT_INIT = 16'h6666;
    SB_CARRY mod_5_add_2143_21 (.CI(n34917), .I0(n3091), .I1(n3116), .CO(n34918));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n34916), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n34916), .I0(n3092), .I1(n3116), .CO(n34917));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n34915), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i39344_3_lut (.I0(n37493), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n42530));
    defparam i39344_3_lut.LUT_INIT = 16'ha6a6;
    SB_CARRY mod_5_add_2143_19 (.CI(n34915), .I0(n3093), .I1(n3116), .CO(n34916));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n34914), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n34914), .I0(n3094), .I1(n3116), .CO(n34915));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n34913), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n34913), .I0(n3095), .I1(n3116), .CO(n34914));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n34912), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n34912), .I0(n3096), .I1(n3116), .CO(n34913));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n34911), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n34911), .I0(n3097), .I1(n3116), .CO(n34912));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n34910), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n34910), .I0(n3098), .I1(n3116), .CO(n34911));
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n42547), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n34909), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n34909), .I0(n3099), .I1(n3116), .CO(n34910));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n34908), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n34908), .I0(n3100), .I1(n3116), .CO(n34909));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n34907), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n34907), .I0(n3101), .I1(n3116), .CO(n34908));
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n34906), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_4_lut (.I0(n42530), .I1(n15228), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_CARRY mod_5_add_2143_10 (.CI(n34906), .I0(n3102), .I1(n3116), .CO(n34907));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n34905), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n34905), .I0(n3103), .I1(n3116), .CO(n34906));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n34904), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n34904), .I0(n3104), .I1(n3116), .CO(n34905));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n34903), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i41177_3_lut_4_lut (.I0(n15228), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n42530), .O(n42682));   // verilog/neopixel.v(22[26:36])
    defparam i41177_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_CARRY mod_5_add_2143_7 (.CI(n34903), .I0(n3105), .I1(n3116), .CO(n34904));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n34902), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n34902), .I0(n3106), .I1(n3116), .CO(n34903));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n34901), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n34901), .I0(n3107), .I1(n3116), .CO(n34902));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n34900), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1189__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_2143_4 (.CI(n34900), .I0(n3108), .I1(n3116), .CO(n34901));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n49784), 
            .I3(n34899), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n34899), .I0(n3109), .I1(n49784), .CO(n34900));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n49784), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n49784), 
            .CO(n34899));
    SB_LUT4 i2_3_lut_adj_1434 (.I0(one_wire_N_399[6]), .I1(one_wire_N_399[5]), 
            .I2(one_wire_N_399[9]), .I3(GND_net), .O(n42660));
    defparam i2_3_lut_adj_1434.LUT_INIT = 16'hfefe;
    SB_LUT4 i34722_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n42605));
    defparam i34722_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut (.I0(n21), .I1(n23), .I2(n22), .I3(n24), .O(n36));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n37));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n29_c), .I2(n36), .I3(n30), .O(n16583));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1435 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n92));
    defparam i1_2_lut_adj_1435.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(one_wire_N_399[2]), .I1(n120), .I2(GND_net), 
            .I3(GND_net), .O(n121));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_399[2]), .I1(one_wire_N_399[3]), .I2(n41871), 
            .I3(one_wire_N_399[4]), .O(n4_adj_4444));
    defparam i1_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i2_4_lut_adj_1437 (.I0(one_wire_N_399[4]), .I1(n4_adj_4444), 
            .I2(n121), .I3(n41871), .O(n43103));
    defparam i2_4_lut_adj_1437.LUT_INIT = 16'hddcd;
    SB_LUT4 i6_4_lut_adj_1438 (.I0(n43103), .I1(one_wire_N_399[11]), .I2(one_wire_N_399[7]), 
            .I3(n16583), .O(n14_adj_4445));
    defparam i6_4_lut_adj_1438.LUT_INIT = 16'h0002;
    SB_LUT4 i2_2_lut (.I0(n42605), .I1(one_wire_N_399[10]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4446));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1439 (.I0(n7_adj_4446), .I1(one_wire_N_399[8]), 
            .I2(n42660), .I3(n14_adj_4445), .O(n49991));
    defparam i4_4_lut_adj_1439.LUT_INIT = 16'hfeff;
    SB_LUT4 i15704_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(16[20:25])
    defparam i15704_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 add_21_18_lut (.I0(n41781), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n34531), .O(n46644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_7_lut (.I0(n41781), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n34520), .O(n46633)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_18 (.CI(n34531), .I0(bit_ctr[16]), .I1(GND_net), .CO(n34532));
    SB_LUT4 i41883_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49784));
    defparam i41883_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n35633), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n35632), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n35632), .I0(n906), .I1(VCC_net), .CO(n35633));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n42682), .I2(VCC_net), 
            .I3(n35631), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n35631), .I0(n42682), .I1(VCC_net), 
            .CO(n35632));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17743), .I2(VCC_net), 
            .I3(n35630), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n35630), .I0(n17743), .I1(VCC_net), 
            .CO(n35631));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n15226), .I2(GND_net), 
            .I3(n35629), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n35629), .I0(n15226), .I1(GND_net), 
            .CO(n35630));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n35629));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4433), .I1(n4_adj_4433), .I2(n1037), 
            .I3(n35628), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n35627), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n35627), .I0(n1005), .I1(n1037), .CO(n35628));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n35626), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n35626), .I0(n1006), .I1(n1037), .CO(n35627));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n35625), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n35625), .I0(n1007), .I1(n1037), .CO(n35626));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n35624), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n35624), .I0(n1008), .I1(n1037), .CO(n35625));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n49786), 
            .I3(n35623), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n35623), .I0(n1009), .I1(n49786), .CO(n35624));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n49786), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n49786), 
            .CO(n35623));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n35622), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n35621), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n35621), .I0(n1104), .I1(n1136), .CO(n35622));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n35620), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n35620), .I0(n1105), .I1(n1136), .CO(n35621));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n35619), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n35619), .I0(n1106), .I1(n1136), .CO(n35620));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n35618), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n35618), .I0(n1107), .I1(n1136), .CO(n35619));
    SB_LUT4 add_21_17_lut (.I0(n41781), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n34530), .O(n46643)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n35617), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n35617), .I0(n1108), .I1(n1136), .CO(n35618));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n49787), 
            .I3(n35616), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n35616), .I0(n1109), .I1(n49787), .CO(n35617));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n49787), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n49787), 
            .CO(n35616));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n35615), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n35614), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n35614), .I0(n1203), .I1(n1235), .CO(n35615));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n35613), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n35613), .I0(n1204), .I1(n1235), .CO(n35614));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n35612), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n35612), .I0(n1205), .I1(n1235), .CO(n35613));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n35611), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_17 (.CI(n34530), .I0(bit_ctr[15]), .I1(GND_net), .CO(n34531));
    SB_CARRY mod_5_add_870_6 (.CI(n35611), .I0(n1206), .I1(n1235), .CO(n35612));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n35610), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n35610), .I0(n1207), .I1(n1235), .CO(n35611));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n35609), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n35609), .I0(n1208), .I1(n1235), .CO(n35610));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n49788), 
            .I3(n35608), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n35608), .I0(n1209), .I1(n49788), .CO(n35609));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n49788), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n49788), 
            .CO(n35608));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n35607), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n35606), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n35606), .I0(n1302), .I1(n1334), .CO(n35607));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n35605), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n35605), .I0(n1303), .I1(n1334), .CO(n35606));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n35604), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n35604), .I0(n1304), .I1(n1334), .CO(n35605));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n35603), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n35603), .I0(n1305), .I1(n1334), .CO(n35604));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n35602), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n35602), .I0(n1306), .I1(n1334), .CO(n35603));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n35601), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n35601), .I0(n1307), .I1(n1334), .CO(n35602));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n35600), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n35600), .I0(n1308), .I1(n1334), .CO(n35601));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n49789), 
            .I3(n35599), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i87_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n42));
    defparam i87_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62_4_lut (.I0(n94), .I1(n92_adj_4447), .I2(n42), .I3(one_wire_N_399[4]), 
            .O(n42563));   // verilog/neopixel.v(16[20:25])
    defparam i62_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i1_4_lut_adj_1440 (.I0(\state[1] ), .I1(start), .I2(n6_adj_4448), 
            .I3(n42563), .O(n35));   // verilog/neopixel.v(16[20:25])
    defparam i1_4_lut_adj_1440.LUT_INIT = 16'haaab;
    SB_CARRY mod_5_add_937_3 (.CI(n35599), .I0(n1309), .I1(n49789), .CO(n35600));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n49789), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n49789), 
            .CO(n35599));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n35598), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n35597), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n35597), .I0(n1401), .I1(n1433), .CO(n35598));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n35596), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n35596), .I0(n1402), .I1(n1433), .CO(n35597));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n35595), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n35595), .I0(n1403), .I1(n1433), .CO(n35596));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n35594), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n35594), .I0(n1404), .I1(n1433), .CO(n35595));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n35593), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n35593), .I0(n1405), .I1(n1433), .CO(n35594));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n35592), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n35592), .I0(n1406), .I1(n1433), .CO(n35593));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n35591), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n35591), .I0(n1407), .I1(n1433), .CO(n35592));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n35590), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n35590), .I0(n1408), .I1(n1433), .CO(n35591));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n49790), 
            .I3(n35589), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n35589), .I0(n1409), .I1(n49790), .CO(n35590));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n49790), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_7 (.CI(n34520), .I0(bit_ctr[5]), .I1(GND_net), .CO(n34521));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n49790), 
            .CO(n35589));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n35140), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n35139), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1441 (.I0(n2887), .I1(n2902), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4449));
    defparam i1_2_lut_adj_1441.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1442 (.I0(n2903), .I1(n2888), .I2(n2901), .I3(n2896), 
            .O(n42_adj_4450));
    defparam i17_4_lut_adj_1442.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2886), .I1(n2898), .I2(n2894), .I3(n2908), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1443 (.I0(n2905), .I1(n2890), .I2(n2904), .I3(n2889), 
            .O(n41));
    defparam i16_4_lut_adj_1443.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2891), .I1(n2892), .I2(n2906), .I3(n2899), 
            .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n2907), .I1(bit_ctr[6]), .I2(n2909), .I3(GND_net), 
            .O(n36_adj_4451));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i19_4_lut_adj_1444 (.I0(n2893), .I1(n2895), .I2(n2897), .I3(n26_adj_4449), 
            .O(n44));
    defparam i19_4_lut_adj_1444.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42_adj_4450), 
            .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_2_lut (.I0(n2885), .I1(n2900), .I2(GND_net), .I3(GND_net), 
            .O(n35_adj_4452));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n35_adj_4452), .I1(n48), .I2(n44), .I3(n36_adj_4451), 
            .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_23 (.CI(n35139), .I0(n2589), .I1(n2621), .CO(n35140));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n35138), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n35138), .I0(n2590), .I1(n2621), .CO(n35139));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n35137), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n35137), .I0(n2591), .I1(n2621), .CO(n35138));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n35136), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n35136), .I0(n2592), .I1(n2621), .CO(n35137));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n35135), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n35135), .I0(n2593), .I1(n2621), .CO(n35136));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n35134), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n35134), .I0(n2594), .I1(n2621), .CO(n35135));
    SB_LUT4 add_21_16_lut (.I0(n41781), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n34529), .O(n46642)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n35133), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n35133), .I0(n2595), .I1(n2621), .CO(n35134));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n35132), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n35132), .I0(n2596), .I1(n2621), .CO(n35133));
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n35131), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n35131), .I0(n2597), .I1(n2621), .CO(n35132));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n35130), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n35130), .I0(n2598), .I1(n2621), .CO(n35131));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n35129), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n35129), .I0(n2599), .I1(n2621), .CO(n35130));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n35128), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n35128), .I0(n2600), .I1(n2621), .CO(n35129));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n35127), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n35127), .I0(n2601), .I1(n2621), .CO(n35128));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n35126), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_10 (.CI(n35126), .I0(n2602), .I1(n2621), .CO(n35127));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n35125), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n35125), .I0(n2603), .I1(n2621), .CO(n35126));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n35124), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n35124), .I0(n2604), .I1(n2621), .CO(n35125));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n35123), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n35123), .I0(n2605), .I1(n2621), .CO(n35124));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n35542), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n35122), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n35122), .I0(n2606), .I1(n2621), .CO(n35123));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n35121), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n35121), .I0(n2607), .I1(n2621), .CO(n35122));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n35541), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n35541), .I0(n1500), .I1(n1532), .CO(n35542));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n35120), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n35540), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n35540), .I0(n1501), .I1(n1532), .CO(n35541));
    SB_CARRY mod_5_add_1808_4 (.CI(n35120), .I0(n2608), .I1(n2621), .CO(n35121));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n35539), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n35539), .I0(n1502), .I1(n1532), .CO(n35540));
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n49791), 
            .I3(n35119), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n35119), .I0(n2609), .I1(n49791), .CO(n35120));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n35538), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n49791), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_9 (.CI(n35538), .I0(n1503), .I1(n1532), .CO(n35539));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n49791), 
            .CO(n35119));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n35537), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n35537), .I0(n1504), .I1(n1532), .CO(n35538));
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n35536), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n35536), .I0(n1505), .I1(n1532), .CO(n35537));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n35535), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n35535), .I0(n1506), .I1(n1532), .CO(n35536));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n35534), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n35534), .I0(n1507), .I1(n1532), .CO(n35535));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n35533), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n35533), .I0(n1508), .I1(n1532), .CO(n35534));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n49792), 
            .I3(n35532), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1071_3 (.CI(n35532), .I0(n1509), .I1(n49792), .CO(n35533));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n49792), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n49792), 
            .CO(n35532));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n35531), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n35530), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n35530), .I0(n1599), .I1(n1631), .CO(n35531));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n35529), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n35529), .I0(n1600), .I1(n1631), .CO(n35530));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n35528), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n35528), .I0(n1601), .I1(n1631), .CO(n35529));
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n35527), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n35527), .I0(n1602), .I1(n1631), .CO(n35528));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n35526), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n35526), .I0(n1603), .I1(n1631), .CO(n35527));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n35525), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n35525), .I0(n1604), .I1(n1631), .CO(n35526));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n35524), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n35524), .I0(n1605), .I1(n1631), .CO(n35525));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n35523), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n35523), .I0(n1606), .I1(n1631), .CO(n35524));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n35522), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_adj_1445 (.I0(one_wire_N_399[4]), .I1(one_wire_N_399[2]), 
            .I2(one_wire_N_399[3]), .I3(GND_net), .O(n92_adj_4447));   // verilog/neopixel.v(53[15:25])
    defparam i2_3_lut_adj_1445.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(one_wire_N_399[7]), .I1(one_wire_N_399[10]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4453));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1447 (.I0(one_wire_N_399[8]), .I1(n16583), .I2(one_wire_N_399[11]), 
            .I3(n6_adj_4453), .O(n1));
    defparam i4_4_lut_adj_1447.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1448 (.I0(one_wire_N_399[9]), .I1(one_wire_N_399[5]), 
            .I2(one_wire_N_399[6]), .I3(GND_net), .O(n128));   // verilog/neopixel.v(53[15:25])
    defparam i2_3_lut_adj_1448.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1138_5 (.CI(n35522), .I0(n1607), .I1(n1631), .CO(n35523));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n35521), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(n121), .I1(one_wire_N_399[3]), .I2(GND_net), 
            .I3(GND_net), .O(n94));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1138_4 (.CI(n35521), .I0(n1608), .I1(n1631), .CO(n35522));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n49793), 
            .I3(n35520), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut_adj_1450 (.I0(n94), .I1(one_wire_N_399[4]), .I2(n128), 
            .I3(n1), .O(n29));
    defparam i3_4_lut_adj_1450.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1451 (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4455));
    defparam i2_2_lut_adj_1451.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48_adj_4456));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1452 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut_adj_1452.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1453 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut_adj_1453.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_3 (.CI(n35520), .I0(n1609), .I1(n49793), .CO(n35521));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n49793), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i16_4_lut_adj_1454 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44_adj_4457));
    defparam i16_4_lut_adj_1454.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1455 (.I0(bit_ctr[3]), .I1(n30_adj_4455), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut_adj_1455.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48_adj_4456), 
            .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44_adj_4457), 
            .O(\state_3__N_248[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1983_3_lut (.I0(n16572), .I1(\state_3__N_248[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4434));
    defparam i1983_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i41175_4_lut (.I0(n20911), .I1(n4434), .I2(\state[0] ), .I3(\state[1] ), 
            .O(n43079));
    defparam i41175_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i41882_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49783));
    defparam i41882_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n49793), 
            .CO(n35520));
    SB_LUT4 i15_4_lut_adj_1456 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_4458));
    defparam i15_4_lut_adj_1456.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1457 (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_4459));
    defparam i19_4_lut_adj_1457.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1458 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_4460));
    defparam i17_4_lut_adj_1458.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1459 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45_adj_4461));
    defparam i18_4_lut_adj_1459.LUT_INIT = 16'hfffe;
    SB_LUT4 i41880_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49781));
    defparam i41880_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1460 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_4462));
    defparam i16_4_lut_adj_1460.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), .I3(GND_net), 
            .O(n40_adj_4463));
    defparam i13_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i21_4_lut_adj_1461 (.I0(n3107), .I1(n42_adj_4458), .I2(n3087), 
            .I3(n3086), .O(n48_adj_4464));
    defparam i21_4_lut_adj_1461.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25_4_lut (.I0(n43_adj_4462), .I1(n45_adj_4461), .I2(n44_adj_4460), 
            .I3(n46_adj_4459), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3095), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n39_adj_4465));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut_adj_1462 (.I0(n39_adj_4465), .I1(n52), .I2(n48_adj_4464), 
            .I3(n40_adj_4463), .O(n3116));
    defparam i26_4_lut_adj_1462.LUT_INIT = 16'hfffe;
    SB_LUT4 i41881_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49782));
    defparam i41881_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n35510), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n35509), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n35509), .I0(n1698), .I1(n1730), .CO(n35510));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n35508), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n35508), .I0(n1699), .I1(n1730), .CO(n35509));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n35507), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4466));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1463 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4467));
    defparam i1_3_lut_adj_1463.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1464 (.I0(n2490), .I1(n34), .I2(n24_adj_4466), 
            .I3(n2494), .O(n38));
    defparam i17_4_lut_adj_1464.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1465 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4468));
    defparam i15_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1466 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4467), 
            .O(n37_adj_4469));
    defparam i16_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1467 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4470));
    defparam i14_4_lut_adj_1467.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1468 (.I0(n35_adj_4470), .I1(n37_adj_4469), .I2(n36_adj_4468), 
            .I3(n38), .O(n2522));
    defparam i20_4_lut_adj_1468.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_12 (.CI(n35507), .I0(n1700), .I1(n1730), .CO(n35508));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n35506), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n35506), .I0(n1701), .I1(n1730), .CO(n35507));
    SB_LUT4 add_21_6_lut (.I0(n41781), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n34519), .O(n46632)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n35505), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n35505), .I0(n1702), .I1(n1730), .CO(n35506));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n35504), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n35504), .I0(n1703), .I1(n1730), .CO(n35505));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n35503), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n35503), .I0(n1704), .I1(n1730), .CO(n35504));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n35502), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n35502), .I0(n1705), .I1(n1730), .CO(n35503));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n35501), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n35501), .I0(n1706), .I1(n1730), .CO(n35502));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n35500), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n35500), .I0(n1707), .I1(n1730), .CO(n35501));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n35499), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n35499), .I0(n1708), .I1(n1730), .CO(n35500));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n49794), 
            .I3(n35498), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n35498), .I0(n1709), .I1(n49794), .CO(n35499));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n49794), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n49794), 
            .CO(n35498));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n35483), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n35482), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n35482), .I0(n1797), .I1(n1829), .CO(n35483));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n35481), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n35481), .I0(n1798), .I1(n1829), .CO(n35482));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n35480), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n35480), .I0(n1799), .I1(n1829), .CO(n35481));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n35479), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n35479), .I0(n1800), .I1(n1829), .CO(n35480));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n35478), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n35478), .I0(n1801), .I1(n1829), .CO(n35479));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n35477), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n35477), .I0(n1802), .I1(n1829), .CO(n35478));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n35476), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n35476), .I0(n1803), .I1(n1829), .CO(n35477));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n35475), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n35475), .I0(n1804), .I1(n1829), .CO(n35476));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n35474), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n35474), .I0(n1805), .I1(n1829), .CO(n35475));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n35473), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n35473), .I0(n1806), .I1(n1829), .CO(n35474));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n35472), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n35472), .I0(n1807), .I1(n1829), .CO(n35473));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n35471), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n35471), .I0(n1808), .I1(n1829), .CO(n35472));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n49795), 
            .I3(n35470), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n35470), .I0(n1809), .I1(n49795), .CO(n35471));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n49795), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n49795), 
            .CO(n35470));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n35469), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n35468), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n35468), .I0(n1896), .I1(n1928), .CO(n35469));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n35467), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n35467), .I0(n1897), .I1(n1928), .CO(n35468));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n35466), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n35466), .I0(n1898), .I1(n1928), .CO(n35467));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n35079), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n35465), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n35465), .I0(n1899), .I1(n1928), .CO(n35466));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n35078), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n35464), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n35464), .I0(n1900), .I1(n1928), .CO(n35465));
    SB_CARRY mod_5_add_1875_24 (.CI(n35078), .I0(n2688), .I1(n2720), .CO(n35079));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n35463), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n35463), .I0(n1901), .I1(n1928), .CO(n35464));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n35077), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n35462), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n35462), .I0(n1902), .I1(n1928), .CO(n35463));
    SB_CARRY mod_5_add_1875_23 (.CI(n35077), .I0(n2689), .I1(n2720), .CO(n35078));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n35461), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n35461), .I0(n1903), .I1(n1928), .CO(n35462));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n35076), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n35460), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n35460), .I0(n1904), .I1(n1928), .CO(n35461));
    SB_CARRY mod_5_add_1875_22 (.CI(n35076), .I0(n2690), .I1(n2720), .CO(n35077));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n35459), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n35459), .I0(n1905), .I1(n1928), .CO(n35460));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n35075), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n35458), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n35458), .I0(n1906), .I1(n1928), .CO(n35459));
    SB_CARRY mod_5_add_1875_21 (.CI(n35075), .I0(n2691), .I1(n2720), .CO(n35076));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n35457), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n35457), .I0(n1907), .I1(n1928), .CO(n35458));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n35074), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n35456), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n35456), .I0(n1908), .I1(n1928), .CO(n35457));
    SB_CARRY mod_5_add_1875_20 (.CI(n35074), .I0(n2692), .I1(n2720), .CO(n35075));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n49796), 
            .I3(n35455), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n35455), .I0(n1909), .I1(n49796), .CO(n35456));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n35073), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n49796), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n49796), 
            .CO(n35455));
    SB_CARRY mod_5_add_1875_19 (.CI(n35073), .I0(n2693), .I1(n2720), .CO(n35074));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n35454), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n35453), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n35072), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n35453), .I0(n1995), .I1(n2027), .CO(n35454));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n35452), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n35072), .I0(n2694), .I1(n2720), .CO(n35073));
    SB_CARRY mod_5_add_1406_16 (.CI(n35452), .I0(n1996), .I1(n2027), .CO(n35453));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n35451), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n35071), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n35451), .I0(n1997), .I1(n2027), .CO(n35452));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n35450), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n35071), .I0(n2695), .I1(n2720), .CO(n35072));
    SB_CARRY mod_5_add_1406_14 (.CI(n35450), .I0(n1998), .I1(n2027), .CO(n35451));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n35449), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n35070), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n35449), .I0(n1999), .I1(n2027), .CO(n35450));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n35448), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n35448), .I0(n2000), .I1(n2027), .CO(n35449));
    SB_CARRY mod_5_add_1875_16 (.CI(n35070), .I0(n2696), .I1(n2720), .CO(n35071));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n35069), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n35447), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n35447), .I0(n2001), .I1(n2027), .CO(n35448));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n35446), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n35069), .I0(n2697), .I1(n2720), .CO(n35070));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n35068), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n35446), .I0(n2002), .I1(n2027), .CO(n35447));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n35445), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n35068), .I0(n2698), .I1(n2720), .CO(n35069));
    SB_CARRY mod_5_add_1406_9 (.CI(n35445), .I0(n2003), .I1(n2027), .CO(n35446));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n35444), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n35067), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n35444), .I0(n2004), .I1(n2027), .CO(n35445));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n35443), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n35067), .I0(n2699), .I1(n2720), .CO(n35068));
    SB_CARRY mod_5_add_1406_7 (.CI(n35443), .I0(n2005), .I1(n2027), .CO(n35444));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n35442), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n35066), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n35442), .I0(n2006), .I1(n2027), .CO(n35443));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n35441), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n35066), .I0(n2700), .I1(n2720), .CO(n35067));
    SB_CARRY mod_5_add_1406_5 (.CI(n35441), .I0(n2007), .I1(n2027), .CO(n35442));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n35440), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n35065), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n35440), .I0(n2008), .I1(n2027), .CO(n35441));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n49798), 
            .I3(n35439), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_11 (.CI(n35065), .I0(n2701), .I1(n2720), .CO(n35066));
    SB_CARRY mod_5_add_1406_3 (.CI(n35439), .I0(n2009), .I1(n49798), .CO(n35440));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n49798), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n35064), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n49798), 
            .CO(n35439));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n35438), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n35064), .I0(n2702), .I1(n2720), .CO(n35065));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n35437), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n35437), .I0(n2094), .I1(n2126), .CO(n35438));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n35436), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n35063), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n35436), .I0(n2095), .I1(n2126), .CO(n35437));
    SB_CARRY mod_5_add_1875_9 (.CI(n35063), .I0(n2703), .I1(n2720), .CO(n35064));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n35062), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n35435), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n35062), .I0(n2704), .I1(n2720), .CO(n35063));
    SB_CARRY mod_5_add_1473_16 (.CI(n35435), .I0(n2096), .I1(n2126), .CO(n35436));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n35434), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n35434), .I0(n2097), .I1(n2126), .CO(n35435));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n35433), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n35061), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n35061), .I0(n2705), .I1(n2720), .CO(n35062));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n35060), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n35060), .I0(n2706), .I1(n2720), .CO(n35061));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n35059), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n35433), .I0(n2098), .I1(n2126), .CO(n35434));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n35432), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n35432), .I0(n2099), .I1(n2126), .CO(n35433));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n35431), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n35059), .I0(n2707), .I1(n2720), .CO(n35060));
    SB_CARRY mod_5_add_1473_12 (.CI(n35431), .I0(n2100), .I1(n2126), .CO(n35432));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n35058), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n35430), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n34529), .I0(bit_ctr[14]), .I1(GND_net), .CO(n34530));
    SB_CARRY mod_5_add_1875_4 (.CI(n35058), .I0(n2708), .I1(n2720), .CO(n35059));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n49797), 
            .I3(n35057), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_11 (.CI(n35430), .I0(n2101), .I1(n2126), .CO(n35431));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n35429), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n34519), .I0(bit_ctr[4]), .I1(GND_net), .CO(n34520));
    SB_CARRY mod_5_add_1473_10 (.CI(n35429), .I0(n2102), .I1(n2126), .CO(n35430));
    SB_LUT4 add_21_15_lut (.I0(n41781), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n34528), .O(n46641)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n35428), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_3 (.CI(n35057), .I0(n2709), .I1(n49797), .CO(n35058));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n49797), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n49797), 
            .CO(n35057));
    SB_CARRY mod_5_add_1473_9 (.CI(n35428), .I0(n2103), .I1(n2126), .CO(n35429));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n35427), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n35427), .I0(n2104), .I1(n2126), .CO(n35428));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n35426), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n35426), .I0(n2105), .I1(n2126), .CO(n35427));
    SB_LUT4 add_21_5_lut (.I0(n41781), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n34518), .O(n46631)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n35425), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n35425), .I0(n2106), .I1(n2126), .CO(n35426));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n35424), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n35424), .I0(n2107), .I1(n2126), .CO(n35425));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n35423), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n35423), .I0(n2108), .I1(n2126), .CO(n35424));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n49799), 
            .I3(n35422), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n35422), .I0(n2109), .I1(n49799), .CO(n35423));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n49799), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n49799), 
            .CO(n35422));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n35421), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n35420), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n35420), .I0(n2193), .I1(n2225), .CO(n35421));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n35419), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n35419), .I0(n2194), .I1(n2225), .CO(n35420));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n35418), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n35418), .I0(n2195), .I1(n2225), .CO(n35419));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n35417), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n35417), .I0(n2196), .I1(n2225), .CO(n35418));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n35416), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n35416), .I0(n2197), .I1(n2225), .CO(n35417));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n35415), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_15 (.CI(n34528), .I0(bit_ctr[13]), .I1(GND_net), .CO(n34529));
    SB_CARRY mod_5_add_1540_14 (.CI(n35415), .I0(n2198), .I1(n2225), .CO(n35416));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n35414), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n35414), .I0(n2199), .I1(n2225), .CO(n35415));
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n35413), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1189__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_DFF timer_1189__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY add_21_5 (.CI(n34518), .I0(bit_ctr[3]), .I1(GND_net), .CO(n34519));
    SB_CARRY mod_5_add_1540_12 (.CI(n35413), .I0(n2200), .I1(n2225), .CO(n35414));
    SB_LUT4 add_21_14_lut (.I0(n41781), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n34527), .O(n46640)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n35412), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n35412), .I0(n2201), .I1(n2225), .CO(n35413));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n35411), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n35411), .I0(n2202), .I1(n2225), .CO(n35412));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n35410), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n35410), .I0(n2203), .I1(n2225), .CO(n35411));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n35409), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n34527), .I0(bit_ctr[12]), .I1(GND_net), .CO(n34528));
    SB_CARRY mod_5_add_1540_8 (.CI(n35409), .I0(n2204), .I1(n2225), .CO(n35410));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n35408), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n35408), .I0(n2205), .I1(n2225), .CO(n35409));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n35407), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n35407), .I0(n2206), .I1(n2225), .CO(n35408));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n35406), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n35406), .I0(n2207), .I1(n2225), .CO(n35407));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n35405), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n35405), .I0(n2208), .I1(n2225), .CO(n35406));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n49800), 
            .I3(n35404), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n35404), .I0(n2209), .I1(n49800), .CO(n35405));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n49800), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n49800), 
            .CO(n35404));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n35403), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n35402), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n35402), .I0(n2292), .I1(n2324), .CO(n35403));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n35401), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n35401), .I0(n2293), .I1(n2324), .CO(n35402));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n35400), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n35400), .I0(n2294), .I1(n2324), .CO(n35401));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n35399), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n35399), .I0(n2295), .I1(n2324), .CO(n35400));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n35026), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(n41781), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n34526), .O(n46639)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n35025), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n35398), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n35025), .I0(n2787), .I1(n2819), .CO(n35026));
    SB_CARRY mod_5_add_1607_16 (.CI(n35398), .I0(n2296), .I1(n2324), .CO(n35399));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n35024), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_4_lut (.I0(n41781), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n34517), .O(n46630)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n35397), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n35397), .I0(n2297), .I1(n2324), .CO(n35398));
    SB_CARRY mod_5_add_1942_24 (.CI(n35024), .I0(n2788), .I1(n2819), .CO(n35025));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n35023), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n35023), .I0(n2789), .I1(n2819), .CO(n35024));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n35396), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n35396), .I0(n2298), .I1(n2324), .CO(n35397));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n35022), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_4 (.CI(n34517), .I0(bit_ctr[2]), .I1(GND_net), .CO(n34518));
    SB_CARRY mod_5_add_1942_22 (.CI(n35022), .I0(n2790), .I1(n2819), .CO(n35023));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n35395), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1189__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1189__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n35021), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n35021), .I0(n2791), .I1(n2819), .CO(n35022));
    SB_CARRY mod_5_add_1607_13 (.CI(n35395), .I0(n2299), .I1(n2324), .CO(n35396));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n35020), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n35394), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n35020), .I0(n2792), .I1(n2819), .CO(n35021));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n35019), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n35019), .I0(n2793), .I1(n2819), .CO(n35020));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n35018), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n35394), .I0(n2300), .I1(n2324), .CO(n35395));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n35393), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n35018), .I0(n2794), .I1(n2819), .CO(n35019));
    SB_CARRY mod_5_add_1607_11 (.CI(n35393), .I0(n2301), .I1(n2324), .CO(n35394));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n35392), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n35017), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n35392), .I0(n2302), .I1(n2324), .CO(n35393));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n35391), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n35017), .I0(n2795), .I1(n2819), .CO(n35018));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n35016), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n35391), .I0(n2303), .I1(n2324), .CO(n35392));
    SB_CARRY mod_5_add_1942_16 (.CI(n35016), .I0(n2796), .I1(n2819), .CO(n35017));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n35015), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n35390), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n35390), .I0(n2304), .I1(n2324), .CO(n35391));
    SB_CARRY mod_5_add_1942_15 (.CI(n35015), .I0(n2797), .I1(n2819), .CO(n35016));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n35389), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n35389), .I0(n2305), .I1(n2324), .CO(n35390));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n35014), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n35014), .I0(n2798), .I1(n2819), .CO(n35015));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n35388), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n35388), .I0(n2306), .I1(n2324), .CO(n35389));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n35013), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n35387), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n35013), .I0(n2799), .I1(n2819), .CO(n35014));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n35012), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n35387), .I0(n2307), .I1(n2324), .CO(n35388));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n35386), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n35386), .I0(n2308), .I1(n2324), .CO(n35387));
    SB_CARRY mod_5_add_1942_12 (.CI(n35012), .I0(n2800), .I1(n2819), .CO(n35013));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n49801), 
            .I3(n35385), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n35011), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_3 (.CI(n35385), .I0(n2309), .I1(n49801), .CO(n35386));
    SB_CARRY mod_5_add_1942_11 (.CI(n35011), .I0(n2801), .I1(n2819), .CO(n35012));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n49801), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n35010), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n49801), 
            .CO(n35385));
    SB_CARRY mod_5_add_1942_10 (.CI(n35010), .I0(n2802), .I1(n2819), .CO(n35011));
    SB_LUT4 timer_1189_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n35384), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1189_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n35383), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n35009), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n35009), .I0(n2803), .I1(n2819), .CO(n35010));
    SB_CARRY timer_1189_add_4_32 (.CI(n35383), .I0(GND_net), .I1(timer[30]), 
            .CO(n35384));
    SB_LUT4 timer_1189_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n35382), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n35008), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n35008), .I0(n2804), .I1(n2819), .CO(n35009));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n35007), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1189_add_4_31 (.CI(n35382), .I0(GND_net), .I1(timer[29]), 
            .CO(n35383));
    SB_LUT4 timer_1189_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n35381), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_30 (.CI(n35381), .I0(GND_net), .I1(timer[28]), 
            .CO(n35382));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17665), .D(state_3__N_248[0]), 
            .S(n17802));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_3_lut (.I0(n41781), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n34516), .O(n46629)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1189_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n35380), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_7 (.CI(n35007), .I0(n2805), .I1(n2819), .CO(n35008));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n35006), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1189_add_4_29 (.CI(n35380), .I0(GND_net), .I1(timer[27]), 
            .CO(n35381));
    SB_LUT4 timer_1189_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n35379), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n35006), .I0(n2806), .I1(n2819), .CO(n35007));
    SB_CARRY timer_1189_add_4_28 (.CI(n35379), .I0(GND_net), .I1(timer[26]), 
            .CO(n35380));
    SB_LUT4 timer_1189_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n35378), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_27 (.CI(n35378), .I0(GND_net), .I1(timer[25]), 
            .CO(n35379));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n35005), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_33_lut (.I0(n41781), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n34546), .O(n46659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_5 (.CI(n35005), .I0(n2807), .I1(n2819), .CO(n35006));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n35004), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1189_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n35377), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n34526), .I0(bit_ctr[11]), .I1(GND_net), .CO(n34527));
    SB_CARRY timer_1189_add_4_26 (.CI(n35377), .I0(GND_net), .I1(timer[24]), 
            .CO(n35378));
    SB_LUT4 add_21_32_lut (.I0(n41781), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n34545), .O(n46658)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1189_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n35376), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_4 (.CI(n35004), .I0(n2808), .I1(n2819), .CO(n35005));
    SB_CARRY timer_1189_add_4_25 (.CI(n35376), .I0(GND_net), .I1(timer[23]), 
            .CO(n35377));
    SB_LUT4 timer_1189_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n35375), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n49802), 
            .I3(n35003), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1189_add_4_24 (.CI(n35375), .I0(GND_net), .I1(timer[22]), 
            .CO(n35376));
    SB_CARRY mod_5_add_1942_3 (.CI(n35003), .I0(n2809), .I1(n49802), .CO(n35004));
    SB_LUT4 timer_1189_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n35374), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n49802), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1189_add_4_23 (.CI(n35374), .I0(GND_net), .I1(timer[21]), 
            .CO(n35375));
    SB_LUT4 add_21_12_lut (.I0(n41781), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n34525), .O(n46638)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n49802), 
            .CO(n35003));
    SB_CARRY add_21_12 (.CI(n34525), .I0(bit_ctr[10]), .I1(GND_net), .CO(n34526));
    SB_LUT4 timer_1189_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n35373), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_22 (.CI(n35373), .I0(GND_net), .I1(timer[20]), 
            .CO(n35374));
    SB_CARRY add_21_32 (.CI(n34545), .I0(bit_ctr[30]), .I1(GND_net), .CO(n34546));
    SB_LUT4 timer_1189_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n35372), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_31_lut (.I0(n41781), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n34544), .O(n46657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1189_add_4_21 (.CI(n35372), .I0(GND_net), .I1(timer[19]), 
            .CO(n35373));
    SB_LUT4 timer_1189_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n35371), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_20 (.CI(n35371), .I0(GND_net), .I1(timer[18]), 
            .CO(n35372));
    SB_LUT4 timer_1189_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n35370), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_19 (.CI(n35370), .I0(GND_net), .I1(timer[17]), 
            .CO(n35371));
    SB_CARRY add_21_31 (.CI(n34544), .I0(bit_ctr[29]), .I1(GND_net), .CO(n34545));
    SB_LUT4 timer_1189_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n35369), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_30_lut (.I0(n41781), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n34543), .O(n46656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1189_add_4_18 (.CI(n35369), .I0(GND_net), .I1(timer[16]), 
            .CO(n35370));
    SB_CARRY add_21_30 (.CI(n34543), .I0(bit_ctr[28]), .I1(GND_net), .CO(n34544));
    SB_LUT4 timer_1189_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n35368), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_17 (.CI(n35368), .I0(GND_net), .I1(timer[15]), 
            .CO(n35369));
    SB_LUT4 timer_1189_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n35367), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_29_lut (.I0(n41781), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n34542), .O(n46655)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1189_add_4_16 (.CI(n35367), .I0(GND_net), .I1(timer[14]), 
            .CO(n35368));
    SB_LUT4 timer_1189_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n35366), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_15 (.CI(n35366), .I0(GND_net), .I1(timer[13]), 
            .CO(n35367));
    SB_LUT4 timer_1189_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n35365), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_14 (.CI(n35365), .I0(GND_net), .I1(timer[12]), 
            .CO(n35366));
    SB_LUT4 timer_1189_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n35364), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_13 (.CI(n35364), .I0(GND_net), .I1(timer[11]), 
            .CO(n35365));
    SB_LUT4 timer_1189_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n35363), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n34542), .I0(bit_ctr[27]), .I1(GND_net), .CO(n34543));
    SB_CARRY timer_1189_add_4_12 (.CI(n35363), .I0(GND_net), .I1(timer[10]), 
            .CO(n35364));
    SB_LUT4 timer_1189_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n35362), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_11 (.CI(n35362), .I0(GND_net), .I1(timer[9]), 
            .CO(n35363));
    SB_LUT4 timer_1189_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n35361), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_28_lut (.I0(n41781), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n34541), .O(n46654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1189_add_4_10 (.CI(n35361), .I0(GND_net), .I1(timer[8]), 
            .CO(n35362));
    SB_LUT4 timer_1189_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n35360), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_9 (.CI(n35360), .I0(GND_net), .I1(timer[7]), 
            .CO(n35361));
    SB_LUT4 timer_1189_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n35359), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_8 (.CI(n35359), .I0(GND_net), .I1(timer[6]), 
            .CO(n35360));
    SB_LUT4 timer_1189_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n35358), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_7 (.CI(n35358), .I0(GND_net), .I1(timer[5]), 
            .CO(n35359));
    SB_LUT4 add_21_11_lut (.I0(n41781), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n34524), .O(n46637)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_28 (.CI(n34541), .I0(bit_ctr[26]), .I1(GND_net), .CO(n34542));
    SB_LUT4 timer_1189_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n35357), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_6 (.CI(n35357), .I0(GND_net), .I1(timer[4]), 
            .CO(n35358));
    SB_LUT4 timer_1189_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n35356), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_27_lut (.I0(n41781), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n34540), .O(n46653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1189_add_4_5 (.CI(n35356), .I0(GND_net), .I1(timer[3]), 
            .CO(n35357));
    SB_LUT4 timer_1189_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n35355), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n34516), .I0(bit_ctr[1]), .I1(GND_net), .CO(n34517));
    SB_CARRY add_21_27 (.CI(n34540), .I0(bit_ctr[25]), .I1(GND_net), .CO(n34541));
    SB_CARRY timer_1189_add_4_4 (.CI(n35355), .I0(GND_net), .I1(timer[2]), 
            .CO(n35356));
    SB_LUT4 timer_1189_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n35354), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_3 (.CI(n35354), .I0(GND_net), .I1(timer[1]), 
            .CO(n35355));
    SB_LUT4 timer_1189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n35354));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n35353), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n35352), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n35352), .I0(n2391), .I1(n2423), .CO(n35353));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n35351), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n35351), .I0(n2392), .I1(n2423), .CO(n35352));
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17984));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n35350), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n35350), .I0(n2393), .I1(n2423), .CO(n35351));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n35349), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n35349), .I0(n2394), .I1(n2423), .CO(n35350));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n35348), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n35348), .I0(n2395), .I1(n2423), .CO(n35349));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n35347), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n35347), .I0(n2396), .I1(n2423), .CO(n35348));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n35346), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n35346), .I0(n2397), .I1(n2423), .CO(n35347));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n35345), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n35345), .I0(n2398), .I1(n2423), .CO(n35346));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n35344), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n35344), .I0(n2399), .I1(n2423), .CO(n35345));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n35343), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n35343), .I0(n2400), .I1(n2423), .CO(n35344));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n35342), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n35342), .I0(n2401), .I1(n2423), .CO(n35343));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n35341), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n35341), .I0(n2402), .I1(n2423), .CO(n35342));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n35340), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n35340), .I0(n2403), .I1(n2423), .CO(n35341));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n35339), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n35339), .I0(n2404), .I1(n2423), .CO(n35340));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n35338), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n35338), .I0(n2405), .I1(n2423), .CO(n35339));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n35337), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_26_lut (.I0(n41781), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n34539), .O(n46652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_11 (.CI(n34524), .I0(bit_ctr[9]), .I1(GND_net), .CO(n34525));
    SB_CARRY add_21_26 (.CI(n34539), .I0(bit_ctr[24]), .I1(GND_net), .CO(n34540));
    SB_CARRY mod_5_add_1674_6 (.CI(n35337), .I0(n2406), .I1(n2423), .CO(n35338));
    SB_LUT4 add_21_25_lut (.I0(n41781), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n34538), .O(n46651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n35336), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n35336), .I0(n2407), .I1(n2423), .CO(n35337));
    SB_CARRY add_21_25 (.CI(n34538), .I0(bit_ctr[23]), .I1(GND_net), .CO(n34539));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n35335), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(n41781), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n34523), .O(n46636)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_4 (.CI(n35335), .I0(n2408), .I1(n2423), .CO(n35336));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n49803), 
            .I3(n35334), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n35334), .I0(n2409), .I1(n49803), .CO(n35335));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n49803), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n49803), 
            .CO(n35334));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n34987), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(n41781), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n34537), .O(n46650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_2_lut (.I0(n41781), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n46628)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_DFFESR one_wire_108 (.Q(PIN_14_c), .C(clk32MHz), .E(n17611), .D(\neo_pixel_transmitter.done_N_462 ), 
            .R(n44172));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_10 (.CI(n34523), .I0(bit_ctr[8]), .I1(GND_net), .CO(n34524));
    SB_CARRY add_21_24 (.CI(n34537), .I0(bit_ctr[22]), .I1(GND_net), .CO(n34538));
    SB_LUT4 add_21_23_lut (.I0(n41781), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n34536), .O(n46649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n34986), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n34986), .I0(n2886), .I1(n2918), .CO(n34987));
    SB_LUT4 add_21_9_lut (.I0(n41781), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n34522), .O(n46635)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n34985), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n34985), .I0(n2887), .I1(n2918), .CO(n34986));
    SB_CARRY add_21_23 (.CI(n34536), .I0(bit_ctr[21]), .I1(GND_net), .CO(n34537));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n34516));
    SB_CARRY add_21_9 (.CI(n34522), .I0(bit_ctr[7]), .I1(GND_net), .CO(n34523));
    SB_LUT4 add_21_22_lut (.I0(n41781), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n34535), .O(n46648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n34984), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_22 (.CI(n34535), .I0(bit_ctr[20]), .I1(GND_net), .CO(n34536));
    SB_LUT4 add_21_21_lut (.I0(n41781), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n34534), .O(n46647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2009_24 (.CI(n34984), .I0(n2888), .I1(n2918), .CO(n34985));
    SB_CARRY add_21_21 (.CI(n34534), .I0(bit_ctr[19]), .I1(GND_net), .CO(n34535));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n34983), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n34983), .I0(n2889), .I1(n2918), .CO(n34984));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n34982), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n34982), .I0(n2890), .I1(n2918), .CO(n34983));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n34981), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n34981), .I0(n2891), .I1(n2918), .CO(n34982));
    SB_LUT4 i1_2_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n29), .I3(GND_net), .O(n16572));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_adj_1469 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n17574), .I3(GND_net), .O(n20911));
    defparam i1_2_lut_3_lut_adj_1469.LUT_INIT = 16'hbfbf;
    SB_LUT4 i223_2_lut (.I0(n26050), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n852));   // verilog/neopixel.v(103[9] 111[12])
    defparam i223_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15680_3_lut (.I0(n20911), .I1(n41777), .I2(\state[0] ), .I3(GND_net), 
            .O(n20959));   // verilog/neopixel.v(16[20:25])
    defparam i15680_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_4_lut_adj_1470 (.I0(\state[0] ), .I1(n20959), .I2(n852), 
            .I3(\state[1] ), .O(n17665));
    defparam i1_4_lut_adj_1470.LUT_INIT = 16'hafcc;
    SB_LUT4 i25_4_lut_adj_1471 (.I0(n20911), .I1(n26050), .I2(\state[1] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n11_adj_4471));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_4_lut_adj_1471.LUT_INIT = 16'h05c5;
    SB_LUT4 i24_4_lut_adj_1472 (.I0(n11_adj_4471), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(n41777), .O(n17802));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_4_lut_adj_1472.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14_4_lut_adj_1473 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4472));
    defparam i14_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1474 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4473));
    defparam i18_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1475 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4474));
    defparam i16_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1476 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4475));
    defparam i17_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1477 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4476));
    defparam i15_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1478 (.I0(n3001), .I1(n2993), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4477));
    defparam i12_2_lut_adj_1478.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4472), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4478));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(\color[2] ), .I2(\color[3] ), 
            .I3(bit_ctr[1]), .O(n49907));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i24_4_lut_adj_1479 (.I0(n41_adj_4476), .I1(n43_adj_4475), .I2(n42_adj_4474), 
            .I3(n44_adj_4473), .O(n50));
    defparam i24_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut_adj_1480 (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), 
            .I3(GND_net), .O(n37_adj_4479));
    defparam i11_3_lut_adj_1480.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut_adj_1481 (.I0(n37_adj_4479), .I1(n50), .I2(n46_adj_4478), 
            .I3(n38_adj_4477), .O(n3017));
    defparam i25_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i29121_2_lut (.I0(bit_ctr[3]), .I1(n26090), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_442[3]));   // verilog/neopixel.v(22[26:36])
    defparam i29121_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34676_2_lut (.I0(one_wire_N_399[2]), .I1(one_wire_N_399[4]), 
            .I2(GND_net), .I3(GND_net), .O(n42557));
    defparam i34676_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1482 (.I0(\state[1] ), .I1(n26050), .I2(GND_net), 
            .I3(GND_net), .O(n41814));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1482.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1483 (.I0(one_wire_N_399[3]), .I1(n42557), .I2(n42), 
            .I3(n92), .O(n60_adj_4480));
    defparam i1_4_lut_adj_1483.LUT_INIT = 16'h7350;
    SB_LUT4 i80_4_lut (.I0(n41814), .I1(n42557), .I2(\neo_pixel_transmitter.done ), 
            .I3(n4_adj_4481), .O(n54_adj_4482));
    defparam i80_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i1_4_lut_adj_1484 (.I0(n29), .I1(n116), .I2(n42), .I3(n60_adj_4480), 
            .O(n57));
    defparam i1_4_lut_adj_1484.LUT_INIT = 16'h3705;
    SB_LUT4 i1_4_lut_adj_1485 (.I0(\state[0] ), .I1(n57), .I2(n54_adj_4482), 
            .I3(n42605), .O(n17611));
    defparam i1_4_lut_adj_1485.LUT_INIT = 16'h50dc;
    SB_LUT4 i50_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_462 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i50_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20785_4_lut (.I0(one_wire_N_399[9]), .I1(n16583), .I2(one_wire_N_399[11]), 
            .I3(one_wire_N_399[10]), .O(n26050));
    defparam i20785_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_adj_1487 (.I0(n26050), .I1(\state[0] ), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n43650));   // verilog/neopixel.v(36[4] 116[11])
    defparam i2_3_lut_adj_1487.LUT_INIT = 16'hfdfd;
    SB_LUT4 i41902_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49803));
    defparam i41902_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2395), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_4484));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1488 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4485));
    defparam i13_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2392), .I1(n2399), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4486));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2407), .I1(n2402), .I2(n2408), .I3(n2396), 
            .O(n31_adj_4487));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1489 (.I0(n2393), .I1(n2406), .I2(n2405), .I3(n2403), 
            .O(n35_adj_4488));
    defparam i15_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1490 (.I0(n33_adj_4485), .I1(n27_adj_4484), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4489));
    defparam i17_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1491 (.I0(n37_adj_4489), .I1(n35_adj_4488), .I2(n31_adj_4487), 
            .I3(n32_adj_4486), .O(n2423));
    defparam i19_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 n49907_bdd_4_lut (.I0(n49907), .I1(\color[1] ), .I2(\color[0] ), 
            .I3(bit_ctr[1]), .O(n44398));
    defparam n49907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i41901_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49802));
    defparam i41901_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20734_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n25994));
    defparam i20734_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1492 (.I0(n3196), .I1(n3208), .I2(n3199), .I3(n3188), 
            .O(n48_adj_4490));
    defparam i20_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1493 (.I0(n3195), .I1(n3202), .I2(n3187), .I3(n3194), 
            .O(n46_adj_4491));
    defparam i18_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1494 (.I0(n3200), .I1(n3185), .I2(n3182), .I3(n3192), 
            .O(n47_adj_4492));
    defparam i19_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1495 (.I0(n3201), .I1(n3197), .I2(n3190), .I3(n3183), 
            .O(n45_adj_4493));
    defparam i17_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1496 (.I0(n3184), .I1(n3205), .I2(n3206), .I3(n3186), 
            .O(n44_adj_4494));
    defparam i16_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1497 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n25994), 
            .O(n43_adj_4495));
    defparam i15_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1498 (.I0(n45_adj_4493), .I1(n47_adj_4492), .I2(n46_adj_4491), 
            .I3(n48_adj_4490), .O(n54_adj_4496));
    defparam i26_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1499 (.I0(n3191), .I1(n3207), .I2(n3204), .I3(n3203), 
            .O(n49_adj_4497));
    defparam i21_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1500 (.I0(n49_adj_4497), .I1(n54_adj_4496), .I2(n43_adj_4495), 
            .I3(n44_adj_4494), .O(n26090));
    defparam i27_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i39442_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n26090), .I3(GND_net), 
            .O(color_bit_N_442[4]));
    defparam i39442_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i40039_4_lut (.I0(n49868), .I1(bit_ctr[2]), .I2(bit_ctr[3]), 
            .I3(n26090), .O(n46586));
    defparam i40039_4_lut.LUT_INIT = 16'h2002;
    SB_LUT4 i20055_4_lut (.I0(n49808), .I1(\state_3__N_248[1] ), .I2(n46586), 
            .I3(color_bit_N_442[4]), .O(state_3__N_248[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i20055_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i41900_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49801));
    defparam i41900_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1501 (.I0(n2803), .I1(n2792), .I2(n2807), .I3(n2801), 
            .O(n40_adj_4498));
    defparam i16_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1502 (.I0(n2808), .I1(n2798), .I2(n2788), .I3(n2796), 
            .O(n38_adj_4499));
    defparam i14_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1503 (.I0(n2794), .I1(n2789), .I2(n2805), .I3(n2797), 
            .O(n39_adj_4500));
    defparam i15_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1504 (.I0(n2804), .I1(n2793), .I2(n2795), .I3(n2802), 
            .O(n37_adj_4501));
    defparam i13_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut_adj_1505 (.I0(n2787), .I1(n2800), .I2(GND_net), 
            .I3(GND_net), .O(n34_adj_4502));
    defparam i10_2_lut_adj_1505.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1506 (.I0(n2791), .I1(n2790), .I2(n2799), .I3(n2806), 
            .O(n42_adj_4503));
    defparam i18_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n37_adj_4501), .I1(n39_adj_4500), .I2(n38_adj_4499), 
            .I3(n40_adj_4498), .O(n46_adj_4504));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2786), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4505));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1507 (.I0(n33_adj_4505), .I1(n46_adj_4504), .I2(n42_adj_4503), 
            .I3(n34_adj_4502), .O(n2819));
    defparam i23_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i20676_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n25936));
    defparam i20676_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut_adj_1508 (.I0(n2303), .I1(n2295), .I2(n2298), .I3(n25936), 
            .O(n30_adj_4506));
    defparam i11_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1509 (.I0(n2307), .I1(n30_adj_4506), .I2(n2296), 
            .I3(n2300), .O(n34_adj_4507));
    defparam i15_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1510 (.I0(n2304), .I1(n2305), .I2(n2299), .I3(n2302), 
            .O(n32_adj_4508));
    defparam i13_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1511 (.I0(n2293), .I1(n2308), .I2(n2294), .I3(n2297), 
            .O(n33_adj_4509));
    defparam i14_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1512 (.I0(n2301), .I1(n2291), .I2(n2306), .I3(n2292), 
            .O(n31_adj_4510));
    defparam i12_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1513 (.I0(n31_adj_4510), .I1(n33_adj_4509), .I2(n32_adj_4508), 
            .I3(n34_adj_4507), .O(n2324));
    defparam i18_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i41899_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49800));
    defparam i41899_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut (.I0(n2202), .I1(n2206), .I2(n2199), .I3(n2208), 
            .O(n28_adj_4511));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1514 (.I0(n2193), .I1(n28_adj_4511), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4512));
    defparam i14_4_lut_adj_1514.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1515 (.I0(n2198), .I1(n2201), .I2(n2207), .I3(n2197), 
            .O(n30_adj_4513));
    defparam i12_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1516 (.I0(n2205), .I1(n2203), .I2(n2194), .I3(n2200), 
            .O(n31_adj_4514));
    defparam i13_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1517 (.I0(n2196), .I1(n2195), .I2(n2192), .I3(n2204), 
            .O(n29_adj_4515));
    defparam i11_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1518 (.I0(n29_adj_4515), .I1(n31_adj_4514), .I2(n30_adj_4513), 
            .I3(n32_adj_4512), .O(n2225));
    defparam i17_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i41898_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49799));
    defparam i41898_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i41896_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49797));
    defparam i41896_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4516));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'heeee;
    SB_LUT4 i20667_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n25927));
    defparam i20667_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1520 (.I0(n2098), .I1(n2102), .I2(n2100), .I3(n18_adj_4516), 
            .O(n30_adj_4517));
    defparam i13_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1521 (.I0(n2108), .I1(n2099), .I2(n2107), .I3(n25927), 
            .O(n28_adj_4518));
    defparam i11_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1522 (.I0(n2094), .I1(n2096), .I2(n2093), .I3(n2101), 
            .O(n29_adj_4519));
    defparam i12_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1523 (.I0(n2105), .I1(n2106), .I2(n2104), .I3(n2095), 
            .O(n27_adj_4520));
    defparam i10_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_41987 (.I0(bit_ctr[0]), .I1(\color[6] ), 
            .I2(\color[7] ), .I3(bit_ctr[1]), .O(n49901));
    defparam bit_ctr_0__bdd_4_lut_41987.LUT_INIT = 16'he4aa;
    SB_LUT4 n49901_bdd_4_lut (.I0(n49901), .I1(\color[5] ), .I2(\color[4] ), 
            .I3(bit_ctr[1]), .O(n44401));
    defparam n49901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16_4_lut_adj_1524 (.I0(n27_adj_4520), .I1(n29_adj_4519), .I2(n28_adj_4518), 
            .I3(n30_adj_4517), .O(n2126));
    defparam i16_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i41897_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49798));
    defparam i41897_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1525 (.I0(n1999), .I1(n2008), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4521));
    defparam i2_2_lut_adj_1525.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1526 (.I0(n2005), .I1(n1995), .I2(n2002), .I3(n2007), 
            .O(n28_adj_4522));
    defparam i12_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1527 (.I0(n1997), .I1(n1998), .I2(n2006), .I3(n2000), 
            .O(n26_adj_4523));
    defparam i10_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1528 (.I0(n1994), .I1(n2001), .I2(n2004), .I3(n1996), 
            .O(n27_adj_4524));
    defparam i11_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1529 (.I0(bit_ctr[15]), .I1(n18_adj_4521), .I2(n2003), 
            .I3(n2009), .O(n25_adj_4525));
    defparam i9_4_lut_adj_1529.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1530 (.I0(n25_adj_4525), .I1(n27_adj_4524), .I2(n26_adj_4523), 
            .I3(n28_adj_4522), .O(n2027));
    defparam i15_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i41895_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49796));
    defparam i41895_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut_adj_1531 (.I0(n2699), .I1(n2687), .I2(n2689), .I3(n2708), 
            .O(n36_adj_4526));
    defparam i13_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1532 (.I0(n2701), .I1(n2695), .I2(n2704), .I3(n2694), 
            .O(n40_adj_4527));
    defparam i17_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[8]), .I1(n2698), .I2(n2709), .I3(GND_net), 
            .O(n31_adj_4528));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1533 (.I0(n2692), .I1(n2688), .I2(n2690), .I3(n2693), 
            .O(n38_adj_4529));
    defparam i15_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1534 (.I0(n2707), .I1(n2691), .I2(n2700), .I3(n2702), 
            .O(n37_adj_4530));
    defparam i14_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1535 (.I0(n2697), .I1(n36_adj_4526), .I2(n2705), 
            .I3(n2706), .O(n41_adj_4531));
    defparam i18_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1536 (.I0(n31_adj_4528), .I1(n40_adj_4527), .I2(n2696), 
            .I3(n2703), .O(n43_adj_4532));
    defparam i20_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1537 (.I0(n43_adj_4532), .I1(n41_adj_4531), .I2(n37_adj_4530), 
            .I3(n38_adj_4529), .O(n2720));
    defparam i22_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1538 (.I0(n1903), .I1(n1899), .I2(n1895), .I3(n1896), 
            .O(n26_adj_4533));
    defparam i11_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1539 (.I0(n1898), .I1(n1902), .I2(n1906), .I3(n1907), 
            .O(n24_adj_4534));
    defparam i9_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1540 (.I0(n1904), .I1(n1905), .I2(n1901), .I3(n1897), 
            .O(n25_adj_4535));
    defparam i10_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1541 (.I0(n1908), .I1(bit_ctr[16]), .I2(n1900), 
            .I3(n1909), .O(n23_adj_4536));
    defparam i8_4_lut_adj_1541.LUT_INIT = 16'hfefa;
    SB_LUT4 i14_4_lut_adj_1542 (.I0(n23_adj_4536), .I1(n25_adj_4535), .I2(n24_adj_4534), 
            .I3(n26_adj_4533), .O(n1928));
    defparam i14_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i41894_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49795));
    defparam i41894_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1543 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4537));
    defparam i10_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1544 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4538));
    defparam i8_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1545 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4539));
    defparam i9_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1546 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4540));
    defparam i7_3_lut_adj_1546.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1547 (.I0(n21_adj_4540), .I1(n23_adj_4539), .I2(n22_adj_4538), 
            .I3(n24_adj_4537), .O(n1829));
    defparam i13_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i41893_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49794));
    defparam i41893_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_41982 (.I0(bit_ctr[0]), .I1(\color[10] ), 
            .I2(\color[11] ), .I3(bit_ctr[1]), .O(n49895));
    defparam bit_ctr_0__bdd_4_lut_41982.LUT_INIT = 16'he4aa;
    SB_LUT4 n49895_bdd_4_lut (.I0(n49895), .I1(\color[9] ), .I2(\color[8] ), 
            .I3(bit_ctr[1]), .O(n44404));
    defparam n49895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1548 (.I0(start), .I1(\state[1] ), .I2(n116), 
            .I3(GND_net), .O(n4_adj_4481));
    defparam i1_2_lut_3_lut_adj_1548.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(n26050), .I3(\state[0] ), .O(n44172));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i2_2_lut_3_lut (.I0(n29), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n41777));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n26074), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n37493));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n26074), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_LUT4 i1_2_lut_4_lut (.I0(one_wire_N_399[4]), .I1(one_wire_N_399[2]), 
            .I2(one_wire_N_399[3]), .I3(n116), .O(n17574));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff80;
    SB_LUT4 i1_2_lut_4_lut_adj_1549 (.I0(n1), .I1(one_wire_N_399[9]), .I2(one_wire_N_399[5]), 
            .I3(one_wire_N_399[6]), .O(n116));
    defparam i1_2_lut_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_41977 (.I0(bit_ctr[0]), .I1(\color[18] ), 
            .I2(\color[19] ), .I3(bit_ctr[1]), .O(n49865));
    defparam bit_ctr_0__bdd_4_lut_41977.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_4_lut (.I0(one_wire_N_399[6]), .I1(one_wire_N_399[5]), 
            .I2(one_wire_N_399[9]), .I3(n1), .O(n6_adj_4448));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3554_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n42530), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3554_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 i9_4_lut_adj_1550 (.I0(n1707), .I1(n1697), .I2(n1702), .I3(n1703), 
            .O(n22_adj_4541));
    defparam i9_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1551 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4542));
    defparam i7_3_lut_adj_1551.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_4_lut_adj_1552 (.I0(n1698), .I1(n1700), .I2(n1705), .I3(n1706), 
            .O(n21_adj_4543));
    defparam i8_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n19_adj_4544));
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i12_4_lut_adj_1553 (.I0(n19_adj_4544), .I1(n21_adj_4543), .I2(n20_adj_4542), 
            .I3(n22_adj_4541), .O(n1730));
    defparam i12_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 n49865_bdd_4_lut (.I0(n49865), .I1(\color[17] ), .I2(\color[16] ), 
            .I3(bit_ctr[1]), .O(n49868));
    defparam n49865_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i41892_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49793));
    defparam i41892_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_41953 (.I0(bit_ctr[0]), .I1(\color[14] ), 
            .I2(\color[15] ), .I3(bit_ctr[1]), .O(n49829));
    defparam bit_ctr_0__bdd_4_lut_41953.LUT_INIT = 16'he4aa;
    SB_LUT4 n49829_bdd_4_lut (.I0(n49829), .I1(\color[13] ), .I2(\color[12] ), 
            .I3(bit_ctr[1]), .O(n48564));
    defparam n49829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1554 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4545));
    defparam i8_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1555 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4546));
    defparam i1_3_lut_adj_1555.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4547));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1556 (.I0(n13_adj_4546), .I1(n20_adj_4545), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4548));
    defparam i10_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1557 (.I0(n1601), .I1(n22_adj_4548), .I2(n18_adj_4547), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i41891_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49792));
    defparam i41891_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i41890_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49791));
    defparam i41890_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1558 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4549));
    defparam i7_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1559 (.I0(n1504), .I1(n18_adj_4549), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4550));
    defparam i9_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), .I3(GND_net), 
            .O(n15_adj_4551));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1560 (.I0(n15_adj_4551), .I1(n20_adj_4550), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n41871));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34666_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n26074), .I2(n608), 
            .I3(bit_ctr[29]), .O(n42547));
    defparam i34666_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n44404), .I2(n48564), 
            .I3(color_bit_N_442[3]), .O(n49805));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49805_bdd_4_lut (.I0(n49805), .I1(n44401), .I2(n44398), .I3(color_bit_N_442[3]), 
            .O(n49808));
    defparam n49805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20809_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n26074));
    defparam i20809_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i39352_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17743));
    defparam i39352_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_LUT4 i14_4_lut_adj_1561 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4552));
    defparam i14_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1562 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4553));
    defparam i3_3_lut_adj_1562.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1563 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4554));
    defparam i12_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1564 (.I0(n25_adj_4553), .I1(n36_adj_4552), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4555));
    defparam i18_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1565 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4556));
    defparam i16_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4554), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4557));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1566 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4558));
    defparam i15_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1567 (.I0(n37_adj_4558), .I1(n39_adj_4557), .I2(n38_adj_4556), 
            .I3(n40_adj_4555), .O(n2621));
    defparam i21_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i41889_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n49790));
    defparam i41889_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n18531, encoder0_position, clk32MHz, 
            n18530, n18529, n18528, n18527, n18526, n18525, n18524, 
            n18523, n18522, n18521, n18520, n18519, n18518, n18517, 
            n18516, n18515, n18514, n18513, n18512, n18511, n18510, 
            n18497, data_o, n2642, GND_net, n17969, count_enable, 
            n18616, reg_B, PIN_23_c_1, PIN_24_c_0, n17971, n44088) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18531;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n18530;
    input n18529;
    input n18528;
    input n18527;
    input n18526;
    input n18525;
    input n18524;
    input n18523;
    input n18522;
    input n18521;
    input n18520;
    input n18519;
    input n18518;
    input n18517;
    input n18516;
    input n18515;
    input n18514;
    input n18513;
    input n18512;
    input n18511;
    input n18510;
    input n18497;
    output [1:0]data_o;
    output [23:0]n2642;
    input GND_net;
    input n17969;
    output count_enable;
    input n18616;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n17971;
    output n44088;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire B_delayed, A_delayed, n2638, n34648, n34647, n34646, n34645, 
        n34644, n34643, n34642, n34641, n34640, n34639, n34638, 
        n34637, n34636, n34635, n34634, n34633, n34632, n34631, 
        n34630, n34629, n34628, n34627, n34626, count_direction, 
        n34625;
    
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n18531));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n18530));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n18529));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n18528));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n18527));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n18526));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n18525));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n18524));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n18523));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n18522));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n18521));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n18520));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n18519));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n18518));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n18517));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n18516));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n18515));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n18514));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n18513));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n18512));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n18511));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n18510));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n18497));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_625_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2638), 
            .I3(n34648), .O(n2642[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_625_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2638), 
            .I3(n34647), .O(n2642[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_24 (.CI(n34647), .I0(encoder0_position[22]), .I1(n2638), 
            .CO(n34648));
    SB_LUT4 add_625_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2638), 
            .I3(n34646), .O(n2642[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_23 (.CI(n34646), .I0(encoder0_position[21]), .I1(n2638), 
            .CO(n34647));
    SB_LUT4 add_625_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2638), 
            .I3(n34645), .O(n2642[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_22 (.CI(n34645), .I0(encoder0_position[20]), .I1(n2638), 
            .CO(n34646));
    SB_LUT4 add_625_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2638), 
            .I3(n34644), .O(n2642[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_21 (.CI(n34644), .I0(encoder0_position[19]), .I1(n2638), 
            .CO(n34645));
    SB_LUT4 add_625_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2638), 
            .I3(n34643), .O(n2642[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_20 (.CI(n34643), .I0(encoder0_position[18]), .I1(n2638), 
            .CO(n34644));
    SB_LUT4 add_625_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2638), 
            .I3(n34642), .O(n2642[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_19 (.CI(n34642), .I0(encoder0_position[17]), .I1(n2638), 
            .CO(n34643));
    SB_LUT4 add_625_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2638), 
            .I3(n34641), .O(n2642[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_18 (.CI(n34641), .I0(encoder0_position[16]), .I1(n2638), 
            .CO(n34642));
    SB_LUT4 add_625_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2638), 
            .I3(n34640), .O(n2642[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_17 (.CI(n34640), .I0(encoder0_position[15]), .I1(n2638), 
            .CO(n34641));
    SB_LUT4 add_625_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2638), 
            .I3(n34639), .O(n2642[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_16 (.CI(n34639), .I0(encoder0_position[14]), .I1(n2638), 
            .CO(n34640));
    SB_LUT4 add_625_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2638), 
            .I3(n34638), .O(n2642[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_15 (.CI(n34638), .I0(encoder0_position[13]), .I1(n2638), 
            .CO(n34639));
    SB_LUT4 add_625_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2638), 
            .I3(n34637), .O(n2642[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_14 (.CI(n34637), .I0(encoder0_position[12]), .I1(n2638), 
            .CO(n34638));
    SB_LUT4 add_625_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2638), 
            .I3(n34636), .O(n2642[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_13 (.CI(n34636), .I0(encoder0_position[11]), .I1(n2638), 
            .CO(n34637));
    SB_LUT4 add_625_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2638), 
            .I3(n34635), .O(n2642[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_12 (.CI(n34635), .I0(encoder0_position[10]), .I1(n2638), 
            .CO(n34636));
    SB_LUT4 add_625_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2638), 
            .I3(n34634), .O(n2642[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_11 (.CI(n34634), .I0(encoder0_position[9]), .I1(n2638), 
            .CO(n34635));
    SB_LUT4 add_625_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2638), 
            .I3(n34633), .O(n2642[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_10 (.CI(n34633), .I0(encoder0_position[8]), .I1(n2638), 
            .CO(n34634));
    SB_LUT4 add_625_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2638), 
            .I3(n34632), .O(n2642[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_9 (.CI(n34632), .I0(encoder0_position[7]), .I1(n2638), 
            .CO(n34633));
    SB_LUT4 add_625_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2638), 
            .I3(n34631), .O(n2642[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_8 (.CI(n34631), .I0(encoder0_position[6]), .I1(n2638), 
            .CO(n34632));
    SB_LUT4 add_625_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2638), 
            .I3(n34630), .O(n2642[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_7 (.CI(n34630), .I0(encoder0_position[5]), .I1(n2638), 
            .CO(n34631));
    SB_LUT4 add_625_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2638), 
            .I3(n34629), .O(n2642[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_6 (.CI(n34629), .I0(encoder0_position[4]), .I1(n2638), 
            .CO(n34630));
    SB_LUT4 add_625_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2638), 
            .I3(n34628), .O(n2642[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_5 (.CI(n34628), .I0(encoder0_position[3]), .I1(n2638), 
            .CO(n34629));
    SB_LUT4 add_625_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2638), 
            .I3(n34627), .O(n2642[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_4 (.CI(n34627), .I0(encoder0_position[2]), .I1(n2638), 
            .CO(n34628));
    SB_LUT4 add_625_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2638), 
            .I3(n34626), .O(n2642[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_3 (.CI(n34626), .I0(encoder0_position[1]), .I1(n2638), 
            .CO(n34627));
    SB_LUT4 add_625_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n34625), .O(n2642[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_625_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_625_2 (.CI(n34625), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n34626));
    SB_CARRY add_625_1 (.CI(GND_net), .I0(n2638), .I1(n2638), .CO(n34625));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17969));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i917_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // quad.v(37[5] 40[8])
    defparam i917_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n18616(n18616), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .PIN_23_c_1(PIN_23_c_1), 
            .PIN_24_c_0(PIN_24_c_0), .n17971(n17971), .n44088(n44088), 
            .GND_net(GND_net)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18616, data_o, clk32MHz, reg_B, PIN_23_c_1, 
            PIN_24_c_0, n17971, n44088, GND_net) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18616;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n17971;
    output n44088;
    input GND_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n1;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3463;
    wire [2:0]n17;
    
    wire n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18616));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_23_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1193__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n1), .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_24_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1193__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1193__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17971));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n44088));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i28881_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i28881_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i28874_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i28874_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44088), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i1443_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i1443_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=48, LSE_LCOL=12, LSE_RCOL=39, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n23171, PWMLimit, clk32MHz, n18460, n18459, n18458, 
            n18457, GND_net, n18456, n18455, n18454, n18453, n18452, 
            n18451, n18450, n18449, n18448, control_mode, rx_data, 
            \data_in_frame[9] , n18447, \data_in_frame[19] , \data_in_frame[14] , 
            \data_in_frame[13] , \data_in_frame[8] , n18329, \data_in_frame[7] , 
            n18328, n18327, n18326, n18325, n18324, n18323, n18369, 
            \data_in_frame[12] , n18667, setpoint, n18666, n18665, 
            n18664, n18663, n18662, n18661, n18660, n18659, n18658, 
            n18657, n18656, n18655, n18654, n18653, n18652, n18651, 
            n18650, n18649, n18648, n18647, n18646, n18645, n18368, 
            n18367, n18366, n18365, n18593, VCC_net, byte_transmit_counter, 
            n18364, n18363, n18362, \data_in_frame[11] , n18550, n18547, 
            n18544, n18541, n18538, n18535, n18509, n50009, \data_in_frame[10] , 
            n18471, n18470, n18469, n18468, n18467, n18466, n23694, 
            n18464, n18463, n18462, n18322, \data_in_frame[6] , \data_in_frame[18] , 
            \data_in_frame[17] , \data_in_frame[5] , n18305, \data_in_frame[4] , 
            n18304, n18303, n18302, n18301, n18300, n18299, n18298, 
            rx_data_ready, \data_in_frame[3] , n18446, n18445, n18444, 
            n18443, n18442, \data_in_frame[2] , \FRAME_MATCHER.state[3] , 
            \FRAME_MATCHER.state[0] , \data_in_frame[1] , Kp_23__N_679, 
            n17503, n37696, n43448, n18266, \data_out_frame[20] , 
            n18265, n18264, n18263, n18262, n18261, n18260, n18259, 
            n18258, \data_out_frame[19] , n18257, n18256, n18255, 
            n18254, n18253, n18252, n18251, n18250, \data_out_frame[18] , 
            n18249, n18248, n18247, n18246, n18245, n18244, n18243, 
            n18242, \data_out_frame[17] , n18241, n18240, n18239, 
            n18238, n18237, n18236, n18235, n18234, \data_out_frame[16] , 
            n18233, n18232, n18231, n41851, n18230, n2857, n41860, 
            n18229, n18228, n18227, n18226, \data_out_frame[15] , 
            n18225, n18224, n18223, n18222, n18221, n18220, n18219, 
            n18218, \data_out_frame[14] , n18217, n18216, n18215, 
            n18214, n18213, n18212, n18211, n18210, \data_out_frame[13] , 
            n18209, n18208, n18207, n18206, n18205, n18204, n18203, 
            n16563, \data_out_frame[5] , \data_out_frame[6] , \data_out_frame[7] , 
            \data_in_frame[20] , \data_in_frame[15] , n18202, \data_out_frame[12] , 
            n18201, n41862, n18507, n4497, n18200, n18199, n18198, 
            n18197, n18196, n18195, n18194, \data_out_frame[11] , 
            n18193, n18192, n18191, n18190, n18189, n18188, n18187, 
            n18186, \data_out_frame[10] , n18185, n18184, n18183, 
            n18533, n18182, n18181, n18180, n18179, n18178, \data_out_frame[9] , 
            n18177, n18176, n18175, n18174, n18173, n18172, n18171, 
            n18170, \data_out_frame[8] , n18169, n18168, n18167, n18536, 
            n18166, n18165, n18164, n18163, n41848, n41857, n18162, 
            n18161, n18160, n18159, n18158, n18157, n18156, n18155, 
            n18154, n18153, n18152, n18151, n18150, n18149, n18148, 
            n18147, n18146, n18145, n18144, n18143, n18393, n18392, 
            n18391, n18390, n18539, n18389, n17862, deadband, n37561, 
            n18433, n18432, n18431, n18430, n18429, n18428, n18427, 
            n18426, n38230, n42079, n37512, n18542, n18545, n18548, 
            n2244, n18142, n18141, n18388, n18387, n18386, n18140, 
            n18139, n18135, \data_in[3] , n18134, n18133, n18132, 
            n18131, n18130, n18129, n18128, n18127, \data_in[2] , 
            n18126, n18125, n18124, n18123, n18122, n18121, n18120, 
            n18119, \data_in[1] , n18118, n18117, n18116, n18115, 
            n18114, n18113, n18112, n18111, \data_in[0] , n18110, 
            n18109, n18108, n18107, n18106, n18105, n18104, gearBoxRatio, 
            n18103, n18102, n18101, n18100, n18099, n18098, n18097, 
            n18096, n18095, n18094, n18093, n18092, n18091, n18090, 
            n18089, n18088, n18087, n18086, n18085, n18084, n18083, 
            n18082, n18081, \Kd[7] , n18080, \Kd[6] , n18079, \Kd[5] , 
            n18078, \Kd[4] , n18077, \Kd[3] , n18076, \Kd[2] , n18075, 
            \Kd[1] , n18074, \Ki[7] , n18073, \Ki[6] , n18072, \Ki[5] , 
            n18071, \Ki[4] , n18070, \Ki[3] , n18069, \Ki[2] , n18068, 
            \Ki[1] , n18067, \Kp[7] , n18066, \Kp[6] , n18065, \Kp[5] , 
            n18064, \Kp[4] , n18063, \Kp[3] , n18062, \Kp[2] , n18061, 
            \Kp[1] , n18060, IntegralLimit, n18059, n18058, n18057, 
            n18056, n18055, n18054, n18053, n18052, n18051, n18050, 
            n18049, n18048, n18047, n18046, n18045, n18044, n18043, 
            n18042, n18041, n18040, n18039, n18038, n18013, n18012, 
            n18011, n18010, n18009, n18008, n18007, n18006, n18005, 
            n18004, n18003, n18002, n18001, n18000, n17999, n17998, 
            n17997, n17996, n17995, n17994, n17993, n17992, n17991, 
            n17983, n40968, n17966, n17965, n17963, n17962, n17961, 
            \Kd[0] , n17960, \Ki[0] , n17959, \Kp[0] , n17958, LED_c, 
            n123, n740, n19921, n16687, n16678, n2484, n16680, 
            n5, n7, n50704, n41916, n28, n42216, n37, n42140, 
            n42342, n42357, n14246, n16683, n42066, n42219, n42330, 
            n42459, n42429, n43056, n15, n13, n14, n42432, n25520, 
            n4446, n4447, n4448, n4449, n4450, n14276, n3, n16675, 
            n6, n4451, n4452, n17283, n4453, n4454, n4455, n4456, 
            n4457, n4458, n4459, n4460, n4461, n42696, n4462, 
            n4463, n4464, n42610, n4465, n4466, n4467, n4469, 
            n4468, n5_adj_15, n4, n19, n41336, n41446, n41444, 
            n41442, n41074, \r_Clock_Count[8] , n41130, \r_Clock_Count[7] , 
            n41224, \r_Clock_Count[6] , n41348, tx_o, tx_enable, n88, 
            n118, \r_SM_Main[2] , n5_adj_16, n44294, n17955, n17977, 
            n17980, n17863, n17866, n17869, n17872, n18575, n17974, 
            n3_adj_17, n17887, r_Bit_Index, n17890, n18701, \r_Clock_Count[0] , 
            r_SM_Main, n18587, n41150, n18583, n18567, \r_Clock_Count[5] , 
            n18555, \r_Clock_Count[1] , \r_SM_Main_2__N_3032[2] , r_Rx_Data, 
            PIN_13_N_50, n27708, n17657, n17707, n17849, n4694, 
            n221, n225, n226, n17897, n17896, n17895, n17894, 
            n17893, n17892, n17891, n16566, n4_adj_19, n25329, n4_adj_20, 
            n4_adj_21, n16432) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n23171;
    output [23:0]PWMLimit;
    input clk32MHz;
    input n18460;
    input n18459;
    input n18458;
    input n18457;
    input GND_net;
    input n18456;
    input n18455;
    input n18454;
    input n18453;
    input n18452;
    input n18451;
    input n18450;
    input n18449;
    input n18448;
    output [7:0]control_mode;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[9] ;
    input n18447;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[8] ;
    input n18329;
    output [7:0]\data_in_frame[7] ;
    input n18328;
    input n18327;
    input n18326;
    input n18325;
    input n18324;
    input n18323;
    input n18369;
    output [7:0]\data_in_frame[12] ;
    input n18667;
    output [23:0]setpoint;
    input n18666;
    input n18665;
    input n18664;
    input n18663;
    input n18662;
    input n18661;
    input n18660;
    input n18659;
    input n18658;
    input n18657;
    input n18656;
    input n18655;
    input n18654;
    input n18653;
    input n18652;
    input n18651;
    input n18650;
    input n18649;
    input n18648;
    input n18647;
    input n18646;
    input n18645;
    input n18368;
    input n18367;
    input n18366;
    input n18365;
    input n18593;
    input VCC_net;
    output [7:0]byte_transmit_counter;
    input n18364;
    input n18363;
    input n18362;
    output [7:0]\data_in_frame[11] ;
    input n18550;
    input n18547;
    input n18544;
    input n18541;
    input n18538;
    input n18535;
    input n18509;
    input n50009;
    output [7:0]\data_in_frame[10] ;
    input n18471;
    input n18470;
    input n18469;
    input n18468;
    input n18467;
    input n18466;
    input n23694;
    input n18464;
    input n18463;
    input n18462;
    input n18322;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[5] ;
    input n18305;
    output [7:0]\data_in_frame[4] ;
    input n18304;
    input n18303;
    input n18302;
    input n18301;
    input n18300;
    input n18299;
    input n18298;
    output rx_data_ready;
    output [7:0]\data_in_frame[3] ;
    input n18446;
    input n18445;
    input n18444;
    input n18443;
    input n18442;
    output [7:0]\data_in_frame[2] ;
    output \FRAME_MATCHER.state[3] ;
    output \FRAME_MATCHER.state[0] ;
    output [7:0]\data_in_frame[1] ;
    output Kp_23__N_679;
    output n17503;
    output n37696;
    output n43448;
    input n18266;
    output [7:0]\data_out_frame[20] ;
    input n18265;
    input n18264;
    input n18263;
    input n18262;
    input n18261;
    input n18260;
    input n18259;
    input n18258;
    output [7:0]\data_out_frame[19] ;
    input n18257;
    input n18256;
    input n18255;
    input n18254;
    input n18253;
    input n18252;
    input n18251;
    input n18250;
    output [7:0]\data_out_frame[18] ;
    input n18249;
    input n18248;
    input n18247;
    input n18246;
    input n18245;
    input n18244;
    input n18243;
    input n18242;
    output [7:0]\data_out_frame[17] ;
    input n18241;
    input n18240;
    input n18239;
    input n18238;
    input n18237;
    input n18236;
    input n18235;
    input n18234;
    output [7:0]\data_out_frame[16] ;
    input n18233;
    input n18232;
    input n18231;
    output n41851;
    input n18230;
    output n2857;
    output n41860;
    input n18229;
    input n18228;
    input n18227;
    input n18226;
    output [7:0]\data_out_frame[15] ;
    input n18225;
    input n18224;
    input n18223;
    input n18222;
    input n18221;
    input n18220;
    input n18219;
    input n18218;
    output [7:0]\data_out_frame[14] ;
    input n18217;
    input n18216;
    input n18215;
    input n18214;
    input n18213;
    input n18212;
    input n18211;
    input n18210;
    output [7:0]\data_out_frame[13] ;
    input n18209;
    input n18208;
    input n18207;
    input n18206;
    input n18205;
    input n18204;
    input n18203;
    output n16563;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[20] ;
    output [7:0]\data_in_frame[15] ;
    input n18202;
    output [7:0]\data_out_frame[12] ;
    input n18201;
    output n41862;
    output n18507;
    output n4497;
    input n18200;
    input n18199;
    input n18198;
    input n18197;
    input n18196;
    input n18195;
    input n18194;
    output [7:0]\data_out_frame[11] ;
    input n18193;
    input n18192;
    input n18191;
    input n18190;
    input n18189;
    input n18188;
    input n18187;
    input n18186;
    output [7:0]\data_out_frame[10] ;
    input n18185;
    input n18184;
    input n18183;
    output n18533;
    input n18182;
    input n18181;
    input n18180;
    input n18179;
    input n18178;
    output [7:0]\data_out_frame[9] ;
    input n18177;
    input n18176;
    input n18175;
    input n18174;
    input n18173;
    input n18172;
    input n18171;
    input n18170;
    output [7:0]\data_out_frame[8] ;
    input n18169;
    input n18168;
    input n18167;
    output n18536;
    input n18166;
    input n18165;
    input n18164;
    input n18163;
    output n41848;
    output n41857;
    input n18162;
    input n18161;
    input n18160;
    input n18159;
    input n18158;
    input n18157;
    input n18156;
    input n18155;
    input n18154;
    input n18153;
    input n18152;
    input n18151;
    input n18150;
    input n18149;
    input n18148;
    input n18147;
    input n18146;
    input n18145;
    input n18144;
    input n18143;
    input n18393;
    input n18392;
    input n18391;
    input n18390;
    output n18539;
    input n18389;
    input n17862;
    output [23:0]deadband;
    input n37561;
    input n18433;
    input n18432;
    input n18431;
    input n18430;
    input n18429;
    input n18428;
    input n18427;
    input n18426;
    output n38230;
    input n42079;
    output n37512;
    output n18542;
    output n18545;
    output n18548;
    output n2244;
    input n18142;
    input n18141;
    input n18388;
    input n18387;
    input n18386;
    input n18140;
    input n18139;
    input n18135;
    output [7:0]\data_in[3] ;
    input n18134;
    input n18133;
    input n18132;
    input n18131;
    input n18130;
    input n18129;
    input n18128;
    input n18127;
    output [7:0]\data_in[2] ;
    input n18126;
    input n18125;
    input n18124;
    input n18123;
    input n18122;
    input n18121;
    input n18120;
    input n18119;
    output [7:0]\data_in[1] ;
    input n18118;
    input n18117;
    input n18116;
    input n18115;
    input n18114;
    input n18113;
    input n18112;
    input n18111;
    output [7:0]\data_in[0] ;
    input n18110;
    input n18109;
    input n18108;
    input n18107;
    input n18106;
    input n18105;
    input n18104;
    output [23:0]gearBoxRatio;
    input n18103;
    input n18102;
    input n18101;
    input n18100;
    input n18099;
    input n18098;
    input n18097;
    input n18096;
    input n18095;
    input n18094;
    input n18093;
    input n18092;
    input n18091;
    input n18090;
    input n18089;
    input n18088;
    input n18087;
    input n18086;
    input n18085;
    input n18084;
    input n18083;
    input n18082;
    input n18081;
    output \Kd[7] ;
    input n18080;
    output \Kd[6] ;
    input n18079;
    output \Kd[5] ;
    input n18078;
    output \Kd[4] ;
    input n18077;
    output \Kd[3] ;
    input n18076;
    output \Kd[2] ;
    input n18075;
    output \Kd[1] ;
    input n18074;
    output \Ki[7] ;
    input n18073;
    output \Ki[6] ;
    input n18072;
    output \Ki[5] ;
    input n18071;
    output \Ki[4] ;
    input n18070;
    output \Ki[3] ;
    input n18069;
    output \Ki[2] ;
    input n18068;
    output \Ki[1] ;
    input n18067;
    output \Kp[7] ;
    input n18066;
    output \Kp[6] ;
    input n18065;
    output \Kp[5] ;
    input n18064;
    output \Kp[4] ;
    input n18063;
    output \Kp[3] ;
    input n18062;
    output \Kp[2] ;
    input n18061;
    output \Kp[1] ;
    input n18060;
    output [23:0]IntegralLimit;
    input n18059;
    input n18058;
    input n18057;
    input n18056;
    input n18055;
    input n18054;
    input n18053;
    input n18052;
    input n18051;
    input n18050;
    input n18049;
    input n18048;
    input n18047;
    input n18046;
    input n18045;
    input n18044;
    input n18043;
    input n18042;
    input n18041;
    input n18040;
    input n18039;
    input n18038;
    input n18013;
    input n18012;
    input n18011;
    input n18010;
    input n18009;
    input n18008;
    input n18007;
    input n18006;
    input n18005;
    input n18004;
    input n18003;
    input n18002;
    input n18001;
    input n18000;
    input n17999;
    input n17998;
    input n17997;
    input n17996;
    input n17995;
    input n17994;
    input n17993;
    input n17992;
    input n17991;
    input n17983;
    input n40968;
    input n17966;
    input n17965;
    input n17963;
    input n17962;
    input n17961;
    output \Kd[0] ;
    input n17960;
    output \Ki[0] ;
    input n17959;
    output \Kp[0] ;
    input n17958;
    output LED_c;
    output n123;
    output n740;
    output n19921;
    output n16687;
    output n16678;
    output n2484;
    output n16680;
    output n5;
    output n7;
    output n50704;
    input n41916;
    input n28;
    input n42216;
    input n37;
    output n42140;
    output n42342;
    output n42357;
    output n14246;
    output n16683;
    input n42066;
    input n42219;
    input n42330;
    output n42459;
    input n42429;
    output n43056;
    input n15;
    input n13;
    input n14;
    output n42432;
    output n25520;
    output n4446;
    output n4447;
    output n4448;
    output n4449;
    output n4450;
    output n14276;
    output n3;
    output n16675;
    output n6;
    output n4451;
    output n4452;
    output n17283;
    output n4453;
    output n4454;
    output n4455;
    output n4456;
    output n4457;
    output n4458;
    output n4459;
    output n4460;
    output n4461;
    output n42696;
    output n4462;
    output n4463;
    output n4464;
    output n42610;
    output n4465;
    output n4466;
    output n4467;
    output n4469;
    output n4468;
    output n5_adj_15;
    input n4;
    input n19;
    input n41336;
    input n41446;
    input n41444;
    input n41442;
    input n41074;
    output \r_Clock_Count[8] ;
    input n41130;
    output \r_Clock_Count[7] ;
    input n41224;
    output \r_Clock_Count[6] ;
    input n41348;
    output tx_o;
    output tx_enable;
    output n88;
    output n118;
    output \r_SM_Main[2] ;
    input n5_adj_16;
    output n44294;
    output n17955;
    output n17977;
    output n17980;
    output n17863;
    output n17866;
    output n17869;
    output n17872;
    output n18575;
    input n17974;
    output n3_adj_17;
    input n17887;
    output [2:0]r_Bit_Index;
    input n17890;
    input n18701;
    output \r_Clock_Count[0] ;
    output [2:0]r_SM_Main;
    input n18587;
    input n41150;
    input n18583;
    input n18567;
    output \r_Clock_Count[5] ;
    input n18555;
    output \r_Clock_Count[1] ;
    output \r_SM_Main_2__N_3032[2] ;
    output r_Rx_Data;
    input PIN_13_N_50;
    output n27708;
    output n17657;
    output n17707;
    output n17849;
    output n4694;
    output n221;
    output n225;
    output n226;
    input n17897;
    input n17896;
    input n17895;
    input n17894;
    input n17893;
    input n17892;
    input n17891;
    output n16566;
    output n4_adj_19;
    output n25329;
    output n4_adj_20;
    output n4_adj_21;
    output n16432;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n34575;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n34576, n2, n34574, n1774, n2_adj_4113, n3_c, n8, n41852, 
        n18338, n18418, n18379, n18378, n18377, n18376, n18337, 
        n18375, n18374, n18373, n18336, n18335, n18334, n34578, 
        n34579, n18333, n18332, n18331, n18330, n2_adj_4114, n34573, 
        n18372, n2_adj_4115, n34572, n18371, n18370, n18339, n18361, 
        n18360, n18359, n18358, n18340, n23932, n18356, n18355, 
        n18354;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(100[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n18353, n18352, n18321, n18320, n18319, n18318, n18317, 
        n18316, n18315, n18411, n18410, n18409, n18408, n18407, 
        n18406, n18405, n18314, n18313, n18312, n18311, n18310, 
        n18309, n18308, n18307, n18306, n18404, n18403, n18402, 
        n18401;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n18400, n18399, n18341, n18342, n18343, n18344, n18345, 
        n18398, n18397, n8_adj_4116, n41861, n18419, n18351, n18420, 
        n18350, n18421, n18349, n18348, n18347, n18422, n18346, 
        n18417, n2_adj_4117, n34571, \FRAME_MATCHER.rx_data_ready_prev , 
        n18297, n18423, n18424, n18396, n18425, n2_adj_4118, n34570, 
        n18296, n2_adj_4119, n3_adj_4120, n2_adj_4121, n34569, n2_adj_4122, 
        n34568, n8_adj_4123, n18295, n2_adj_4124, n34567, n2_adj_4125, 
        n34566, n10, n41876, n2_adj_4126, n34565, n16608, n16468, 
        n8_adj_4127;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n18439, n41874, n18412, n18294, n18293, n18292, n18291, 
        n18290, n2_adj_4128, n34564, n18289, n2_adj_4129, n34563, 
        n18288, n18287, n25285, n16446, n44325, n16682, n25611, 
        n44377, n44376;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n44374, n44373, n44371, n44370, n31, n25297, n25299;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n4_c, n41996, n41891, n16804, n5_c, n17168, n41993, n16893, 
        n41977, n6_c, n44368, n49964, n16307, n6_adj_4130, n16, 
        Kp_23__N_809, n4_adj_4131, n42229, n17035, n41898, n16898, 
        n42262, n42384, n2_adj_4132, n34562, n6_adj_4133, n16827, 
        n18, n44359, n44358, n44362, n49976, n41999, n41925, n15066, 
        Kp_23__N_676, n16_adj_4134, n17, n44365, n49970, n6_adj_4135, 
        n2_adj_4136, n34561, n41956, n17037, n37571, n43394, n8_adj_4137, 
        n18382, n37621, n15_c, n18383, Kp_23__N_729, n8_adj_4138, 
        n16851, n2_adj_4139, n34560, n16903, n1, n28_c, n16889, 
        n26, n17185, n27, n25, n7_c, n144, n26154, n31_adj_4140, 
        n25630, n13947, n18384;
    wire [7:0]\data_in_frame[14]_c ;   // verilog/coms.v(94[12:25])
    
    wire n18380, n2_adj_4141, n34559, n18286, n2_adj_4142, n34558, 
        n18285, n18385, n18284, n18381, n18283, n18282, n18441, 
        n2_adj_4143, n34557, n18440, n18281, n18280, n24, n18279, 
        n18278, n41843, n2_adj_4144, n34556, n18277, n18276, n18275, 
        n18274, n18273, n18272, n18271, n18270, n18269, n18268, 
        n18267, n3_adj_4145, n34555, n18416, n2_adj_4146, n34554, 
        n22, n18438, n10_adj_4147, n18437, n18395, n18436, n3_adj_4148, 
        n3_adj_4149, n3_adj_4150, n3_adj_4151, n3_adj_4152, n3_adj_4153, 
        n3_adj_4154, n3_adj_4155, n3_adj_4156, n3_adj_4157, n3_adj_4158, 
        n3_adj_4159, n3_adj_4160, n3_adj_4161, n3_adj_4162, n3_adj_4163, 
        n3_adj_4164, n3_adj_4165, n2_adj_4166, n3_adj_4167, n2_adj_4168, 
        n3_adj_4169, n2_adj_4170, n3_adj_4171, n2_adj_4172, n3_adj_4173, 
        n2_adj_4174, n3_adj_4175, n2_adj_4176, n3_adj_4177, n2_adj_4178, 
        n3_adj_4179, n2_adj_4180, n3_adj_4181, n2_adj_4182, n3_adj_4183, 
        n2_adj_4184, n3_adj_4185, n43355, n17676;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n43374, n43377, n44061, n43198, n44072, n43875, n43169, 
        n43711;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n42290, n42412, n43317, n43126, n42174, n43726, n43199, 
        n40980, n50161, n40984, n41172, n41264, n40986, n41266, 
        n41046, n41268, n41044, n41270, n41042, n41282, n41052, 
        n41334, n41060, n41342, n40966, n41344, n41050, n41346, 
        n41040, n7_adj_4186, n8_adj_4187, n7_adj_4188, n8_adj_4189, 
        n7_adj_4190, n8_adj_4191, n41240, n40988, n7_adj_4192, n8_adj_4193, 
        n41242, n41038, n41244, n41036, n41246, n41034, n25288, 
        n41032, n41248, n41030, n7_adj_4194, n25290, n41250, n41028, 
        n41252, n41026, n7_adj_4195, n8_adj_4196, n7_adj_4197, n8_adj_4198, 
        n7_adj_4199, n8_adj_4200, n41254, n40982, n41144, n40964, 
        n7_adj_4201, n8_adj_4202, n26_adj_4203, n25_adj_4204, n14_c, 
        n14_adj_4205, n13_c, n13_adj_4206, n164, n42251, n17415, 
        n42393, n10_adj_4207, n41962, n16971, n43667, n43329, n38220, 
        n18_adj_4208, n19_c, n6_adj_4209, n5_adj_4210, n44379, n18_adj_4211, 
        n30, n49952, n44380, n45195, n44357, n17325, n42408, n28_adj_4212, 
        n49946, n49862, n42372, n42447, n42167, n27_adj_4213, n34553, 
        n34552, n34551, n46769;
    wire [2:0]r_SM_Main_2__N_3106;
    
    wire n42491, n18394, n18415, n49985, n49988, n44336, n44337, 
        n49973, n44334, n44333, n44342, n44343, n49967, n44340, 
        n44339, n44348, n44349, n49961, n44346, n44345, n49955, 
        n49958, n49949, n42097, n16750, n42308, n10_adj_4214, n16268, 
        n38270, n42070, n18414, n34550, n49943, n18435, n42345, 
        n6_adj_4215, n18434, n42152, n43335, n42179, n43390, n42351, 
        n10_adj_4216, n37587, n8_adj_4217, n42149, n43441, Kp_23__N_1213, 
        n37485, n43365, n22_adj_4218, n41959, n42245, n42959, n42076, 
        n44278, n42825, n42158, n27_adj_4219, n42390, Kp_23__N_1201, 
        n42188, n14_adj_4220, n42360, n17509, n17497, n13_adj_4221, 
        n43446, n17396, n42299, n20, n29, n42883, n42085, n38228, 
        n19_adj_4222, n44218, n20_adj_4223, n34549, n19_adj_4224, 
        n46604, n49937, n34548, n34547, n17_adj_4225, n16_adj_4226, 
        n49940, n8_adj_4227, n42248, n44282, n30_adj_4228, n25_adj_4229, 
        n19_adj_4230, n46590, n49931, tx_transmit_N_2998, n34584, 
        n34583, n18138;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    
    wire n18137, n34582, n18136, n34581, n34580, n17_adj_4231, n16_adj_4232, 
        n49934, n17964, n34577, n3735, n6_adj_4233, n17672, n19_adj_4234, 
        n46589, n49925, n17_adj_4235, n16_adj_4236, n49928, n16676, 
        n42487, n18413, n42058, n1716, n42305, n6_adj_4237, n3_adj_4238, 
        n6_adj_4239, n42274, n42035, n42092, n42146, n42094, n6_adj_4240, 
        n4_adj_4241, n6_adj_4242, n6_adj_4243, n6_adj_4244, n42283, 
        n1287, n42339, n37473, n28_adj_4245, n42049, n42203, n3761, 
        n16_adj_4246, n17_adj_4247, n16541, n16476, n16_adj_4248, 
        n17_adj_4249, n63, n16538, n18_adj_4250, n37409, n42302, 
        n42091, n20_adj_4251, n15_adj_4252, n63_adj_4253, n42155, 
        n17116, n42, n40, n41, n39, n38, n37_c, n48, n43, 
        n46588, n5_adj_4254, n49913, n4_adj_4255, n41704, n46678, 
        n888, n10_adj_4256, n16611, n14_adj_4257, n15_adj_4258, n10_adj_4259, 
        n14_adj_4260, n41833, n20_adj_4261, n19_adj_4262, n44308, 
        n63_adj_4263, n16558, n16677, n10_adj_4264, n16684, n17103, 
        Kp_23__N_1210, n42222, n42375, n12, n42438, n38274, n10_adj_4268, 
        n41913, n38259, n6_adj_4269, n42128, n31_adj_4270, n42381, 
        n17126, n6_adj_4271, n16253, n6_adj_4272, n6_adj_4273, n42414, 
        n6_adj_4274, n41983, n37982, n16310, n42072, n42289, n42235, 
        Kp_23__N_1136, n8_adj_4275, n7_adj_4276, n42268, n41941, n42405, 
        n42411, n16_adj_4278, n15_adj_4279, n42023, n17_adj_4280, 
        n38283;
    wire [31:0]n93;
    
    wire n17421, n12_adj_4281, n10_adj_4282, n42100, n14_adj_4283, 
        n59, n42462, n6_adj_4284, n42399, n17145, n42232, n17535, 
        n4_adj_4285, n4_adj_4286, n141, n10_adj_4287, n42131, n42016, 
        n28_adj_4288, n26_adj_4289, n27_adj_4290, n41968, n25_adj_4291, 
        n44019, n42435, n38_adj_4292, n42286, n36, n37_adj_4293, 
        n40_adj_4294, n35, n44, n39_adj_4295, n10_adj_4296, n16_adj_4297, 
        n12_adj_4298, n42444, Kp_23__N_588, n10_adj_4299, n42200, 
        n38325, n10_adj_4300, n42121, n42296, n13_adj_4304, n42213, 
        n8_adj_4305, n7_adj_4306, n10_adj_4307, n41888, n42311, n14_adj_4308, 
        n16521, n9, n47, n42396, n13980, n25891, n25307, n6_adj_4309, 
        n42134, n42336, n14_adj_4310, n10_adj_4311, n42327, n42116, 
        n12_adj_4312, n41910, n10_adj_4313, n16_adj_4314, n17_adj_4315, 
        n46582, n19_adj_4316, n16_adj_4317, n17_adj_4318, n46583, 
        n19_adj_4319, n16_adj_4320, n17_adj_4321, n46584, n19_adj_4322, 
        n16_adj_4323, n17_adj_4324, n46585, n19_adj_4325, tx_active;
    wire [2:0]r_SM_Main_c;   // verilog/uart_tx.v(31[16:25])
    
    wire n10142, n4_adj_4326, n41424, n4_adj_4327, n26_adj_4328;
    wire [31:0]\FRAME_MATCHER.state_31__N_2275 ;
    
    wire n4_adj_4329, n49916, n16679, n16772, n6_adj_4331, n42450, 
        n10_adj_4332, n37697, n41965, n42280, n47196, n5_adj_4333, 
        n44375, n49874, n49838, n49826, n16994, n42456, n47191, 
        n5_adj_4334, n44372, n49880, n49850, n49844, n42241, n47184, 
        n5_adj_4335, n44369, n49886, n49856, n42039, n49820, n48582, 
        n48586, n42210, n49892, n46613, n6_adj_4336, n5_adj_4337, 
        n44366, n17004, n6_adj_4338, n41971, n6_adj_4339, n46610, 
        n6_adj_4340, n5_adj_4341, n44363, n42225, n47168, n5_adj_4342, 
        n44360, n41952, n34, n39_adj_4344, n42109, n42314, n42292, 
        n42271, n42366, n42019, n16_adj_4345, n17304, n17301, n4_adj_4346, 
        n26152, n2_adj_4347, n44320, n42664, n26156, n49889, n7_adj_4348, 
        n16938, n42784, n5_adj_4349, n6_adj_4350;
    wire [31:0]\FRAME_MATCHER.state_31__N_2243 ;
    
    wire n37905, n6_adj_4351, n42265, n42441, n42137, n22_adj_4352, 
        n42387, n20_adj_4353, n42465, n24_adj_4354, n42207, n16249, 
        n42420, n42426, n10_adj_4355, n42321, n16691, n42402, n10_adj_4356, 
        n42423, n10_adj_4357, n42173, n17424, n42363, n41885, n16_adj_4358, 
        n42046, n17_adj_4359, n1185, n42029, n20_adj_4360, n41980, 
        n19_adj_4361, n17430, n21, n42026, n1515, n6_adj_4363, n37540, 
        n37514, n10_adj_4364, n14_adj_4365, n16815, n42277, n37471, 
        n42009, n26_adj_4366, n42197, n16989, n41986, n29_adj_4367, 
        n28_adj_4368, n32, n42161, n27_adj_4369, n28_adj_4370, n35_adj_4371, 
        n42194, n40_adj_4372, n42182, n38_adj_4373, n42164, n37_adj_4374, 
        n17289, n42378, n43449, n10_adj_4375, n38252, n42191, n11, 
        n13_adj_4376, n17138, n42317, n16768, n42354, n6_adj_4377, 
        n12_adj_4378, n8_adj_4379, n17375, n38226, n7_adj_4380, n42259, 
        n43760, n16862, n6_adj_4381, n16873, n42052, n17142, n37575, 
        n42176, n42185, n1379, n42055, n42112, n41895, n17198, 
        n42417, n10_adj_4382, n43751, n42324, n42453, n41919, n41929, 
        n41974, n41938, n30_adj_4383, n16778, n34_adj_4384, n32_adj_4385, 
        n36_adj_4386, n42032, n31_adj_4387, n18_adj_4388, n24_adj_4389, 
        n22_adj_4390, n26_adj_4391, n17206, n10_adj_4392, n41946, 
        n14_adj_4393, n37877, n18_adj_4394, n24_adj_4395, n22_adj_4396, 
        n26_adj_4397, n12_adj_4398, n10_adj_4399, n14_adj_4400, n49883, 
        n12_adj_4401, n49877, n49871, n10_adj_4402, n49859, n49853, 
        n49847, n49841, n42103, n49835, n16_adj_4404, n22_adj_4405, 
        n49823, n20_adj_4406, n24_adj_4408, n49817, n10_adj_4409, 
        n14_adj_4410, n13_adj_4411, n22_adj_4412, n27_adj_4413, n26_adj_4414, 
        n44231, n44302, n31_adj_4415;
    
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n23171));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18460));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18459));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18458));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18457));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_24 (.CI(n34575), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n34576));
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18456));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18455));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18454));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18453));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18452));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18451));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18450));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18449));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_23_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n34574), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_4113), .S(n3_c));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n18448));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_23 (.CI(n34574), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n34575));
    SB_LUT4 i13054_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n18338));
    defparam i13054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n18447));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18418));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n18379));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18378));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18377));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18376));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18337));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18375));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18374));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18373));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18336));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18335));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18334));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_27 (.CI(n34578), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n34579));
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18333));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18332));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n18331));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n18330));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_22_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n34573), .O(n2_adj_4114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n18329));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n18328));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18372));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n18327));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_22 (.CI(n34573), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n34574));
    SB_LUT4 add_44_21_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n34572), .O(n2_adj_4115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n18326));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n18325));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18371));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n18324));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n18323));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18370));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18369));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n18667));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n18666));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n18665));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n18664));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n18663));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n18662));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n18661));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n18660));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n18659));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n18658));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n18657));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n18656));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n18655));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n18654));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n18653));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n18652));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n18651));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n18650));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n18649));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n18648));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n18647));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n18646));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n18645));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13055_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n18339));
    defparam i13055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18368));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18367));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18366));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18365));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n18593));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18364));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18363));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18362));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18361));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18360));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18359));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18358));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13056_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n18340));
    defparam i13056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n23932));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18356));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18355));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18354));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter_c[1]), .C(clk32MHz), 
            .E(VCC_net), .D(n18550));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter_c[2]), .C(clk32MHz), 
            .E(VCC_net), .D(n18547));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), .C(clk32MHz), 
            .E(VCC_net), .D(n18544));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), .C(clk32MHz), 
            .E(VCC_net), .D(n18541));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), .C(clk32MHz), 
            .E(VCC_net), .D(n18538));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
            .E(VCC_net), .D(n18535));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
            .E(VCC_net), .D(n18509));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n50009));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18353));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18352));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18471));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18470));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18469));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18468));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18467));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18466));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n23694));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18464));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18463));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18462));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n18322));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n18321));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n18320));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n18319));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n18318));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n18317));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n18316));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n18315));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18411));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18410));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18409));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18408));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18407));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18406));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18405));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n18314));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n18313));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n18312));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n18311));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n18310));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n18309));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n18308));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n18307));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n18306));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n18305));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18404));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n18304));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n18303));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n18302));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n18301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n18300));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n18299));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18403));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18402));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18401));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18400));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18399));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13057_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n18341));
    defparam i13057_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13058_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n18342));
    defparam i13058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13059_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n18343));
    defparam i13059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13060_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n18344));
    defparam i13060_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13061_3_lut_4_lut (.I0(n8), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n18345));
    defparam i13061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18398));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18397));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13135_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18419));
    defparam i13135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18351));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13136_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18420));
    defparam i13136_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18350));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13137_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18421));
    defparam i13137_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18348));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18347));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13138_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18422));
    defparam i13138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18346));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n18298));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18417));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_21 (.CI(n34572), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n34573));
    SB_LUT4 add_44_20_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n34571), .O(n2_adj_4117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_20 (.CI(n34571), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n34572));
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n18297));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13139_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18423));
    defparam i13139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18345));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13140_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18424));
    defparam i13140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18396));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n18446));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n18445));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18344));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n18444));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13141_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18425));
    defparam i13141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_19_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n34570), .O(n2_adj_4118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13134_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41861), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18418));
    defparam i13134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_19 (.CI(n34570), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n34571));
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n18296));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4119), .S(n3_adj_4120));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_18_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n34569), .O(n2_adj_4121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_18 (.CI(n34569), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n34570));
    SB_LUT4 add_44_17_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n34568), .O(n2_adj_4122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 equal_75_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4123));   // verilog/coms.v(154[7:23])
    defparam equal_75_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4116));   // verilog/coms.v(154[7:23])
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n18443));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n18295));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_17 (.CI(n34568), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n34569));
    SB_LUT4 add_44_16_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n34567), .O(n2_adj_4124)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_16 (.CI(n34567), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n34568));
    SB_LUT4 add_44_15_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n34566), .O(n2_adj_4125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_15 (.CI(n34566), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n34567));
    SB_LUT4 i5_3_lut (.I0(\FRAME_MATCHER.state [9]), .I1(n10), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n41876));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_44_14_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n34565), .O(n2_adj_4126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_14 (.CI(n34565), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n34566));
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n16608), .I3(\FRAME_MATCHER.i [4]), .O(n16468));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13155_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n18439));
    defparam i13155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n18442));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [4]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n41874));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18412));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n18294));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n18293));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n18292));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n18291));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n18290));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_13_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n34564), .O(n2_adj_4128)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_13 (.CI(n34564), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n34565));
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n18289));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_12_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n34563), .O(n2_adj_4129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n18288));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n18287));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_887 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n25285), .O(n41861));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_887.LUT_INIT = 16'hefff;
    SB_LUT4 i36424_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n16446), .I2(GND_net), 
            .I3(GND_net), .O(n44325));
    defparam i36424_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16682));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20352_1_lut (.I0(n25611), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1774));
    defparam i20352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44377), .I3(n44376), 
            .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44374), .I3(n44373), 
            .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44371), .I3(n44370), 
            .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i20040_2_lut (.I0(n31), .I1(n25297), .I2(GND_net), .I3(GND_net), 
            .O(n25299));
    defparam i20040_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_888 (.I0(\data_in_frame[5] [5]), .I1(n41996), .I2(n41891), 
            .I3(\data_in_frame[1] [3]), .O(n16804));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_CARRY add_44_12 (.CI(n34563), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n34564));
    SB_LUT4 i2_3_lut_adj_889 (.I0(\data_in_frame[4] [5]), .I1(n5_c), .I2(n4_c), 
            .I3(GND_net), .O(n17168));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_889.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_890 (.I0(\data_in_frame[1] [6]), .I1(n41993), .I2(\data_in_frame[4] [2]), 
            .I3(GND_net), .O(n16893));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_890.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n41996));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_in_frame[3] [3]), .I1(n41977), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44368), .I3(n49964), 
            .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i4_4_lut (.I0(n16307), .I1(n6_adj_4130), .I2(\data_in_frame[3] [0]), 
            .I3(n6_c), .O(Kp_23__N_679));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1187_i16_2_lut (.I0(Kp_23__N_679), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/coms.v(230[9:81])
    defparam equal_1187_i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_893 (.I0(Kp_23__N_809), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17503));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_894 (.I0(n4_adj_4131), .I1(n42229), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n17035));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_895 (.I0(\data_in_frame[4] [3]), .I1(n41898), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[2] [1]), .O(n16898));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_896 (.I0(n42262), .I1(\data_in_frame[0] [7]), .I2(n42384), 
            .I3(GND_net), .O(n42229));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_896.LUT_INIT = 16'h9696;
    SB_LUT4 add_44_11_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n34562), .O(n2_adj_4132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_11 (.CI(n34562), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n34563));
    SB_LUT4 i4_4_lut_adj_897 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[3] [2]), .I3(n6_adj_4133), .O(n41977));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n41898));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16827));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_900 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n6_adj_4130));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_900.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [24]), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/coms.v(206[5:16])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_901 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_c));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_901.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44359), .I3(n44358), 
            .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44362), .I3(n49976), 
            .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\data_in_frame[1] [3]), .I1(n41999), .I2(n41925), 
            .I3(n16827), .O(n42262));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_903 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n41993));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_904 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [5]), .I3(n42262), .O(n42384));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_905 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n15066));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_905.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(Kp_23__N_676), .I1(n42384), .I2(n41993), .I3(\data_in_frame[0] [3]), 
            .O(n16_adj_4134));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[1] [5]), .I1(n41898), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[2] [3]), .O(n17));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in_frame[2] [6]), .I2(n16_adj_4134), 
            .I3(\data_in_frame[0] [6]), .O(n16307));   // verilog/coms.v(76[16:27])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44365), .I3(n49970), 
            .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_adj_906 (.I0(n16307), .I1(n15066), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4135));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_10_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n34561), .O(n2_adj_4136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_10 (.CI(n34561), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n34562));
    SB_LUT4 i4_4_lut_adj_907 (.I0(n41977), .I1(n41891), .I2(\data_in_frame[1] [2]), 
            .I3(n6_adj_4135), .O(n41956));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n17037), .I1(n41956), .I2(GND_net), 
            .I3(GND_net), .O(n37571));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_909 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[2] [6]), .O(n43394));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_910 (.I0(\data_in_frame[0] [7]), .I1(n43394), .I2(\data_in_frame[3] [0]), 
            .I3(\data_in_frame[1] [0]), .O(n17037));
    defparam i3_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_911 (.I0(\data_in_frame[5] [2]), .I1(n17037), .I2(\data_in_frame[3] [1]), 
            .I3(GND_net), .O(n37696));
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i13098_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18382));
    defparam i13098_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_912 (.I0(n42229), .I1(n41956), .I2(\data_in_frame[5] [1]), 
            .I3(GND_net), .O(n37621));
    defparam i2_3_lut_adj_912.LUT_INIT = 16'h9696;
    SB_LUT4 equal_1187_i15_2_lut (.I0(Kp_23__N_676), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // verilog/coms.v(230[9:81])
    defparam equal_1187_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13099_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18383));
    defparam i13099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n41999));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 equal_1187_i8_2_lut (.I0(Kp_23__N_729), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4138));   // verilog/coms.v(230[9:81])
    defparam equal_1187_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_914 (.I0(\data_in_frame[3] [6]), .I1(n41999), .I2(\data_in_frame[3] [7]), 
            .I3(\data_in_frame[4] [0]), .O(n16851));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_9_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n34560), .O(n2_adj_4139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_915 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [4]), 
            .I2(n4_c), .I3(n41898), .O(n16903));   // verilog/coms.v(166[9:87])
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_CARRY add_44_9 (.CI(n34560), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n34561));
    SB_LUT4 i12_4_lut (.I0(n15_c), .I1(n37621), .I2(n1), .I3(n37696), 
            .O(n28_c));
    defparam i12_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut (.I0(n16903), .I1(n16889), .I2(n16851), .I3(n8_adj_4138), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n16893), .I1(n17185), .I2(n17168), .I3(n16804), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_916 (.I0(n16898), .I1(n17035), .I2(n17503), .I3(n16), 
            .O(n25));
    defparam i9_4_lut_adj_916.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28_c), .O(n31));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_917 (.I0(n7_c), .I1(n41876), .I2(n144), .I3(n41874), 
            .O(n26154));
    defparam i4_4_lut_adj_917.LUT_INIT = 16'hfffe;
    SB_LUT4 i20370_4_lut (.I0(n25297), .I1(n31_adj_4140), .I2(n31), .I3(\FRAME_MATCHER.state [1]), 
            .O(n25630));
    defparam i20370_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_3_lut (.I0(n25630), .I1(n13947), .I2(n26154), .I3(GND_net), 
            .O(n43448));
    defparam i3_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i13100_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18384));
    defparam i13100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13096_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[14]_c [2]), .O(n18380));
    defparam i13096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_8_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n34559), .O(n2_adj_4141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_8 (.CI(n34559), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n34560));
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n18286));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_7_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n34558), .O(n2_adj_4142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n18285));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13101_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[14]_c [7]), .O(n18385));
    defparam i13101_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_7 (.CI(n34558), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n34559));
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n18284));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13097_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[3]), 
            .I3(\data_in_frame[14]_c [3]), .O(n18381));
    defparam i13097_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13094_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18378));
    defparam i13094_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13095_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n18379));
    defparam i13095_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n18283));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n18282));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18441));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_6_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n34557), .O(n2_adj_4143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18440));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18439));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n18281));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_6 (.CI(n34557), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n34558));
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n18280));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10_4_lut_adj_918 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [19]), 
            .O(n24));   // verilog/coms.v(206[5:16])
    defparam i10_4_lut_adj_918.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n18279));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n18278));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_919 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n25285), .O(n41843));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_919.LUT_INIT = 16'hfeff;
    SB_LUT4 add_44_5_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n34556), .O(n2_adj_4144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n18277));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n18276));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n18275));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n18274));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n18273));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n18272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n18271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n18270));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n18269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n18268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n18267));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n18266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n18265));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n18264));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n18263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n18262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n18261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n18260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n18259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n18258));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n18257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n18256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n18255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n18254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n18253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n18252));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_920 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n25285), .O(n41852));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_920.LUT_INIT = 16'hefff;
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n18251));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n18250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n18249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n18248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n18247));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n18246));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_5 (.CI(n34556), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n34557));
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n18245));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4144), .S(n3_adj_4145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n18244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n18243));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_4_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n34555), .O(n2_adj_4119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n18242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n18241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n18240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n18239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n18238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n18237));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n18236));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n18235));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n18234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n18233));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n18232));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n18231));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_4 (.CI(n34555), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n34556));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n41843), .I3(\FRAME_MATCHER.i [0]), .O(n41851));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18416));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_71_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4137));
    defparam equal_71_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 add_44_3_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n34554), .O(n2_adj_4146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(\FRAME_MATCHER.state [17]), 
            .O(n22));   // verilog/coms.v(206[5:16])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18438));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n18230));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20162_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n16468), .I3(\FRAME_MATCHER.i [31]), .O(n2857));
    defparam i20162_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i1981_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_4147));
    defparam i1981_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_921 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n41852), .I3(\FRAME_MATCHER.i [0]), .O(n41860));
    defparam i1_2_lut_3_lut_4_lut_adj_921.LUT_INIT = 16'hf7ff;
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18437));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n18229));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13086_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n18370));
    defparam i13086_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n18228));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18395));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18436));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4143), .S(n3_adj_4148));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13087_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n18371));
    defparam i13087_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4142), .S(n3_adj_4149));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4141), .S(n3_adj_4150));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4139), .S(n3_adj_4151));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4136), .S(n3_adj_4152));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4132), .S(n3_adj_4153));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4129), .S(n3_adj_4154));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4128), .S(n3_adj_4155));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4126), .S(n3_adj_4156));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4125), .S(n3_adj_4157));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4124), .S(n3_adj_4158));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4122), .S(n3_adj_4159));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4121), .S(n3_adj_4160));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4118), .S(n3_adj_4161));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4117), .S(n3_adj_4162));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4115), .S(n3_adj_4163));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4114), .S(n3_adj_4164));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_4165));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4166), .S(n3_adj_4167));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4168), .S(n3_adj_4169));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4170), .S(n3_adj_4171));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4172), .S(n3_adj_4173));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4174), .S(n3_adj_4175));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4176), .S(n3_adj_4177));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4178), .S(n3_adj_4179));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4180), .S(n3_adj_4181));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4182), .S(n3_adj_4183));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4184), .S(n3_adj_4185));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n17676), .D(n43355));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n17676), .D(n43374));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n17676), .D(n43377));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n17676), .D(n44061));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n17676), .D(n43198));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n17676), .D(n44072));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n17676), .D(n43875));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n17676), .D(n43169));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n17676), .D(n43711));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n17676), .D(n42290));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n17676), .D(n42412));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n17676), .D(n43317));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n17676), .D(n43126));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n17676), .D(n42174));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n17676), .D(n43726));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n17676), .D(n43199));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n18227));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n18226));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n18225));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n18224));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n18223));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n18222));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n18221));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n18220));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n18219));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n18218));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n18217));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n18216));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n18215));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n40980), .S(n50161));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n40984), .S(n41172));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n41264), .S(n40986));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n41266), .S(n41046));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n41268), .S(n41044));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n41270), .S(n41042));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n41282), .S(n41052));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n41334), .S(n41060));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n41342), .S(n40966));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n41344), .S(n41050));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n41346), .S(n41040));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n7_adj_4186), .S(n8_adj_4187));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n7_adj_4188), .S(n8_adj_4189));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_4190), .S(n8_adj_4191));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n41240), .S(n40988));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n7_adj_4192), .S(n8_adj_4193));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n41242), .S(n41038));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n41244), .S(n41036));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n41246), .S(n41034));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n25288), .S(n41032));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n41248), .S(n41030));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_4194), .S(n25290));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n41250), .S(n41028));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n41252), .S(n41026));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n7_adj_4195), .S(n8_adj_4196));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_4197), .S(n8_adj_4198));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n7_adj_4199), .S(n8_adj_4200));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n41254), .S(n40982));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n41144), .S(n40964));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4201), .S(n8_adj_4202));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n18214));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13088_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n18372));
    defparam i13088_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_922 (.I0(\FRAME_MATCHER.state [29]), .I1(n24), 
            .I2(n18), .I3(\FRAME_MATCHER.state [30]), .O(n26_adj_4203));   // verilog/coms.v(206[5:16])
    defparam i12_4_lut_adj_922.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n18213));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n18212));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i11_3_lut (.I0(\FRAME_MATCHER.state [21]), .I1(n22), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n25_adj_4204));   // verilog/coms.v(206[5:16])
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n18211));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n18210));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n18209));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n18208));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n18207));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n18206));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n18205));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n18204));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n18203));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut (.I0(\FRAME_MATCHER.state [28]), .I1(n25_adj_4204), 
            .I2(\FRAME_MATCHER.state [26]), .I3(n26_adj_4203), .O(n7_c));   // verilog/coms.v(206[5:16])
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_923 (.I0(n7_c), .I1(n41874), .I2(n41876), .I3(n144), 
            .O(n16446));   // verilog/coms.v(206[5:16])
    defparam i4_4_lut_adj_923.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\FRAME_MATCHER.state [1]), .I1(n16446), 
            .I2(GND_net), .I3(GND_net), .O(n16563));   // verilog/coms.v(195[5:24])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_925 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_c));
    defparam i6_4_lut_adj_925.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_926 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_4205));   // verilog/coms.v(232[13:35])
    defparam i6_4_lut_adj_926.LUT_INIT = 16'hfffe;
    SB_LUT4 i13089_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n18373));
    defparam i13089_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13090_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n18374));
    defparam i13090_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_c));
    defparam i5_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_927 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_4206));   // verilog/coms.v(232[13:35])
    defparam i5_4_lut_adj_927.LUT_INIT = 16'hfffe;
    SB_LUT4 i20038_4_lut (.I0(n13_adj_4206), .I1(n13_c), .I2(n14_adj_4205), 
            .I3(n14_c), .O(n25297));
    defparam i20038_4_lut.LUT_INIT = 16'h32fa;
    SB_LUT4 i13091_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n18375));
    defparam i13091_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_928 (.I0(n42251), .I1(n17415), .I2(\data_in_frame[21] [6]), 
            .I3(n42393), .O(n10_adj_4207));   // verilog/coms.v(71[16:42])
    defparam i4_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_929 (.I0(n41962), .I1(n10_adj_4207), .I2(n16971), 
            .I3(GND_net), .O(n43667));   // verilog/coms.v(71[16:42])
    defparam i5_3_lut_adj_929.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_930 (.I0(n43329), .I1(n38220), .I2(\data_in_frame[16] [7]), 
            .I3(\data_in_frame[18] [5]), .O(n18_adj_4208));
    defparam i7_4_lut_adj_930.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_c));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4209));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'ha300;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4210));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36477_4_lut (.I0(n19_c), .I1(\data_out_frame[22] [0]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n44379));
    defparam i36477_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[20] [5]), .I3(n18_adj_4211), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i36478_3_lut (.I0(n49952), .I1(n44379), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44380));
    defparam i36478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36455_3_lut (.I0(n5_adj_4210), .I1(n6_adj_4209), .I2(n45195), 
            .I3(GND_net), .O(n44357));
    defparam i36455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_931 (.I0(\data_in_frame[7] [1]), .I1(n17325), 
            .I2(n37571), .I3(n42408), .O(n28_adj_4212));
    defparam i11_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i36457_4_lut (.I0(n44357), .I1(n44380), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44359));
    defparam i36457_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36456_3_lut (.I0(n49946), .I1(n49862), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44358));
    defparam i36456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13093_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n18377));
    defparam i13093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17279_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41852), .I2(\data_in_frame[13] [6]), 
            .I3(rx_data[6]), .O(n18376));
    defparam i17279_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i10_4_lut_adj_932 (.I0(n42372), .I1(n42447), .I2(\data_in_frame[15] [7]), 
            .I3(n42167), .O(n27_adj_4213));
    defparam i10_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_CARRY add_44_3 (.CI(n34554), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n34555));
    SB_LUT4 add_44_2_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n2_adj_4113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n18202));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n18201));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n34554));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_933 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n41861), .I3(\FRAME_MATCHER.i [0]), .O(n41862));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_933.LUT_INIT = 16'hfffb;
    SB_LUT4 add_639_9_lut (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4497), .I3(n34553), .O(n18507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_9_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n18200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n18199));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n18198));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n18197));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n18196));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n18195));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n18194));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n18193));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n18192));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n18191));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n18190));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n18189));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n18188));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n18187));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n18186));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n18185));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n18184));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n18183));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_639_8_lut (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[6]), 
            .I2(n4497), .I3(n34552), .O(n18533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_8_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n18182));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n18181));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n18180));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n18179));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n18178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n18177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n18176));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n18175));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n18174));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n18173));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n18172));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n18171));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n18170));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n18169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n18168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n18167));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_639_8 (.CI(n34552), .I0(byte_transmit_counter_c[6]), .I1(n4497), 
            .CO(n34553));
    SB_LUT4 add_639_7_lut (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[5]), 
            .I2(n4497), .I3(n34551), .O(n18536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_7_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n18166));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n18165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n18164));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3227 (.Q(r_SM_Main_2__N_3106[0]), .C(clk32MHz), 
            .D(n46769), .R(n42491));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n18163));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_934 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n41843), .I3(\FRAME_MATCHER.i [0]), .O(n41848));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_934.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_935 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n41852), .I3(\FRAME_MATCHER.i [0]), .O(n41857));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_935.LUT_INIT = 16'hfffb;
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n18162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n18161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n18160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n18159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n18158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n18157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n18156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n18155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18394));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18415));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n18154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n18153));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49985));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49985_bdd_4_lut (.I0(n49985), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49988));
    defparam n49985_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n18152));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n18151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n18150));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n18149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n18148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n18147));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n18146));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter_c[1]), 
            .I1(n44336), .I2(n44337), .I3(byte_transmit_counter_c[2]), 
            .O(n49973));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49973_bdd_4_lut (.I0(n49973), .I1(n44334), .I2(n44333), .I3(byte_transmit_counter_c[2]), 
            .O(n49976));
    defparam n49973_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42042 (.I0(byte_transmit_counter_c[1]), 
            .I1(n44342), .I2(n44343), .I3(byte_transmit_counter_c[2]), 
            .O(n49967));
    defparam byte_transmit_counter_1__bdd_4_lut_42042.LUT_INIT = 16'he4aa;
    SB_LUT4 n49967_bdd_4_lut (.I0(n49967), .I1(n44340), .I2(n44339), .I3(byte_transmit_counter_c[2]), 
            .O(n49970));
    defparam n49967_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42037 (.I0(byte_transmit_counter_c[1]), 
            .I1(n44348), .I2(n44349), .I3(byte_transmit_counter_c[2]), 
            .O(n49961));
    defparam byte_transmit_counter_1__bdd_4_lut_42037.LUT_INIT = 16'he4aa;
    SB_LUT4 n49961_bdd_4_lut (.I0(n49961), .I1(n44346), .I2(n44345), .I3(byte_transmit_counter_c[2]), 
            .O(n49964));
    defparam n49961_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_42051 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49955));
    defparam byte_transmit_counter_0__bdd_4_lut_42051.LUT_INIT = 16'he4aa;
    SB_LUT4 n49955_bdd_4_lut (.I0(n49955), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n49958));
    defparam n49955_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_42027 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49949));
    defparam byte_transmit_counter_0__bdd_4_lut_42027.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18342));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n18145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n18144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n18143));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18341));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18340));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18393));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_936 (.I0(n42097), .I1(n16750), .I2(\data_in_frame[20] [2]), 
            .I3(n42308), .O(n10_adj_4214));
    defparam i4_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18392));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18339));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[21] [1]), .I1(n16268), .I2(n38270), 
            .I3(GND_net), .O(n42070));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18391));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49949_bdd_4_lut (.I0(n49949), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49952));
    defparam n49949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18390));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_639_7 (.CI(n34551), .I0(byte_transmit_counter_c[5]), .I1(n4497), 
            .CO(n34552));
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18414));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_639_6_lut (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[4]), 
            .I2(n4497), .I3(n34550), .O(n18539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_6_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14]_c [3]), .C(clk32MHz), 
           .D(n18381));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_42022 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49943));
    defparam byte_transmit_counter_0__bdd_4_lut_42022.LUT_INIT = 16'he4aa;
    SB_LUT4 equal_64_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4127));   // verilog/coms.v(154[7:23])
    defparam equal_64_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_CARRY add_639_6 (.CI(n34550), .I0(byte_transmit_counter_c[4]), .I1(n4497), 
            .CO(n34551));
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18389));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i0 (.Q(deadband[0]), .C(clk32MHz), .D(n17862));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18435));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_937 (.I0(n37561), .I1(n42345), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4215));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18434));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18433));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18432));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18431));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18430));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18429));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18428));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18427));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18426));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18425));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18424));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18423));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18422));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49943_bdd_4_lut (.I0(n49943), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49946));
    defparam n49943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_938 (.I0(\data_in_frame[20] [6]), .I1(n38230), 
            .I2(n42152), .I3(n6_adj_4215), .O(n43335));
    defparam i4_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_939 (.I0(n42179), .I1(\data_in_frame[20] [0]), 
            .I2(n43390), .I3(n42351), .O(n10_adj_4216));
    defparam i4_4_lut_adj_939.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_940 (.I0(\data_in_frame[20] [3]), .I1(n37587), 
            .I2(n42079), .I3(GND_net), .O(n8_adj_4217));
    defparam i3_3_lut_adj_940.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_941 (.I0(\data_in_frame[21] [2]), .I1(n42149), 
            .I2(\data_in_frame[19] [1]), .I3(n16268), .O(n43441));
    defparam i3_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_942 (.I0(Kp_23__N_1213), .I1(n10_adj_4216), .I2(n37485), 
            .I3(GND_net), .O(n43365));
    defparam i5_3_lut_adj_942.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_943 (.I0(\data_in_frame[18] [2]), .I1(n43441), 
            .I2(n8_adj_4217), .I3(n17325), .O(n22_adj_4218));
    defparam i6_4_lut_adj_943.LUT_INIT = 16'hb77b;
    SB_LUT4 i2_3_lut_adj_944 (.I0(n41959), .I1(n42245), .I2(\data_in_frame[21] [4]), 
            .I3(GND_net), .O(n42959));
    defparam i2_3_lut_adj_944.LUT_INIT = 16'h9696;
    SB_LUT4 i36383_4_lut (.I0(\data_in_frame[20] [1]), .I1(n43667), .I2(n42076), 
            .I3(\data_in_frame[19] [7]), .O(n44278));
    defparam i36383_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_4_lut_adj_945 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[19] [1]), 
            .I2(n16268), .I3(n42245), .O(n42825));
    defparam i2_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_946 (.I0(\data_in_frame[20] [4]), .I1(n22_adj_4218), 
            .I2(n43365), .I3(n42158), .O(n27_adj_4219));
    defparam i11_4_lut_adj_946.LUT_INIT = 16'hdfef;
    SB_LUT4 i6_4_lut_adj_947 (.I0(n42390), .I1(Kp_23__N_1201), .I2(n42188), 
            .I3(\data_in_frame[15] [4]), .O(n14_adj_4220));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_948 (.I0(\data_in_frame[21] [7]), .I1(n42360), 
            .I2(n17509), .I3(n17497), .O(n13_adj_4221));   // verilog/coms.v(71[16:42])
    defparam i5_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_949 (.I0(n16268), .I1(n42149), .I2(n38270), .I3(\data_in_frame[21] [0]), 
            .O(n43446));
    defparam i2_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_950 (.I0(n37512), .I1(n18_adj_4208), .I2(n17396), 
            .I3(n42299), .O(n20));
    defparam i9_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n27_adj_4213), .I1(n29), .I2(n28_adj_4212), 
            .I3(n30), .O(n42883));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_951 (.I0(n42085), .I1(\data_in_frame[20] [7]), 
            .I2(n38228), .I3(n38270), .O(n19_adj_4222));
    defparam i8_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i36329_3_lut (.I0(n43446), .I1(n13_adj_4221), .I2(n14_adj_4220), 
            .I3(GND_net), .O(n44218));
    defparam i36329_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i4_4_lut_adj_952 (.I0(n37587), .I1(n42070), .I2(n10_adj_4214), 
            .I3(n17415), .O(n20_adj_4223));
    defparam i4_4_lut_adj_952.LUT_INIT = 16'hedde;
    SB_LUT4 add_639_5_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[3]), 
            .I2(n4497), .I3(n34549), .O(n18542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42032 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4224), .I2(n46604), .I3(byte_transmit_counter_c[2]), 
            .O(n49937));
    defparam byte_transmit_counter_1__bdd_4_lut_42032.LUT_INIT = 16'he4aa;
    SB_CARRY add_639_5 (.CI(n34549), .I0(byte_transmit_counter_c[3]), .I1(n4497), 
            .CO(n34550));
    SB_LUT4 add_639_4_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[2]), 
            .I2(n4497), .I3(n34548), .O(n18545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_639_4 (.CI(n34548), .I0(byte_transmit_counter_c[2]), .I1(n4497), 
            .CO(n34549));
    SB_LUT4 add_639_3_lut (.I0(byte_transmit_counter_c[1]), .I1(byte_transmit_counter_c[1]), 
            .I2(n4497), .I3(n34547), .O(n18548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 n49937_bdd_4_lut (.I0(n49937), .I1(n17_adj_4225), .I2(n16_adj_4226), 
            .I3(byte_transmit_counter_c[2]), .O(n49940));
    defparam n49937_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13046_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n18330));
    defparam i13046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_639_3 (.CI(n34547), .I0(byte_transmit_counter_c[1]), .I1(n4497), 
            .CO(n34548));
    SB_LUT4 i36386_4_lut (.I0(n41959), .I1(n43335), .I2(n42248), .I3(\data_in_frame[21] [5]), 
            .O(n44282));
    defparam i36386_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i14_4_lut (.I0(n27_adj_4219), .I1(n42825), .I2(n44278), .I3(n42959), 
            .O(n30_adj_4228));
    defparam i14_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i9_4_lut_adj_953 (.I0(n44218), .I1(n19_adj_4222), .I2(n42883), 
            .I3(n20), .O(n25_adj_4229));
    defparam i9_4_lut_adj_953.LUT_INIT = 16'h7fdf;
    SB_LUT4 i15_4_lut_adj_954 (.I0(n25_adj_4229), .I1(n30_adj_4228), .I2(n44282), 
            .I3(n20_adj_4223), .O(n31_adj_4140));
    defparam i15_4_lut_adj_954.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42012 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4230), .I2(n46590), .I3(byte_transmit_counter_c[2]), 
            .O(n49931));
    defparam byte_transmit_counter_1__bdd_4_lut_42012.LUT_INIT = 16'he4aa;
    SB_LUT4 add_639_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_2998), .I3(GND_net), .O(n2244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13047_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n18331));
    defparam i13047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_639_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2998), 
            .CO(n34547));
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n18142));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13048_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18332));
    defparam i13048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n18141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18388));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13049_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18333));
    defparam i13049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18387));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18386));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14]_c [7]), .C(clk32MHz), 
           .D(n18385));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n18140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n18139));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_33_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n34584), .O(n2_adj_4184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_32_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n34583), .O(n2_adj_4182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_32 (.CI(n34583), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n34584));
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18421));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0] [4]), .C(clk32MHz), 
           .D(n18138));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0] [3]), .C(clk32MHz), 
           .D(n18137));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_31_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n34582), .O(n2_adj_4180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_31 (.CI(n34582), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n34583));
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0] [2]), .C(clk32MHz), 
           .D(n18136));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n18135));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n18134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n18133));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n18132));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n18131));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n18130));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n18129));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n18128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n18127));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n18126));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_30_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n34581), .O(n2_adj_4178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_30 (.CI(n34581), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n34582));
    SB_LUT4 add_44_29_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n34580), .O(n2_adj_4176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_29 (.CI(n34580), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n34581));
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n18125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n18124));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n18123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n18122));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49931_bdd_4_lut (.I0(n49931), .I1(n17_adj_4231), .I2(n16_adj_4232), 
            .I3(byte_transmit_counter_c[2]), .O(n49934));
    defparam n49931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n18121));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n18120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n18119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n18118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n18117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n18116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n18115));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n18114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n18113));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n18112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n18111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n18110));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_28_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n34579), .O(n2_adj_4174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_28 (.CI(n34579), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n34580));
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n18109));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n18108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n18107));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12990_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n18274));
    defparam i12990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12991_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n18275));
    defparam i12991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12992_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n18276));
    defparam i12992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n18106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n18105));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n18104));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12993_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n18277));
    defparam i12993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12994_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n18278));
    defparam i12994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12995_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n18279));
    defparam i12995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n18103));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13050_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18334));
    defparam i13050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12996_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n18280));
    defparam i12996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n18102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n18101));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12997_3_lut_4_lut (.I0(n8), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n18281));
    defparam i12997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n18100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n18099));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n18098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n18097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n18096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14]_c [2]), .C(clk32MHz), 
           .D(n18380));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18384));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n18095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n18094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n18093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n18092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n18091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n18090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n18089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n18088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n18087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n18086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n18085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n18084));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n18083));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n18082));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i7 (.Q(\Kd[7] ), .C(clk32MHz), .D(n18081));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i6 (.Q(\Kd[6] ), .C(clk32MHz), .D(n18080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i5 (.Q(\Kd[5] ), .C(clk32MHz), .D(n18079));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12680_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n17964));
    defparam i12680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kd_i4 (.Q(\Kd[4] ), .C(clk32MHz), .D(n18078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i3 (.Q(\Kd[3] ), .C(clk32MHz), .D(n18077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i2 (.Q(\Kd[2] ), .C(clk32MHz), .D(n18076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i1 (.Q(\Kd[1] ), .C(clk32MHz), .D(n18075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n18074));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12983_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n18267));
    defparam i12983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12984_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n18268));
    defparam i12984_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n18073));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n18072));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n18071));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n18070));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n18069));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n18068));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n18067));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n18066));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n18065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n18064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n18063));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n18062));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n18061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n18060));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18338));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n18059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n18058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n18057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n18056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n18055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n18054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n18053));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n18052));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12985_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n18269));
    defparam i12985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n18051));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n18050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n18049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n18048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n18047));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n18046));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n18045));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n18044));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n18043));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n18042));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_26_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n34577), .O(n2_adj_4170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n18041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n18040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n18039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n18038));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12986_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n18270));
    defparam i12986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i1 (.Q(deadband[1]), .C(clk32MHz), .D(n18013));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12987_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n18271));
    defparam i12987_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12988_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n18272));
    defparam i12988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12989_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n18273));
    defparam i12989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i2 (.Q(deadband[2]), .C(clk32MHz), .D(n18012));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i3 (.Q(deadband[3]), .C(clk32MHz), .D(n18011));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i4 (.Q(deadband[4]), .C(clk32MHz), .D(n18010));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i5 (.Q(deadband[5]), .C(clk32MHz), .D(n18009));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i6 (.Q(deadband[6]), .C(clk32MHz), .D(n18008));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i7 (.Q(deadband[7]), .C(clk32MHz), .D(n18007));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i8 (.Q(deadband[8]), .C(clk32MHz), .D(n18006));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i9 (.Q(deadband[9]), .C(clk32MHz), .D(n18005));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i10 (.Q(deadband[10]), .C(clk32MHz), .D(n18004));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i11 (.Q(deadband[11]), .C(clk32MHz), .D(n18003));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i12 (.Q(deadband[12]), .C(clk32MHz), .D(n18002));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i13 (.Q(deadband[13]), .C(clk32MHz), .D(n18001));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i14 (.Q(deadband[14]), .C(clk32MHz), .D(n18000));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i15 (.Q(deadband[15]), .C(clk32MHz), .D(n17999));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i16 (.Q(deadband[16]), .C(clk32MHz), .D(n17998));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i17 (.Q(deadband[17]), .C(clk32MHz), .D(n17997));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i18 (.Q(deadband[18]), .C(clk32MHz), .D(n17996));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i19 (.Q(deadband[19]), .C(clk32MHz), .D(n17995));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13051_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18335));
    defparam i13051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i20 (.Q(deadband[20]), .C(clk32MHz), .D(n17994));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i21 (.Q(deadband[21]), .C(clk32MHz), .D(n17993));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i22 (.Q(deadband[22]), .C(clk32MHz), .D(n17992));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i23 (.Q(deadband[23]), .C(clk32MHz), .D(n17991));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_955 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n3735), .I3(n6_adj_4233), .O(n17672));   // verilog/coms.v(110[11:16])
    defparam i2_3_lut_4_lut_adj_955.LUT_INIT = 16'he000;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17983));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42007 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4234), .I2(n46589), .I3(byte_transmit_counter_c[2]), 
            .O(n49925));
    defparam byte_transmit_counter_1__bdd_4_lut_42007.LUT_INIT = 16'he4aa;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n40968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n17963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n17962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i0 (.Q(\Kd[0] ), .C(clk32MHz), .D(n17961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n17960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n17958));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13156_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n18440));
    defparam i13156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49925_bdd_4_lut (.I0(n49925), .I1(n17_adj_4235), .I2(n16_adj_4236), 
            .I3(byte_transmit_counter_c[2]), .O(n49928));
    defparam n49925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_44_26 (.CI(n34577), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n34578));
    SB_LUT4 add_44_25_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n34576), .O(n2_adj_4168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_25 (.CI(n34576), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n34577));
    SB_LUT4 add_44_27_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n34578), .O(n2_adj_4172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13052_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18336));
    defparam i13052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_24_lut (.I0(n1774), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n34575), .O(n2_adj_4166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_DFFE LED_3230 (.Q(LED_c), .C(clk32MHz), .E(n42487), .D(n16676));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13053_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18337));
    defparam i13053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18413));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12854_3_lut_4_lut (.I0(n3735), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17672), .I3(\data_out_frame[0] [4]), .O(n18138));
    defparam i12854_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i12852_3_lut_4_lut (.I0(n3735), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17672), .I3(\data_out_frame[0] [2]), .O(n18136));
    defparam i12852_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i12853_3_lut_4_lut (.I0(n3735), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17672), .I3(\data_out_frame[0] [3]), .O(n18137));
    defparam i12853_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18383));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_76_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_76_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18382));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n42058), .I1(\data_out_frame[20] [6]), .I2(\data_out_frame[16] [4]), 
            .I3(n1716), .O(n42305));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18420));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_956 (.I0(n42058), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[16] [3]), 
            .O(n6_adj_4237));
    defparam i1_2_lut_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4146), .S(n3_adj_4238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18419));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[13] [5]), .I3(GND_net), .O(n6_adj_4239));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_957 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[14] [0]), .I3(GND_net), .O(n42274));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_957.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(\data_out_frame[18] [5]), .I1(n42035), 
            .I2(n42092), .I3(n42146), .O(n43374));
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_959 (.I0(\data_out_frame[18] [5]), .I1(n42035), 
            .I2(n42305), .I3(n42094), .O(n43199));
    defparam i2_3_lut_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 equal_77_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4227));   // verilog/coms.v(154[7:23])
    defparam equal_77_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_960 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n6_adj_4240));
    defparam i1_2_lut_3_lut_adj_960.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[9] [4]), 
            .I2(n4_adj_4241), .I3(\data_out_frame[7] [4]), .O(n6_adj_4242));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_961 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n6_adj_4243));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_962 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n6_adj_4244));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_962.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_963 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n42283));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_963.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_964 (.I0(\data_out_frame[8] [5]), .I1(n1287), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[11] [2]), .O(n42339));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i9_2_lut_3_lut (.I0(\data_out_frame[10] [2]), .I1(n37473), .I2(\data_out_frame[10] [1]), 
            .I3(GND_net), .O(n28_adj_4245));
    defparam i9_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_965 (.I0(\data_out_frame[10] [2]), .I1(n37473), 
            .I2(\data_out_frame[14] [6]), .I3(n42049), .O(n42203));
    defparam i2_3_lut_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i20169_4_lut (.I0(n10_adj_4147), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n16608), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i20169_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i6_4_lut_adj_966 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4246));
    defparam i6_4_lut_adj_966.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_967 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4247));
    defparam i7_4_lut_adj_967.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_968 (.I0(n17_adj_4247), .I1(\data_in[1] [6]), .I2(n16_adj_4246), 
            .I3(\data_in[3] [7]), .O(n16541));
    defparam i9_4_lut_adj_968.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_969 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n16476), .O(n16_adj_4248));
    defparam i6_4_lut_adj_969.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_970 (.I0(n16541), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4249));
    defparam i7_4_lut_adj_970.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_971 (.I0(n17_adj_4249), .I1(\data_in[3] [5]), .I2(n16_adj_4248), 
            .I3(\data_in[3] [3]), .O(n63));
    defparam i9_4_lut_adj_971.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_972 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n16538), .I3(\data_in[1] [0]), .O(n18_adj_4250));
    defparam i7_4_lut_adj_972.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_4_lut_adj_973 (.I0(\data_out_frame[17] [2]), .I1(n37409), 
            .I2(n42302), .I3(n42091), .O(n43198));
    defparam i2_3_lut_4_lut_adj_973.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_974 (.I0(\data_in[1] [4]), .I1(n18_adj_4250), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [3]), .O(n20_adj_4251));
    defparam i9_4_lut_adj_974.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_975 (.I0(n15_adj_4252), .I1(n20_adj_4251), .I2(n16541), 
            .I3(\data_in[0] [6]), .O(n63_adj_4253));
    defparam i10_4_lut_adj_975.LUT_INIT = 16'hfeff;
    SB_LUT4 i20105_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4253), 
            .I2(n63), .I3(GND_net), .O(n123));   // verilog/coms.v(139[4] 142[7])
    defparam i20105_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(\data_out_frame[17] [2]), .I1(n37409), 
            .I2(n42155), .I3(n17116), .O(n43875));
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_977 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [16]), .O(n40));
    defparam i15_4_lut_adj_977.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_978 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut_adj_978.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_979 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39));
    defparam i14_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_c));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [27]), .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_42002 (.I0(byte_transmit_counter_c[1]), 
            .I1(n46588), .I2(n5_adj_4254), .I3(byte_transmit_counter_c[2]), 
            .O(n49913));
    defparam byte_transmit_counter_1__bdd_4_lut_42002.LUT_INIT = 16'he4aa;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48), .I2(n37_c), .I3(n38), .O(n16608));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_980 (.I0(n16468), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4255));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_LUT4 i20161_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_4255), .I3(\FRAME_MATCHER.i [1]), .O(n740));   // verilog/coms.v(157[9:60])
    defparam i20161_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i37293_2_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n45195));
    defparam i37293_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_981 (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[5]), .I3(GND_net), .O(n41704));
    defparam i2_3_lut_adj_981.LUT_INIT = 16'hfefe;
    SB_LUT4 i39524_3_lut (.I0(n41704), .I1(n45195), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n46678));
    defparam i39524_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(n19921), .I1(n41704), .I2(n46678), .I3(byte_transmit_counter_c[4]), 
            .O(n888));
    defparam i1_4_lut.LUT_INIT = 16'hafbb;
    SB_LUT4 i4_4_lut_adj_982 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4256));
    defparam i4_4_lut_adj_982.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_983 (.I0(\data_in[3] [4]), .I1(n10_adj_4256), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n16611));
    defparam i5_3_lut_adj_983.LUT_INIT = 16'hdfdf;
    SB_LUT4 i5_3_lut_adj_984 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4257));
    defparam i5_3_lut_adj_984.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_985 (.I0(\data_in[0] [6]), .I1(n16611), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4258));
    defparam i6_4_lut_adj_985.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_986 (.I0(n15_adj_4258), .I1(\data_in[3] [0]), .I2(n14_adj_4257), 
            .I3(\data_in[2] [2]), .O(n16476));
    defparam i8_4_lut_adj_986.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4259));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_987 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4260));
    defparam i6_4_lut_adj_987.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_988 (.I0(\data_in[3] [6]), .I1(n14_adj_4260), .I2(n10_adj_4259), 
            .I3(\data_in[2] [1]), .O(n16538));
    defparam i7_4_lut_adj_988.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_989 (.I0(n16687), .I1(n888), .I2(GND_net), .I3(GND_net), 
            .O(n41833));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'h4444;
    SB_LUT4 i8_4_lut_adj_990 (.I0(n16538), .I1(\data_in[1] [3]), .I2(n16476), 
            .I3(\data_in[1] [2]), .O(n20_adj_4261));
    defparam i8_4_lut_adj_990.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_991 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_4262));
    defparam i7_4_lut_adj_991.LUT_INIT = 16'hfeff;
    SB_LUT4 i36410_4_lut (.I0(\data_in[2] [5]), .I1(\data_in[2] [0]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n44308));
    defparam i36410_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_992 (.I0(n44308), .I1(n19_adj_4262), .I2(n20_adj_4261), 
            .I3(GND_net), .O(n63_adj_4263));
    defparam i11_3_lut_adj_992.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_adj_993 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16446), .I3(GND_net), .O(n16558));   // verilog/coms.v(225[5:23])
    defparam i2_3_lut_adj_993.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_adj_994 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n16558), .I3(GND_net), .O(n16687));   // verilog/coms.v(206[5:16])
    defparam i1_3_lut_adj_994.LUT_INIT = 16'hf7f7;
    SB_LUT4 i4_4_lut_adj_995 (.I0(n16687), .I1(n25611), .I2(n16678), .I3(n16677), 
            .O(n10_adj_4264));
    defparam i4_4_lut_adj_995.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_996 (.I0(\FRAME_MATCHER.state[0] ), .I1(n10_adj_4264), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n44325), .O(n2484));
    defparam i5_4_lut_adj_996.LUT_INIT = 16'hcc8c;
    SB_LUT4 select_366_Select_2_i5_4_lut (.I0(n123), .I1(n16680), .I2(n2857), 
            .I3(n63_adj_4263), .O(n5));
    defparam select_366_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 select_366_Select_2_i7_4_lut (.I0(n123), .I1(n16684), .I2(n3761), 
            .I3(n63_adj_4263), .O(n7));
    defparam select_366_Select_2_i7_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i20101_rep_362_2_lut (.I0(n123), .I1(n63_adj_4263), .I2(GND_net), 
            .I3(GND_net), .O(n50704));   // verilog/coms.v(143[4] 146[7])
    defparam i20101_rep_362_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_997 (.I0(n17103), .I1(Kp_23__N_1210), .I2(\data_in_frame[14]_c [7]), 
            .I3(GND_net), .O(n17509));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_997.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_998 (.I0(n42222), .I1(n42375), .I2(\data_in_frame[19] [0]), 
            .I3(n41916), .O(n12));
    defparam i5_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_999 (.I0(n28), .I1(n12), .I2(n42438), .I3(n38274), 
            .O(n38220));
    defparam i6_4_lut_adj_999.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1000 (.I0(n42216), .I1(n16), .I2(\data_in_frame[18] [7]), 
            .I3(n42299), .O(n10_adj_4268));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1001 (.I0(n41913), .I1(n10_adj_4268), .I2(n38259), 
            .I3(GND_net), .O(n16268));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_adj_1001.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4269));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1003 (.I0(n16898), .I1(n42128), .I2(n31_adj_4270), 
            .I3(n6_adj_4269), .O(n42381));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1004 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[17] [3]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[17] [5]), .O(n42360));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1005 (.I0(\data_in_frame[12] [7]), .I1(n17126), 
            .I2(n42381), .I3(n6_adj_4271), .O(n17497));   // verilog/coms.v(71[16:42])
    defparam i4_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1006 (.I0(\data_out_frame[15] [7]), .I1(n16253), 
            .I2(\data_out_frame[18] [3]), .I3(\data_out_frame[16] [3]), 
            .O(n6_adj_4272));
    defparam i1_2_lut_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[19] [7]), .I1(n42360), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4273));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1008 (.I0(\data_in_frame[13] [0]), .I1(n42414), 
            .I2(n17497), .I3(n6_adj_4273), .O(n42179));
    defparam i4_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1009 (.I0(\data_out_frame[15] [7]), .I1(n16253), 
            .I2(\data_out_frame[18] [3]), .I3(\data_out_frame[13] [5]), 
            .O(n6_adj_4274));
    defparam i1_2_lut_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1010 (.I0(n41983), .I1(n37982), .I2(n16310), 
            .I3(n42072), .O(n42289));
    defparam i2_3_lut_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(\data_in_frame[7] [7]), .I1(n42235), 
            .I2(n16804), .I3(GND_net), .O(n17396));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1012 (.I0(\data_in_frame[15] [3]), .I1(n42390), 
            .I2(n42248), .I3(Kp_23__N_1213), .O(n41962));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42097));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1014 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[17] [7]), .I3(\data_in_frame[15] [3]), .O(n42351));
    defparam i3_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1136));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1015 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4275));
    defparam i2_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1016 (.I0(Kp_23__N_1201), .I1(n7_adj_4276), .I2(n42097), 
            .I3(n8_adj_4275), .O(n42076));
    defparam i5_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1017 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[8] [4]), 
            .I2(\data_in_frame[14]_c [7]), .I3(GND_net), .O(n42268));
    defparam i2_3_lut_adj_1017.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1018 (.I0(\data_in_frame[8] [2]), .I1(n41941), 
            .I2(n17503), .I3(GND_net), .O(n42405));
    defparam i2_3_lut_adj_1018.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1019 (.I0(n16310), .I1(\data_out_frame[20] [1]), 
            .I2(n42411), .I3(GND_net), .O(n42412));
    defparam i1_2_lut_3_lut_adj_1019.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1020 (.I0(n37), .I1(\data_in_frame[12] [6]), .I2(n42268), 
            .I3(\data_in_frame[6] [1]), .O(n16_adj_4278));
    defparam i6_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4279));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1021 (.I0(n37561), .I1(n42023), .I2(n42405), 
            .I3(\data_in_frame[10] [5]), .O(n17_adj_4280));
    defparam i7_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1022 (.I0(n16310), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(n38283), .O(n43317));
    defparam i2_3_lut_4_lut_adj_1022.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(\data_in_frame[19] [2]), .I1(n17_adj_4280), 
            .I2(n15_adj_4279), .I3(n16_adj_4278), .O(n42245));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1024 (.I0(n93[1]), .I1(n63_adj_4263), .I2(n41833), 
            .I3(n2484), .O(n40980));   // verilog/coms.v(143[4] 146[7])
    defparam i1_3_lut_4_lut_adj_1024.LUT_INIT = 16'hbbb0;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17421));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i20623_2_lut_3_lut (.I0(n63), .I1(n63_adj_4253), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n93[1]));
    defparam i20623_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5_4_lut_adj_1026 (.I0(\data_in_frame[12] [3]), .I1(n8_adj_4138), 
            .I2(\data_in_frame[10] [1]), .I3(n17035), .O(n12_adj_4281));   // verilog/coms.v(70[16:41])
    defparam i5_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1027 (.I0(\data_in_frame[8] [1]), .I1(n12_adj_4281), 
            .I2(\data_in_frame[7] [5]), .I3(n17421), .O(n42140));   // verilog/coms.v(70[16:41])
    defparam i6_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1028 (.I0(n42140), .I1(n16804), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4282));
    defparam i2_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1029 (.I0(n42342), .I1(n38259), .I2(n42100), 
            .I3(\data_in_frame[14] [4]), .O(n14_adj_4283));
    defparam i6_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1030 (.I0(\data_in_frame[14]_c [3]), .I1(n14_adj_4283), 
            .I2(n10_adj_4282), .I3(n16), .O(n43329));
    defparam i7_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42357));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42188));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut (.I0(n63), .I1(n63_adj_4253), .I2(n63_adj_4263), 
            .I3(GND_net), .O(n14246));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i75_2_lut_3_lut (.I0(n740), .I1(n14246), .I2(n16683), .I3(GND_net), 
            .O(n59));   // verilog/coms.v(157[6] 159[9])
    defparam i75_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3_4_lut_adj_1033 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[8] [0]), 
            .I2(n16851), .I3(\data_in_frame[12] [4]), .O(n42462));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1034 (.I0(\data_in_frame[14]_c [2]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[12] [0]), .I3(\data_in_frame[14]_c [3]), 
            .O(n42375));
    defparam i3_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4284));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1036 (.I0(n42399), .I1(Kp_23__N_679), .I2(n17145), 
            .I3(n6_adj_4284), .O(n38274));
    defparam i4_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(n38274), .I1(n42375), .I2(GND_net), 
            .I3(GND_net), .O(n42152));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42251));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1039 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[8] [5]), .I3(GND_net), .O(n42232));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1039.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(n16804), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42372));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42447));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1042 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[6] [2]), .I3(GND_net), .O(n41941));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1042.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17535));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1044 (.I0(n740), .I1(n14246), .I2(n16563), 
            .I3(\FRAME_MATCHER.state[3] ), .O(n4_adj_4285));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1044.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut_adj_1045 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n7_adj_4201));
    defparam i1_2_lut_3_lut_adj_1045.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1046 (.I0(\data_in_frame[8] [3]), .I1(n17535), 
            .I2(n16889), .I3(n41941), .O(n10_adj_4287));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1047 (.I0(\data_in_frame[8] [1]), .I1(n10_adj_4287), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n42235));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1048 (.I0(\data_in_frame[16] [7]), .I1(n42235), 
            .I2(n42100), .I3(\data_in_frame[16] [5]), .O(n41913));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1049 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [5]), 
            .I2(\data_in_frame[10] [7]), .I3(\data_in_frame[12] [7]), .O(n42131));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42016));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1051 (.I0(n17185), .I1(Kp_23__N_729), .I2(\data_in_frame[5] [6]), 
            .I3(\data_in_frame[4] [7]), .O(n28_adj_4288));
    defparam i12_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1052 (.I0(\data_in_frame[13] [3]), .I1(n42016), 
            .I2(n42131), .I3(n41913), .O(n26_adj_4289));
    defparam i10_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1053 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_809), .I3(\data_in_frame[5] [7]), .O(n27_adj_4290));
    defparam i11_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1054 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n41144));
    defparam i1_2_lut_3_lut_adj_1054.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_1055 (.I0(\data_in_frame[9] [3]), .I1(n41968), 
            .I2(\data_in_frame[13] [7]), .I3(n42066), .O(n25_adj_4291));
    defparam i9_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1056 (.I0(n25_adj_4291), .I1(n27_adj_4290), .I2(n26_adj_4289), 
            .I3(n28_adj_4288), .O(n44019));
    defparam i15_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1057 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[13] [4]), .I3(n42435), .O(n38_adj_4292));
    defparam i15_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1058 (.I0(n42372), .I1(n42286), .I2(n42232), 
            .I3(n42219), .O(n36));
    defparam i13_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1059 (.I0(n42330), .I1(n42222), .I2(n42251), 
            .I3(n42152), .O(n37_adj_4293));
    defparam i14_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1060 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[7] [6]), .I3(\data_in_frame[9] [7]), .O(n40_adj_4294));
    defparam i17_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n35), .I1(n37_adj_4293), .I2(n36), .I3(n38_adj_4292), 
            .O(n44));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1061 (.I0(\data_in_frame[14]_c [7]), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[16] [2]), .I3(\data_in_frame[11] [2]), .O(n39_adj_4295));
    defparam i16_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1062 (.I0(n39_adj_4295), .I1(\data_in_frame[15] [0]), 
            .I2(n44), .I3(n40_adj_4294), .O(n10_adj_4296));
    defparam i1_4_lut_adj_1062.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1063 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[17] [0]), 
            .I2(n16750), .I3(n10_adj_4296), .O(n16_adj_4297));
    defparam i7_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1064 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n41254));
    defparam i1_2_lut_3_lut_adj_1064.LUT_INIT = 16'he0e0;
    SB_LUT4 i8_4_lut_adj_1065 (.I0(n42357), .I1(n16_adj_4297), .I2(n12_adj_4298), 
            .I3(\data_in_frame[15] [2]), .O(n43390));
    defparam i8_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i13157_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n18441));
    defparam i13157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42414));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16971));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42408));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1069 (.I0(\data_in_frame[9] [2]), .I1(n1), .I2(\data_in_frame[7] [1]), 
            .I3(GND_net), .O(n42286));
    defparam i2_3_lut_adj_1069.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[6] [5]), .I1(n16898), 
            .I2(GND_net), .I3(GND_net), .O(n42444));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42308));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1072 (.I0(\data_in_frame[11] [3]), .I1(n42444), 
            .I2(n42286), .I3(Kp_23__N_588), .O(n10_adj_4299));
    defparam i4_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(n37696), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42200));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1074 (.I0(\data_in_frame[7] [2]), .I1(n38325), 
            .I2(\data_in_frame[7] [0]), .I3(\data_in_frame[11] [4]), .O(n42167));
    defparam i3_4_lut_adj_1074.LUT_INIT = 16'h9669;
    SB_LUT4 data_in_frame_6__7__I_0_3242_2_lut (.I0(\data_in_frame[6] [7]), 
            .I1(\data_in_frame[6] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_588));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_6__7__I_0_3242_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1075 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n7_adj_4199));
    defparam i1_2_lut_3_lut_adj_1075.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1076 (.I0(\data_in_frame[9] [2]), .I1(n16903), 
            .I2(n37621), .I3(n42167), .O(n10_adj_4300));
    defparam i4_4_lut_adj_1076.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17145));   // verilog/coms.v(77[16:35])
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1078 (.I0(\data_in_frame[5] [1]), .I1(n41956), 
            .I2(n4_adj_4131), .I3(\data_in_frame[5] [3]), .O(n42459));
    defparam i3_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1079 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n7_adj_4197));
    defparam i1_2_lut_3_lut_adj_1079.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1080 (.I0(\data_in_frame[11] [6]), .I1(n42459), 
            .I2(n42429), .I3(n42399), .O(n43056));
    defparam i3_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(\data_in_frame[16] [2]), .I1(n15), .I2(n13), 
            .I3(n14), .O(n42121));
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1082 (.I0(\data_in_frame[18] [4]), .I1(n42121), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n42345));   // verilog/coms.v(83[17:63])
    defparam i2_3_lut_adj_1082.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1083 (.I0(n16971), .I1(n42414), .I2(n42296), 
            .I3(\data_in_frame[17] [5]), .O(n13_adj_4304));
    defparam i5_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1084 (.I0(n42121), .I1(n42079), .I2(n42213), 
            .I3(GND_net), .O(n8_adj_4305));
    defparam i3_3_lut_adj_1084.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1085 (.I0(\data_in_frame[18] [2]), .I1(n7_adj_4306), 
            .I2(\data_in_frame[18] [3]), .I3(n8_adj_4305), .O(n42158));
    defparam i2_4_lut_adj_1085.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1086 (.I0(n42158), .I1(n37587), .I2(n37485), 
            .I3(n42345), .O(n10_adj_4307));
    defparam i4_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_in_frame[19] [1]), .I1(n42245), 
            .I2(GND_net), .I3(GND_net), .O(n41888));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1088 (.I0(n42311), .I1(\data_in_frame[15] [4]), 
            .I2(n41962), .I3(\data_in_frame[19] [3]), .O(n14_adj_4308));
    defparam i6_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1089 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16521));
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(n42076), .I1(n41888), .I2(n10_adj_4307), 
            .I3(Kp_23__N_1136), .O(n9));
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1091 (.I0(n9), .I1(n14_adj_4308), .I2(n42179), 
            .I3(\data_in_frame[14] [6]), .O(n38270));
    defparam i7_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[13] [7]), .I1(n43056), 
            .I2(GND_net), .I3(GND_net), .O(n38228));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1093 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[14]_c [2]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n42085));
    defparam i2_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n16893), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42128));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1095 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n7_adj_4195));
    defparam i1_2_lut_3_lut_adj_1095.LUT_INIT = 16'he0e0;
    SB_LUT4 i15_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47));
    defparam i15_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1096 (.I0(n15_c), .I1(\data_in_frame[9] [1]), .I2(\data_in_frame[7] [0]), 
            .I3(\data_in_frame[11] [2]), .O(n42396));   // verilog/coms.v(70[16:41])
    defparam i3_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n13980));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1098 (.I0(\data_in_frame[6] [5]), .I1(n42396), 
            .I2(n41968), .I3(\data_in_frame[6] [7]), .O(n17103));   // verilog/coms.v(77[16:35])
    defparam i3_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_in_frame[13] [4]), .I1(n17103), 
            .I2(GND_net), .I3(GND_net), .O(n42432));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1100 (.I0(n25891), .I1(n25307), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n6_adj_4309));
    defparam i2_4_lut_adj_1100.LUT_INIT = 16'h5d55;
    SB_LUT4 i1_2_lut_3_lut_adj_1101 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n41252));
    defparam i1_2_lut_3_lut_adj_1101.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1102 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n41250));
    defparam i1_2_lut_3_lut_adj_1102.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(n26154), .I1(n6_adj_4309), .I2(n25299), 
            .I3(n16521), .O(n4497));
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1104 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n7_adj_4194));
    defparam i1_2_lut_3_lut_adj_1104.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1105 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n41248));
    defparam i1_2_lut_3_lut_adj_1105.LUT_INIT = 16'he0e0;
    SB_LUT4 i20260_3_lut (.I0(n4497), .I1(\FRAME_MATCHER.state[0] ), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n25520));
    defparam i20260_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42134));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i20030_2_lut_3_lut (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n25288));
    defparam i20030_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42336));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1108 (.I0(n42336), .I1(n17168), .I2(n42134), 
            .I3(n31_adj_4270), .O(n14_adj_4310));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1109 (.I0(\data_in_frame[8] [7]), .I1(n14_adj_4310), 
            .I2(n10_adj_4311), .I3(\data_in_frame[11] [0]), .O(Kp_23__N_1210));   // verilog/coms.v(73[16:43])
    defparam i7_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_in_frame[6] [7]), .I1(n17168), 
            .I2(GND_net), .I3(GND_net), .O(n42327));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_in_frame[7] [3]), .I1(n37621), 
            .I2(GND_net), .I3(GND_net), .O(n38259));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(n37696), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42116));
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1113 (.I0(\data_in_frame[7] [1]), .I1(n42116), 
            .I2(\data_in_frame[11] [5]), .I3(n38259), .O(n12_adj_4312));
    defparam i5_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1114 (.I0(\data_in_frame[5] [0]), .I1(n12_adj_4312), 
            .I2(n42327), .I3(n38325), .O(n37512));
    defparam i6_4_lut_adj_1114.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(n37512), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42213));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_in_frame[13] [5]), .I1(n42296), 
            .I2(GND_net), .I3(GND_net), .O(n41910));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(Kp_23__N_1210), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17415));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1118 (.I0(n41910), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[16] [0]), .I3(n42213), .O(n10_adj_4313));
    defparam i4_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[17] [7]), 
            .I2(n10_adj_4313), .I3(\data_in_frame[13] [6]), .O(n37587));
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4314));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4315));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39138_2_lut (.I0(\data_out_frame[22] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46582));
    defparam i39138_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4316));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4317));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4318));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39292_2_lut (.I0(\data_out_frame[22] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46583));
    defparam i39292_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4319));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4320));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4321));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39287_2_lut (.I0(\data_out_frame[22] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46584));
    defparam i39287_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4322));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4323));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1120 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n41246));
    defparam i1_2_lut_3_lut_adj_1120.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4324));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39281_2_lut (.I0(\data_out_frame[22] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46585));
    defparam i39281_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1121 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n41244));
    defparam i1_2_lut_3_lut_adj_1121.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4325));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4254));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39431_2_lut (.I0(\data_out_frame[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46588));
    defparam i39431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1122 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n41242));
    defparam i1_2_lut_3_lut_adj_1122.LUT_INIT = 16'he0e0;
    SB_LUT4 i41185_2_lut (.I0(n14246), .I1(n16676), .I2(GND_net), .I3(GND_net), 
            .O(n42487));
    defparam i41185_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n7_adj_4192));
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n41240));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n7_adj_4190));
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1126 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n7_adj_4188));
    defparam i1_2_lut_3_lut_adj_1126.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n7_adj_4186));
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n41346));
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4236));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4235));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n41344));
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1130 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n41342));
    defparam i1_2_lut_3_lut_adj_1130.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n41334));
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1132 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n41282));
    defparam i1_2_lut_3_lut_adj_1132.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1133 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n41270));
    defparam i1_2_lut_3_lut_adj_1133.LUT_INIT = 16'he0e0;
    SB_LUT4 i12_4_lut_adj_1134 (.I0(tx_active), .I1(r_SM_Main_c[1]), .I2(n10142), 
            .I3(n4_adj_4326), .O(n41424));   // verilog/uart_tx.v(31[16:25])
    defparam i12_4_lut_adj_1134.LUT_INIT = 16'h32aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1135 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n41268));
    defparam i1_2_lut_3_lut_adj_1135.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n41266));
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'he0e0;
    SB_LUT4 i39278_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46589));
    defparam i39278_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4234));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1137 (.I0(n4_adj_4286), .I1(n141), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n41264));
    defparam i1_2_lut_3_lut_adj_1137.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1138 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [31]), .O(n8_adj_4202));
    defparam i1_2_lut_4_lut_adj_1138.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1139 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [30]), .O(n40964));
    defparam i1_2_lut_4_lut_adj_1139.LUT_INIT = 16'hfe00;
    SB_LUT4 i12998_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n18282));
    defparam i12998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12999_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n18283));
    defparam i12999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13000_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n18284));
    defparam i13000_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13001_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n18285));
    defparam i13001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1140 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [27]), .O(n8_adj_4198));
    defparam i1_2_lut_4_lut_adj_1140.LUT_INIT = 16'hfe00;
    SB_LUT4 i20031_2_lut_4_lut (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [23]), .O(n25290));
    defparam i20031_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i13002_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n18286));
    defparam i13002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1141 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [15]), .O(n8_adj_4191));
    defparam i1_2_lut_4_lut_adj_1141.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1142 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [14]), .O(n8_adj_4189));
    defparam i1_2_lut_4_lut_adj_1142.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1143 (.I0(n4_adj_4327), .I1(n59), .I2(n26_adj_4328), 
            .I3(\FRAME_MATCHER.state [13]), .O(n8_adj_4187));
    defparam i1_2_lut_4_lut_adj_1143.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1144 (.I0(n59), .I1(n26_adj_4328), .I2(n4_adj_4327), 
            .I3(\FRAME_MATCHER.state [28]), .O(n8_adj_4200));
    defparam i1_2_lut_4_lut_adj_1144.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1145 (.I0(n59), .I1(n26_adj_4328), .I2(n4_adj_4327), 
            .I3(\FRAME_MATCHER.state [26]), .O(n8_adj_4196));
    defparam i1_2_lut_4_lut_adj_1145.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1146 (.I0(n59), .I1(n26_adj_4328), .I2(n4_adj_4327), 
            .I3(\FRAME_MATCHER.state [17]), .O(n8_adj_4193));
    defparam i1_2_lut_4_lut_adj_1146.LUT_INIT = 16'hfe00;
    SB_LUT4 select_331_Select_1_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n3_adj_4238));
    defparam select_331_Select_1_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_31_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [31]), .I3(GND_net), .O(n3_adj_4185));
    defparam select_331_Select_31_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_30_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [30]), .I3(GND_net), .O(n3_adj_4183));
    defparam select_331_Select_30_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13003_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n18287));
    defparam i13003_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_331_Select_29_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [29]), .I3(GND_net), .O(n3_adj_4181));
    defparam select_331_Select_29_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_28_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [28]), .I3(GND_net), .O(n3_adj_4179));
    defparam select_331_Select_28_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_27_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [27]), .I3(GND_net), .O(n3_adj_4177));
    defparam select_331_Select_27_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_26_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [26]), .I3(GND_net), .O(n3_adj_4175));
    defparam select_331_Select_26_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_25_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [25]), .I3(GND_net), .O(n3_adj_4173));
    defparam select_331_Select_25_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_24_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [24]), .I3(GND_net), .O(n3_adj_4171));
    defparam select_331_Select_24_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_23_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [23]), .I3(GND_net), .O(n3_adj_4169));
    defparam select_331_Select_23_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_22_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [22]), .I3(GND_net), .O(n3_adj_4167));
    defparam select_331_Select_22_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_21_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [21]), .I3(GND_net), .O(n3_adj_4165));
    defparam select_331_Select_21_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_20_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [20]), .I3(GND_net), .O(n3_adj_4164));
    defparam select_331_Select_20_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_19_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [19]), .I3(GND_net), .O(n3_adj_4163));
    defparam select_331_Select_19_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13004_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n18288));
    defparam i13004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_331_Select_18_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [18]), .I3(GND_net), .O(n3_adj_4162));
    defparam select_331_Select_18_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_17_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [17]), .I3(GND_net), .O(n3_adj_4161));
    defparam select_331_Select_17_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_16_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [16]), .I3(GND_net), .O(n3_adj_4160));
    defparam select_331_Select_16_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_15_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [15]), .I3(GND_net), .O(n3_adj_4159));
    defparam select_331_Select_15_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_14_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [14]), .I3(GND_net), .O(n3_adj_4158));
    defparam select_331_Select_14_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_13_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [13]), .I3(GND_net), .O(n3_adj_4157));
    defparam select_331_Select_13_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_12_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [12]), .I3(GND_net), .O(n3_adj_4156));
    defparam select_331_Select_12_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_11_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [11]), .I3(GND_net), .O(n3_adj_4155));
    defparam select_331_Select_11_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4232));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4231));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_331_Select_10_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [10]), .I3(GND_net), .O(n3_adj_4154));
    defparam select_331_Select_10_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_9_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [9]), .I3(GND_net), .O(n3_adj_4153));
    defparam select_331_Select_9_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_8_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n3_adj_4152));
    defparam select_331_Select_8_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13005_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n18289));
    defparam i13005_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_331_Select_7_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [7]), .I3(GND_net), .O(n3_adj_4151));
    defparam select_331_Select_7_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_6_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [6]), .I3(GND_net), .O(n3_adj_4150));
    defparam select_331_Select_6_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_5_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n3_adj_4149));
    defparam select_331_Select_5_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i17_3_lut (.I0(n25630), .I1(\FRAME_MATCHER.state_31__N_2275 [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n6_adj_4233));
    defparam i17_3_lut.LUT_INIT = 16'h5c5c;
    SB_LUT4 mux_1090_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n4446));
    defparam mux_1090_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_331_Select_4_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n3_adj_4148));
    defparam select_331_Select_4_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_1090_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16] [1]), .O(n4447));
    defparam mux_1090_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1090_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n4448));
    defparam mux_1090_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_331_Select_3_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n3_adj_4145));
    defparam select_331_Select_3_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_1090_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n4449));
    defparam mux_1090_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_331_Select_2_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n3_adj_4120));
    defparam select_331_Select_2_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_331_Select_0_i3_2_lut_3_lut (.I0(n25611), .I1(n16676), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n3_c));
    defparam select_331_Select_0_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_1090_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n4450));
    defparam mux_1090_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i39276_2_lut (.I0(\data_out_frame[22] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46590));
    defparam i39276_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4230));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20028_2_lut_2_lut_3_lut (.I0(n25611), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n25285));
    defparam i20028_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1147 (.I0(\FRAME_MATCHER.state_31__N_2275 [3]), 
            .I1(\FRAME_MATCHER.state [2]), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n3735), .O(n14276));
    defparam i2_3_lut_4_lut_adj_1147.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n4_adj_4329));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0504;
    SB_LUT4 n49913_bdd_4_lut_4_lut (.I0(\data_out_frame[0] [4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter_c[2]), .I3(n49913), .O(n49916));
    defparam n49913_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4226));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4225));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1148 (.I0(n16851), .I1(n16889), .I2(n8_adj_4138), 
            .I3(\data_in_frame[8] [3]), .O(n17126));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1149 (.I0(n16851), .I1(n16889), .I2(\data_in_frame[6] [2]), 
            .I3(GND_net), .O(n31_adj_4270));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 i38949_2_lut (.I0(\data_out_frame[22] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46604));
    defparam i38949_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4224));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_339_i3_3_lut_4_lut (.I0(n31_adj_4140), .I1(n25297), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n16679), .O(n3));
    defparam equal_339_i3_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1150 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(n42128), .O(n41968));   // verilog/coms.v(77[16:35])
    defparam i1_2_lut_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1151 (.I0(\data_in_frame[15] [1]), .I1(n17103), 
            .I2(Kp_23__N_1210), .I3(\data_in_frame[14]_c [7]), .O(n42393));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(n16903), .O(n10_adj_4311));   // verilog/coms.v(77[16:35])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1152 (.I0(n16772), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(\data_out_frame[14] [0]), 
            .O(n6_adj_4331));
    defparam i1_2_lut_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_1153 (.I0(n42450), .I1(n42308), .I2(n43390), 
            .I3(n13_adj_4304), .O(n37485));
    defparam i1_4_lut_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1154 (.I0(n16772), .I1(n10_adj_4332), .I2(\data_out_frame[5] [5]), 
            .I3(n42049), .O(n37697));
    defparam i1_2_lut_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1155 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n41965));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_3_lut_adj_1155.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1156 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n42280));
    defparam i1_2_lut_3_lut_adj_1156.LUT_INIT = 16'h9696;
    SB_LUT4 i39293_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n47196));   // verilog/coms.v(104[34:55])
    defparam i39293_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4333));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36473_4_lut (.I0(n5_adj_4333), .I1(n47196), .I2(n45195), 
            .I3(byte_transmit_counter[0]), .O(n44375));
    defparam i36473_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i36475_4_lut (.I0(n44375), .I1(n49874), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44377));
    defparam i36475_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36474_3_lut (.I0(n49838), .I1(n49826), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44376));
    defparam i36474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1157 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(n16994), .I3(n42203), .O(n42456));
    defparam i2_3_lut_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i39288_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47191));   // verilog/coms.v(104[34:55])
    defparam i39288_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4334));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16675));   // verilog/coms.v(148[5:9])
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'heeee;
    SB_LUT4 i36470_4_lut (.I0(n5_adj_4334), .I1(n47191), .I2(n45195), 
            .I3(byte_transmit_counter[0]), .O(n44372));
    defparam i36470_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i36472_4_lut (.I0(n44372), .I1(n49880), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44374));
    defparam i36472_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36471_3_lut (.I0(n49850), .I1(n49844), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44373));
    defparam i36471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1159 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[6] [2]), .O(n42241));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n47184));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4335));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36467_4_lut (.I0(n5_adj_4335), .I1(byte_transmit_counter[0]), 
            .I2(n45195), .I3(n47184), .O(n44369));
    defparam i36467_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i36469_4_lut (.I0(n44369), .I1(n49886), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44371));
    defparam i36469_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36468_3_lut (.I0(n49988), .I1(n49856), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44370));
    defparam i36468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1160 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[11] [5]), .O(n42039));
    defparam i2_3_lut_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i40679_3_lut (.I0(n49958), .I1(n49820), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n48582));
    defparam i40679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40683_3_lut (.I0(n49916), .I1(n48582), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n48586));   // verilog/coms.v(104[34:55])
    defparam i40683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1161 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n42210));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i40684_4_lut (.I0(n48586), .I1(n49892), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i40684_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i38989_2_lut (.I0(\data_out_frame[0] [3]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46613));   // verilog/coms.v(104[34:55])
    defparam i38989_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n46613), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_4336));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4337));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36464_3_lut (.I0(n5_adj_4337), .I1(n6_adj_4336), .I2(n45195), 
            .I3(GND_net), .O(n44366));
    defparam i36464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n17004));
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 i36466_4_lut (.I0(n44366), .I1(n49928), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44368));
    defparam i36466_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1163 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[6] [2]), .O(n6_adj_4338));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1164 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[12] [6]), 
            .I2(n41971), .I3(GND_net), .O(n6_adj_4339));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1165 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n42462), .I3(\data_in_frame[16] [6]), .O(n42222));
    defparam i2_3_lut_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i39439_2_lut (.I0(\data_out_frame[0] [2]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46610));   // verilog/coms.v(104[34:55])
    defparam i39439_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(n46610), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_4340));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4341));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36461_3_lut (.I0(n5_adj_4341), .I1(n6_adj_4340), .I2(n45195), 
            .I3(GND_net), .O(n44363));
    defparam i36461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36463_4_lut (.I0(n44363), .I1(n49934), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44365));
    defparam i36463_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut_adj_1166 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n42225));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1167 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n42200), .I3(n17185), .O(n38230));
    defparam i2_3_lut_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1168 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[11] [7]), .I3(\data_in_frame[10] [0]), .O(n42342));
    defparam i1_2_lut_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i39266_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47168));   // verilog/coms.v(104[34:55])
    defparam i39266_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4342));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36458_4_lut (.I0(n5_adj_4342), .I1(n47168), .I2(n45195), 
            .I3(byte_transmit_counter[0]), .O(n44360));
    defparam i36458_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i36460_4_lut (.I0(n44360), .I1(n49940), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44362));
    defparam i36460_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n41952));
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1170 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n42219), .I3(\data_in_frame[10] [0]), .O(n6));
    defparam i1_2_lut_3_lut_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i17_3_lut_4_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(n34), .I3(\data_out_frame[18] [3]), .O(n39_adj_4344));
    defparam i17_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1171 (.I0(n42109), .I1(n42314), .I2(\data_out_frame[17] [4]), 
            .I3(\data_out_frame[20] [0]), .O(n42292));
    defparam i1_2_lut_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1172 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[13] [2]), .I3(\data_out_frame[13] [3]), 
            .O(n42271));
    defparam i2_3_lut_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1173 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[11] [2]), .O(n42366));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1174 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n42019));
    defparam i1_2_lut_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_out_frame[9] [2]), .I1(n42283), .I2(\data_out_frame[8] [7]), 
            .I3(\data_out_frame[13] [3]), .O(n16_adj_4345));   // verilog/coms.v(73[16:27])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1175 (.I0(n37982), .I1(n17304), .I2(n42289), 
            .I3(GND_net), .O(n42290));
    defparam i1_2_lut_3_lut_adj_1175.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1176 (.I0(\data_out_frame[20] [3]), .I1(n17304), 
            .I2(n17301), .I3(\data_out_frame[20] [2]), .O(n43126));
    defparam i2_3_lut_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1177 (.I0(\FRAME_MATCHER.state[3] ), .I1(n14246), 
            .I2(n2484), .I3(n141), .O(n40984));
    defparam i1_3_lut_4_lut_adj_1177.LUT_INIT = 16'haa80;
    SB_LUT4 mux_1090_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n4451));
    defparam mux_1090_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i36443_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44345));
    defparam i36443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36444_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44346));
    defparam i36444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36447_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44349));
    defparam i36447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36446_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44348));
    defparam i36446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1090_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n4452));
    defparam mux_1090_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i36437_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44339));
    defparam i36437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36438_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44340));
    defparam i36438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36441_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44343));
    defparam i36441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36440_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44342));
    defparam i36440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36431_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44333));
    defparam i36431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36432_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44334));
    defparam i36432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36435_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44337));
    defparam i36435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36434_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n44336));
    defparam i36434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n17283), .I1(n42450), .I2(\data_in_frame[13] [7]), 
            .I3(n43056), .O(n7_adj_4306));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1178 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n26154), .I3(GND_net), .O(n4_adj_4346));
    defparam i1_2_lut_3_lut_adj_1178.LUT_INIT = 16'hfefe;
    SB_LUT4 i13070_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n18354));
    defparam i13070_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_714_i1_3_lut_4_lut (.I0(n31), .I1(n25297), .I2(tx_transmit_N_2998), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n26152));   // verilog/coms.v(147[4] 288[11])
    defparam mux_714_i1_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 mux_1090_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n4453));
    defparam mux_1090_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i34617_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n26154), .I3(n2_adj_4347), .O(n42491));
    defparam i34617_4_lut_4_lut.LUT_INIT = 16'hfbf8;
    SB_LUT4 i1_2_lut_3_lut_adj_1179 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n2_adj_4347));
    defparam i1_2_lut_3_lut_adj_1179.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13071_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n18355));
    defparam i13071_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36420_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[3]), 
            .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter_c[1]), 
            .O(n44320));   // verilog/coms.v(100[12:33])
    defparam i36420_3_lut_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 i13072_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n18356));
    defparam i13072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18665_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(\data_in_frame[11] [3]), 
            .I3(rx_data[3]), .O(n23932));
    defparam i18665_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13074_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n18358));
    defparam i13074_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[7]), .I3(GND_net), .O(n42664));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'hfefe;
    SB_LUT4 i41873_4_lut (.I0(n42664), .I1(r_SM_Main_2__N_3106[0]), .I2(n44320), 
            .I3(tx_active), .O(tx_transmit_N_2998));
    defparam i41873_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_732_i1_4_lut (.I0(n25307), .I1(n26152), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n26156));   // verilog/coms.v(147[4] 288[11])
    defparam mux_732_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i38867_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n26156), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n4_adj_4346), .O(n46769));   // verilog/coms.v(147[4] 288[11])
    defparam i38867_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i13075_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n18359));
    defparam i13075_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1090_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n4454));
    defparam mux_1090_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13076_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n18360));
    defparam i13076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1090_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n4455));
    defparam mux_1090_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13077_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n18361));
    defparam i13077_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1090_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n4456));
    defparam mux_1090_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1181 (.I0(n17283), .I1(n42450), .I2(n42351), 
            .I3(\data_in_frame[13] [5]), .O(n7_adj_4276));
    defparam i1_3_lut_4_lut_adj_1181.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1090_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n4457));
    defparam mux_1090_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1090_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n4458));
    defparam mux_1090_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1090_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n4459));
    defparam mux_1090_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1090_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n4460));
    defparam mux_1090_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_41992 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4325), .I2(n46585), .I3(byte_transmit_counter_c[2]), 
            .O(n49889));
    defparam byte_transmit_counter_1__bdd_4_lut_41992.LUT_INIT = 16'he4aa;
    SB_LUT4 n49889_bdd_4_lut (.I0(n49889), .I1(n17_adj_4324), .I2(n16_adj_4323), 
            .I3(byte_transmit_counter_c[2]), .O(n49892));
    defparam n49889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1090_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n4461));
    defparam mux_1090_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\FRAME_MATCHER.state [29]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n40982));
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h8888;
    SB_LUT4 i34810_2_lut_4_lut (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[7]), .I3(n44320), .O(n42696));
    defparam i34810_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1183 (.I0(n17037), .I1(n41956), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n38325));
    defparam i1_2_lut_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1184 (.I0(Kp_23__N_1213), .I1(\data_in_frame[13] [4]), 
            .I2(n17103), .I3(\data_in_frame[13] [3]), .O(n42296));
    defparam i2_3_lut_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i20631_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n25891));
    defparam i20631_4_lut_4_lut.LUT_INIT = 16'h4046;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\FRAME_MATCHER.state [25]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41026));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\FRAME_MATCHER.state [24]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41028));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1187 (.I0(Kp_23__N_676), .I1(\data_in_frame[4] [6]), 
            .I2(n42435), .I3(n1), .O(n42399));
    defparam i2_3_lut_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1188 (.I0(\data_in_frame[7] [2]), .I1(n37696), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n42435));
    defparam i1_2_lut_3_lut_adj_1188.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[5] [0]), .I1(n10_adj_4300), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[6] [6]), .O(n17283));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1189 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(n10_adj_4299), .I3(n16), .O(n42450));
    defparam i5_3_lut_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\FRAME_MATCHER.state [22]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41030));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h8888;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n12_adj_4298));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(\FRAME_MATCHER.state [21]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41032));
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h8888;
    SB_LUT4 i12_3_lut_4_lut (.I0(\data_in_frame[12] [3]), .I1(n44019), .I2(\data_in_frame[10] [6]), 
            .I3(\data_in_frame[11] [1]), .O(n35));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\FRAME_MATCHER.state [20]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41034));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1193 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n42100));
    defparam i1_2_lut_3_lut_adj_1193.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\FRAME_MATCHER.state [19]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41036));
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\FRAME_MATCHER.state [18]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41038));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1196 (.I0(n17283), .I1(\data_in_frame[13] [5]), 
            .I2(n42296), .I3(\data_in_frame[15] [4]), .O(n16750));
    defparam i2_3_lut_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1090_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14] [0]), .O(n4462));
    defparam mux_1090_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1197 (.I0(n41983), .I1(n37982), .I2(\data_out_frame[20] [4]), 
            .I3(\data_out_frame[20] [3]), .O(n42174));
    defparam i1_2_lut_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(\FRAME_MATCHER.state [16]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n40988));
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1199 (.I0(\data_in_frame[7] [7]), .I1(n42235), 
            .I2(n16804), .I3(\data_in_frame[19] [5]), .O(n42390));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1200 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[8] [5]), .I3(n42405), .O(n6_adj_4271));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(\data_in_frame[14]_c [3]), .I1(\data_in_frame[17] [0]), 
            .I2(n42066), .I3(GND_net), .O(n42299));
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1202 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n38220), .I3(GND_net), .O(n42149));
    defparam i1_2_lut_3_lut_adj_1202.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1203 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[6] [0]), .O(n42438));
    defparam i1_2_lut_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1204 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n17325));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1205 (.I0(n16903), .I1(\data_in_frame[6] [5]), 
            .I2(n16898), .I3(GND_net), .O(n16938));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(\FRAME_MATCHER.state [12]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41040));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\FRAME_MATCHER.state [11]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41050));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\FRAME_MATCHER.state [10]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n40966));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\FRAME_MATCHER.state [9]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41060));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\FRAME_MATCHER.state [8]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41052));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\FRAME_MATCHER.state [7]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41042));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1090_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14] [1]), .O(n4463));
    defparam mux_1090_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\FRAME_MATCHER.state [6]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41044));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\FRAME_MATCHER.state [5]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n41046));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1214 (.I0(n26_adj_4328), .I1(n4_adj_4327), .I2(n16682), 
            .I3(n4_adj_4285), .O(n7_adj_4348));
    defparam i2_4_lut_adj_1214.LUT_INIT = 16'hefee;
    SB_LUT4 mux_1090_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14]_c [2]), .O(n4464));
    defparam mux_1090_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\FRAME_MATCHER.state [4]), .I1(n7_adj_4348), 
            .I2(GND_net), .I3(GND_net), .O(n40986));
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1216 (.I0(n3761), .I1(n16684), .I2(n14246), .I3(GND_net), 
            .O(n141));   // verilog/coms.v(244[5:25])
    defparam i1_3_lut_adj_1216.LUT_INIT = 16'h1010;
    SB_LUT4 i159_2_lut (.I0(n14246), .I1(n2484), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4327));
    defparam i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i155_3_lut (.I0(n16687), .I1(n888), .I2(n14246), .I3(GND_net), 
            .O(n4_adj_4286));   // verilog/coms.v(113[11:12])
    defparam i155_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_4_lut_adj_1217 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16446), .I3(n16675), .O(n16678));   // verilog/coms.v(195[5:24])
    defparam i2_3_lut_4_lut_adj_1217.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_3_lut_adj_1218 (.I0(n16680), .I1(n2857), .I2(n14246), .I3(GND_net), 
            .O(n26_adj_4328));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1218.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_adj_1219 (.I0(n26_adj_4328), .I1(n59), .I2(n4_adj_4286), 
            .I3(GND_net), .O(n42784));
    defparam i2_3_lut_adj_1219.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1220 (.I0(\FRAME_MATCHER.state_31__N_2275 [3]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n16677), .I3(n42784), .O(n41172));
    defparam i1_4_lut_adj_1220.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1221 (.I0(n16558), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n16677));   // verilog/coms.v(161[5:29])
    defparam i1_2_lut_3_lut_adj_1221.LUT_INIT = 16'hfefe;
    SB_LUT4 i34727_2_lut (.I0(n16684), .I1(n3761), .I2(GND_net), .I3(GND_net), 
            .O(n42610));
    defparam i34727_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1090_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14]_c [3]), .O(n4465));
    defparam mux_1090_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in[3] [4]), .I1(n10_adj_4256), .I2(\data_in[2] [7]), 
            .I3(\data_in[3] [0]), .O(n15_adj_4252));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_3_lut_adj_1222 (.I0(n16558), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n16684));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_3_lut_adj_1222.LUT_INIT = 16'hefef;
    SB_LUT4 select_366_Select_1_i5_4_lut (.I0(n63_adj_4263), .I1(n16680), 
            .I2(n2857), .I3(n93[1]), .O(n5_adj_4349));
    defparam select_366_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i2_4_lut_adj_1223 (.I0(n93[1]), .I1(n5_adj_4349), .I2(n42610), 
            .I3(n63_adj_4263), .O(n6_adj_4350));
    defparam i2_4_lut_adj_1223.LUT_INIT = 16'hcecf;
    SB_LUT4 i3_4_lut_adj_1224 (.I0(n16678), .I1(n6_adj_4350), .I2(\FRAME_MATCHER.state_31__N_2243 [1]), 
            .I3(n16683), .O(n50161));
    defparam i3_4_lut_adj_1224.LUT_INIT = 16'hddfd;
    SB_LUT4 mux_1090_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[14] [4]), .O(n4466));
    defparam mux_1090_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1090_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14] [5]), .O(n4467));
    defparam mux_1090_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(n37905), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42094));
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1226 (.I0(\data_out_frame[20] [4]), .I1(n42094), 
            .I2(n17301), .I3(n41983), .O(n43726));
    defparam i2_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1227 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[8] [4]), .O(n6_adj_4351));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1090_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14]_c [7]), .O(n4469));
    defparam mux_1090_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1228 (.I0(n17304), .I1(n42265), .I2(n42441), 
            .I3(n42137), .O(n22_adj_4352));   // verilog/coms.v(73[16:27])
    defparam i9_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[17] [5]), .I1(n42387), .I2(\data_out_frame[10] [6]), 
            .I3(GND_net), .O(n20_adj_4353));   // verilog/coms.v(73[16:27])
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1229 (.I0(n42109), .I1(n22_adj_4352), .I2(n16_adj_4345), 
            .I3(n42465), .O(n24_adj_4354));   // verilog/coms.v(73[16:27])
    defparam i11_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i41182_2_lut_3_lut_3_lut (.I0(n3735), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n17676));
    defparam i41182_2_lut_3_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i12_4_lut_adj_1230 (.I0(\data_out_frame[6] [5]), .I1(n24_adj_4354), 
            .I2(n20_adj_4353), .I3(\data_out_frame[6] [4]), .O(n16310));   // verilog/coms.v(73[16:27])
    defparam i12_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42265));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1232 (.I0(\data_out_frame[9] [2]), .I1(n42283), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n42207));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(n42207), .I1(n42366), .I2(\data_out_frame[7] [0]), 
            .I3(GND_net), .O(n16249));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1234 (.I0(n42420), .I1(n16249), .I2(\data_out_frame[13] [7]), 
            .I3(n42426), .O(n10_adj_4355));
    defparam i4_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1235 (.I0(n42321), .I1(n10_adj_4355), .I2(n16691), 
            .I3(GND_net), .O(n37982));
    defparam i5_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(n37982), .I1(n17304), .I2(GND_net), 
            .I3(GND_net), .O(n38283));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1237 (.I0(n42292), .I1(n16249), .I2(n42019), 
            .I3(n42402), .O(n10_adj_4356));
    defparam i4_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1238 (.I0(n42423), .I1(n10_adj_4356), .I2(n42265), 
            .I3(GND_net), .O(n42411));
    defparam i5_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(n42289), .I1(n42411), .I2(n38283), 
            .I3(GND_net), .O(n43711));
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[19] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42465));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1090_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n25299), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14] [6]), .O(n4468));
    defparam mux_1090_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1241 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n42137));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1242 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[16] [0]), .I3(n42137), .O(n10_adj_4357));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1243 (.I0(n42339), .I1(n10_adj_4357), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n42321));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_adj_1243.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42173));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1245 (.I0(n17424), .I1(\data_out_frame[6] [2]), 
            .I2(n41952), .I3(n6_adj_4351), .O(n42423));
    defparam i4_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42402));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1247 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[13] [5]), .I3(GND_net), .O(n42363));
    defparam i2_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1248 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[3] [7]), .O(n6_adj_4133));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1249 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[18] [2]), 
            .I2(n42274), .I3(n41885), .O(n16_adj_4358));   // verilog/coms.v(70[16:41])
    defparam i6_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1250 (.I0(\data_out_frame[13] [4]), .I1(n42046), 
            .I2(n42366), .I3(\data_out_frame[16] [0]), .O(n17_adj_4359));   // verilog/coms.v(70[16:41])
    defparam i7_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1251 (.I0(n17_adj_4359), .I1(\data_out_frame[16] [1]), 
            .I2(n16_adj_4358), .I3(n1185), .O(n17301));   // verilog/coms.v(70[16:41])
    defparam i9_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1252 (.I0(\data_out_frame[6] [3]), .I1(n42029), 
            .I2(n42363), .I3(\data_out_frame[13] [4]), .O(n20_adj_4360));   // verilog/coms.v(72[16:27])
    defparam i8_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1253 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[18] [0]), 
            .I2(n42271), .I3(n41980), .O(n19_adj_4361));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1254 (.I0(n17430), .I1(\data_out_frame[11] [0]), 
            .I2(n42225), .I3(\data_out_frame[8] [4]), .O(n21));   // verilog/coms.v(72[16:27])
    defparam i9_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1255 (.I0(n21), .I1(n19_adj_4361), .I2(n20_adj_4360), 
            .I3(GND_net), .O(n17304));   // verilog/coms.v(72[16:27])
    defparam i11_3_lut_adj_1255.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1256 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[1] [3]), .O(Kp_23__N_729));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(n17304), .I1(n17301), .I2(GND_net), 
            .I3(GND_net), .O(n42026));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_4_lut_adj_1258 (.I0(n63_adj_4263), .I1(n740), .I2(n41833), 
            .I3(n16683), .O(n5_adj_15));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut_adj_1258.LUT_INIT = 16'ha0a2;
    SB_LUT4 i20630_2_lut_3_lut (.I0(n63_adj_4263), .I1(n740), .I2(n93[1]), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2243 [1]));   // verilog/coms.v(157[6] 159[9])
    defparam i20630_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_out_frame[15] [5]), .I1(n1515), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4363));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1260 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(n37540), .I3(n6_adj_4363), .O(n42420));
    defparam i4_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1261 (.I0(n37514), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[18] [4]), .I3(n6_adj_4272), .O(n37905));
    defparam i4_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1262 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[9] [1]), .I3(GND_net), .O(n42046));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1263 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4364));   // verilog/coms.v(83[17:70])
    defparam i2_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1264 (.I0(n42046), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[7] [2]), .O(n14_adj_4365));   // verilog/coms.v(83[17:70])
    defparam i6_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1265 (.I0(\data_out_frame[5] [1]), .I1(n14_adj_4365), 
            .I2(n10_adj_4364), .I3(\data_out_frame[9] [3]), .O(n1515));   // verilog/coms.v(83[17:70])
    defparam i7_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[13] [5]), .I1(n16815), 
            .I2(GND_net), .I3(GND_net), .O(n41885));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(\data_out_frame[13] [6]), .I1(n42035), 
            .I2(n1515), .I3(GND_net), .O(n42277));
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1268 (.I0(n37471), .I1(n42277), .I2(n42009), 
            .I3(n41885), .O(n37514));
    defparam i3_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i9_3_lut (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [2]), 
            .I2(n37514), .I3(GND_net), .O(n26_adj_4366));
    defparam i9_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1269 (.I0(n42197), .I1(n16989), .I2(n41986), 
            .I3(\data_out_frame[15] [4]), .O(n29_adj_4367));
    defparam i12_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1270 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[15] [3]), .I3(n42420), .O(n28_adj_4368));
    defparam i11_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1271 (.I0(n29_adj_4367), .I1(\data_out_frame[15] [2]), 
            .I2(n26_adj_4366), .I3(\data_out_frame[17] [4]), .O(n32));
    defparam i15_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1272 (.I0(n42363), .I1(n42456), .I2(\data_out_frame[12] [5]), 
            .I3(n42161), .O(n27_adj_4369));
    defparam i10_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1273 (.I0(n27_adj_4369), .I1(n42302), .I2(n32), 
            .I3(n28_adj_4368), .O(n28_adj_4370));
    defparam i6_4_lut_adj_1273.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1274 (.I0(\data_out_frame[20] [5]), .I1(n42423), 
            .I2(n42173), .I3(\data_out_frame[20] [1]), .O(n35_adj_4371));
    defparam i13_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1275 (.I0(n37905), .I1(\data_out_frame[20] [2]), 
            .I2(n42305), .I3(n42146), .O(n34));
    defparam i12_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1276 (.I0(n35_adj_4371), .I1(n42058), .I2(n28_adj_4370), 
            .I3(n42194), .O(n40_adj_4372));
    defparam i18_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1277 (.I0(n42271), .I1(n42155), .I2(n42182), 
            .I3(n42026), .O(n38_adj_4373));
    defparam i16_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1278 (.I0(n42164), .I1(\data_out_frame[18] [5]), 
            .I2(n42019), .I3(n42321), .O(n37_adj_4374));
    defparam i15_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1279 (.I0(n37_adj_4374), .I1(n39_adj_4344), .I2(n38_adj_4373), 
            .I3(n40_adj_4372), .O(n42072));
    defparam i21_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1280 (.I0(n42277), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [1]), .I3(n6_adj_4274), .O(n41983));   // verilog/coms.v(69[16:62])
    defparam i4_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(n17289), .I1(n42378), .I2(\data_out_frame[14] [7]), 
            .I3(\data_out_frame[15] [1]), .O(n43449));
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1282 (.I0(n42072), .I1(\data_out_frame[17] [3]), 
            .I2(n43449), .I3(n42292), .O(n10_adj_4375));
    defparam i4_4_lut_adj_1282.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1283 (.I0(n41983), .I1(n10_adj_4375), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n43169));
    defparam i5_3_lut_adj_1283.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1284 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[13] [2]), .I3(GND_net), .O(n42109));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42155));
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1286 (.I0(n42109), .I1(n42314), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n17116));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42197));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1288 (.I0(\data_out_frame[19] [3]), .I1(n42197), 
            .I2(\data_out_frame[19] [4]), .I3(n38252), .O(n44072));
    defparam i3_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42302));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41925));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i3_2_lut (.I0(n42191), .I1(\data_out_frame[12] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n11));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1291 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[19] [1]), 
            .O(n13_adj_4376));
    defparam i5_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1292 (.I0(n13_adj_4376), .I1(n11), .I2(\data_out_frame[14] [7]), 
            .I3(n42092), .O(n44061));
    defparam i7_4_lut_adj_1292.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1293 (.I0(n17138), .I1(n42317), .I2(\data_out_frame[14] [2]), 
            .I3(GND_net), .O(n42009));
    defparam i2_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1294 (.I0(\data_out_frame[11] [6]), .I1(n16768), 
            .I2(n42210), .I3(n6_adj_4242), .O(n16815));
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1295 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[18] [7]), .I3(GND_net), .O(n42182));
    defparam i2_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1296 (.I0(n16815), .I1(n42009), .I2(n16989), 
            .I3(GND_net), .O(n1716));
    defparam i2_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_out_frame[18] [6]), .I1(n42354), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4377));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1298 (.I0(n1716), .I1(\data_out_frame[16] [4]), 
            .I2(n42182), .I3(n6_adj_4377), .O(n43377));
    defparam i4_4_lut_adj_1298.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16768));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1300 (.I0(n16768), .I1(n42039), .I2(\data_out_frame[12] [0]), 
            .I3(\data_out_frame[9] [6]), .O(n12_adj_4378));
    defparam i5_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1301 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[13] [7]), 
            .I2(n12_adj_4378), .I3(n8_adj_4379), .O(n42035));
    defparam i1_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17375));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\data_out_frame[14] [5]), .I1(n38226), 
            .I2(GND_net), .I3(GND_net), .O(n42161));
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1304 (.I0(\data_out_frame[19] [0]), .I1(n37473), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4380));
    defparam i2_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1305 (.I0(n7_adj_4380), .I1(n42259), .I2(n43760), 
            .I3(n42161), .O(n42354));
    defparam i4_4_lut_adj_1305.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16862));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42441));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4381));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1309 (.I0(n16873), .I1(\data_out_frame[9] [7]), 
            .I2(n42052), .I3(n6_adj_4381), .O(n41986));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_out_frame[12] [4]), .I1(n41986), 
            .I2(GND_net), .I3(GND_net), .O(n42259));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1311 (.I0(\data_out_frame[14] [5]), .I1(n42259), 
            .I2(\data_out_frame[16] [7]), .I3(n17142), .O(n42191));
    defparam i3_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1312 (.I0(n37575), .I1(n42441), .I2(n42225), 
            .I3(\data_out_frame[6] [3]), .O(n42378));
    defparam i3_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1313 (.I0(\data_out_frame[12] [7]), .I1(n16994), 
            .I2(\data_out_frame[15] [2]), .I3(\data_out_frame[11] [0]), 
            .O(n41971));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\data_out_frame[12] [6]), .I1(n41971), 
            .I2(GND_net), .I3(GND_net), .O(n17289));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(\data_out_frame[11] [1]), .I1(n1287), 
            .I2(n16862), .I3(n6_adj_4339), .O(n42314));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1316 (.I0(n41971), .I1(n42378), .I2(n42191), 
            .I3(n42176), .O(n38252));
    defparam i3_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42185));
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42176));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1319 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[8] [2]), .I3(n6_adj_4338), .O(n16994));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1320 (.I0(n16994), .I1(n37473), .I2(\data_out_frame[12] [5]), 
            .I3(GND_net), .O(n37575));
    defparam i2_3_lut_adj_1320.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1321 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[9] [3]), 
            .I2(n17004), .I3(n6_adj_4244), .O(n1379));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1322 (.I0(n42055), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[8] [4]), .I3(n6_adj_4243), .O(n17142));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_out_frame[11] [5]), .I1(n1379), 
            .I2(GND_net), .I3(GND_net), .O(n42112));
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1324 (.I0(n1185), .I1(n42210), .I2(n41895), .I3(n17198), 
            .O(n16253));
    defparam i3_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1325 (.I0(n42112), .I1(n17142), .I2(\data_out_frame[12] [7]), 
            .I3(n42417), .O(n10_adj_4382));
    defparam i4_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1326 (.I0(\data_out_frame[12] [6]), .I1(n10_adj_4382), 
            .I2(\data_out_frame[12] [4]), .I3(GND_net), .O(n43751));
    defparam i5_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1327 (.I0(n37575), .I1(n42112), .I2(\data_out_frame[13] [0]), 
            .I3(n43751), .O(n42426));
    defparam i3_4_lut_adj_1327.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1328 (.I0(n42426), .I1(n42324), .I2(n16253), 
            .I3(GND_net), .O(n37540));
    defparam i2_3_lut_adj_1328.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16691));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(n16893), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42023));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1331 (.I0(\data_in_frame[3] [7]), .I1(n41925), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[4] [1]), .O(n16889));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1332 (.I0(\data_out_frame[13] [3]), .I1(n16691), 
            .I2(\data_out_frame[13] [4]), .I3(n6_adj_4239), .O(n42324));
    defparam i4_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1333 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42055));
    defparam i1_2_lut_adj_1333.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1334 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42453));
    defparam i1_2_lut_adj_1334.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42317));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41919));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i395_2_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1185));   // verilog/coms.v(69[16:27])
    defparam i395_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1337 (.I0(\data_out_frame[10] [3]), .I1(n41965), 
            .I2(n41929), .I3(\data_out_frame[8] [2]), .O(n37473));   // verilog/coms.v(69[16:62])
    defparam i3_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i531_2_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1287));   // verilog/coms.v(69[16:27])
    defparam i531_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16873));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1339 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n41929));   // verilog/coms.v(69[16:62])
    defparam i2_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1340 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[6] [4]), .O(n41980));
    defparam i3_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17424));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1342 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [3]), .I3(n1379), .O(n8_adj_4379));
    defparam i1_2_lut_3_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1343 (.I0(n16889), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[8] [6]), .I3(n42023), .O(n41974));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n41938));
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_LUT4 i12_3_lut_4_lut_adj_1345 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(n42342), .I3(n16938), .O(n29));
    defparam i12_3_lut_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1346 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[14]_c [2]), .I3(\data_in_frame[14] [1]), 
            .O(n18_adj_4211));
    defparam i1_2_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1347 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [5]), .I3(n6_adj_4240), .O(n41895));
    defparam i4_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1348 (.I0(n41938), .I1(\data_out_frame[7] [6]), 
            .I2(n42283), .I3(n17424), .O(n30_adj_4383));
    defparam i11_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1349 (.I0(\data_out_frame[11] [4]), .I1(n30_adj_4383), 
            .I2(n16778), .I3(\data_out_frame[9] [0]), .O(n34_adj_4384));
    defparam i15_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1350 (.I0(n42339), .I1(n41980), .I2(n42039), 
            .I3(n41929), .O(n32_adj_4385));
    defparam i13_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1351 (.I0(n1185), .I1(n34_adj_4384), .I2(n28_adj_4245), 
            .I3(\data_out_frame[10] [4]), .O(n36_adj_4386));
    defparam i17_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1352 (.I0(n42032), .I1(\data_out_frame[9] [1]), 
            .I2(n41919), .I3(n37697), .O(n31_adj_4387));
    defparam i12_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1353 (.I0(n42317), .I1(n31_adj_4387), .I2(n36_adj_4386), 
            .I3(n32_adj_4385), .O(n42417));
    defparam i2_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1354 (.I0(\data_out_frame[6] [4]), .I1(n42456), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4388));
    defparam i4_2_lut_adj_1354.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1355 (.I0(n42417), .I1(n41895), .I2(n42241), 
            .I3(\data_out_frame[5] [2]), .O(n24_adj_4389));
    defparam i10_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1356 (.I0(n42453), .I1(n42055), .I2(\data_out_frame[6] [3]), 
            .I3(\data_out_frame[7] [0]), .O(n22_adj_4390));
    defparam i8_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1357 (.I0(n42324), .I1(n24_adj_4389), .I2(n18_adj_4388), 
            .I3(\data_out_frame[7] [3]), .O(n26_adj_4391));
    defparam i12_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i13062_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n18346));
    defparam i13062_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1358 (.I0(\data_out_frame[8] [5]), .I1(n26_adj_4391), 
            .I2(n22_adj_4390), .I3(n37540), .O(n37409));
    defparam i13_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1359 (.I0(\data_out_frame[10] [5]), .I1(n42241), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n42387));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4241));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1361 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(n17206), .I3(\data_out_frame[10] [1]), .O(n42052));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1362 (.I0(n42052), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4392));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1363 (.I0(n42280), .I1(\data_out_frame[12] [1]), 
            .I2(n41946), .I3(\data_out_frame[12] [2]), .O(n14_adj_4393));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1364 (.I0(\data_out_frame[14] [3]), .I1(n14_adj_4393), 
            .I2(n10_adj_4392), .I3(\data_out_frame[5] [1]), .O(n16989));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42194));
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1366 (.I0(\data_out_frame[12] [4]), .I1(n42203), 
            .I2(n37575), .I3(GND_net), .O(n37877));
    defparam i2_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1367 (.I0(n37877), .I1(n38226), .I2(n42194), 
            .I3(\data_out_frame[16] [6]), .O(n42091));
    defparam i3_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1368 (.I0(n16989), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4394));   // verilog/coms.v(72[16:27])
    defparam i4_2_lut_adj_1368.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1369 (.I0(n38226), .I1(n42387), .I2(n37409), 
            .I3(\data_out_frame[11] [1]), .O(n24_adj_4395));   // verilog/coms.v(72[16:27])
    defparam i10_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1370 (.I0(\data_out_frame[13] [1]), .I1(n41919), 
            .I2(n42185), .I3(\data_out_frame[16] [5]), .O(n22_adj_4396));   // verilog/coms.v(72[16:27])
    defparam i8_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i13063_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n18347));
    defparam i13063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1371 (.I0(n38252), .I1(n24_adj_4395), .I2(n18_adj_4394), 
            .I3(n42314), .O(n26_adj_4397));   // verilog/coms.v(72[16:27])
    defparam i12_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1372 (.I0(n41952), .I1(n26_adj_4397), .I2(n22_adj_4396), 
            .I3(\data_out_frame[8] [7]), .O(n43760));   // verilog/coms.v(72[16:27])
    defparam i13_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(n43760), .I1(n42091), .I2(GND_net), 
            .I3(GND_net), .O(n42092));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1374 (.I0(\data_out_frame[16] [5]), .I1(n37877), 
            .I2(n42354), .I3(\data_out_frame[20] [7]), .O(n12_adj_4398));   // verilog/coms.v(69[16:62])
    defparam i5_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1375 (.I0(n17375), .I1(n12_adj_4398), .I2(n42185), 
            .I3(\data_out_frame[16] [7]), .O(n42146));   // verilog/coms.v(69[16:62])
    defparam i6_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i13064_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n18348));
    defparam i13064_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1376 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41946));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1376.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1377 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17206));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1377.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1378 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4399));   // verilog/coms.v(69[16:62])
    defparam i2_2_lut_adj_1378.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1379 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [6]), .I3(n41965), .O(n14_adj_4400));   // verilog/coms.v(69[16:62])
    defparam i6_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1380 (.I0(\data_out_frame[5] [6]), .I1(n14_adj_4400), 
            .I2(n10_adj_4399), .I3(\data_out_frame[6] [0]), .O(n42049));   // verilog/coms.v(69[16:62])
    defparam i7_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1381 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[10] [0]), .I3(n41946), .O(n10_adj_4332));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1382 (.I0(n16772), .I1(n10_adj_4332), .I2(\data_out_frame[5] [5]), 
            .I3(GND_net), .O(n17138));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16778));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1384 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n17198));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1385 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n16772));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42029));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1387 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [4]), 
            .I2(n42029), .I3(\data_out_frame[9] [5]), .O(n42032));
    defparam i3_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1388 (.I0(\data_out_frame[11] [4]), .I1(n17198), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n17430));
    defparam i2_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1389 (.I0(n17430), .I1(\data_out_frame[5] [0]), 
            .I2(n42032), .I3(n6_adj_4331), .O(n37471));
    defparam i4_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1390 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[18] [4]), 
            .I2(n37471), .I3(GND_net), .O(n42058));
    defparam i2_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42164));
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1392 (.I0(\data_out_frame[14] [4]), .I1(n16778), 
            .I2(\data_out_frame[10] [2]), .I3(n37697), .O(n38226));
    defparam i3_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1393 (.I0(n38226), .I1(\data_out_frame[20] [7]), 
            .I2(n42164), .I3(n6_adj_4237), .O(n43355));
    defparam i4_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i13065_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n18349));
    defparam i13065_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_41972 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4322), .I2(n46584), .I3(byte_transmit_counter_c[2]), 
            .O(n49883));
    defparam byte_transmit_counter_1__bdd_4_lut_41972.LUT_INIT = 16'he4aa;
    SB_LUT4 i13066_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n18350));
    defparam i13066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49883_bdd_4_lut (.I0(n49883), .I1(n17_adj_4321), .I2(n16_adj_4320), 
            .I3(byte_transmit_counter_c[2]), .O(n49886));
    defparam n49883_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1394 (.I0(\data_in_frame[6] [1]), .I1(n42131), 
            .I2(n16938), .I3(n16889), .O(n12_adj_4401));   // verilog/coms.v(73[16:43])
    defparam i5_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_41967 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4319), .I2(n46583), .I3(byte_transmit_counter_c[2]), 
            .O(n49877));
    defparam byte_transmit_counter_1__bdd_4_lut_41967.LUT_INIT = 16'he4aa;
    SB_LUT4 n49877_bdd_4_lut (.I0(n49877), .I1(n17_adj_4318), .I2(n16_adj_4317), 
            .I3(byte_transmit_counter_c[2]), .O(n49880));
    defparam n49877_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1395 (.I0(\data_in_frame[8] [6]), .I1(n12_adj_4401), 
            .I2(n42336), .I3(n17126), .O(Kp_23__N_1201));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_41962 (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_4316), .I2(n46582), .I3(byte_transmit_counter_c[2]), 
            .O(n49871));
    defparam byte_transmit_counter_1__bdd_4_lut_41962.LUT_INIT = 16'he4aa;
    SB_LUT4 n49871_bdd_4_lut (.I0(n49871), .I1(n17_adj_4315), .I2(n16_adj_4314), 
            .I3(byte_transmit_counter_c[2]), .O(n49874));
    defparam n49871_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1396 (.I0(n42327), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[8] [5]), .I3(n42396), .O(n10_adj_4402));   // verilog/coms.v(77[16:35])
    defparam i4_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i13067_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n18351));
    defparam i13067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13068_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n18352));
    defparam i13068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1397 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n16446), .I3(n16682), .O(n16683));   // verilog/coms.v(148[5:9])
    defparam i1_2_lut_3_lut_4_lut_adj_1397.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n16446), .I3(n16675), .O(n16676));   // verilog/coms.v(148[5:9])
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1399 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n16446), .I3(\FRAME_MATCHER.state [2]), 
            .O(n16679));   // verilog/coms.v(148[5:9])
    defparam i1_2_lut_3_lut_4_lut_adj_1399.LUT_INIT = 16'hfeff;
    SB_LUT4 i13069_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41852), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n18353));
    defparam i13069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8691_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n13947));
    defparam i8691_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i13030_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n18314));
    defparam i13030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(\data_in_frame[5] [0]), .I1(n17037), 
            .I2(n41956), .I3(GND_net), .O(n1));
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_LUT4 i13150_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n18434));
    defparam i13150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13031_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n18315));
    defparam i13031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13151_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n18435));
    defparam i13151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1401 (.I0(n41974), .I1(n10_adj_4402), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(Kp_23__N_1213));   // verilog/coms.v(77[16:35])
    defparam i5_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_42017 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49859));
    defparam byte_transmit_counter_0__bdd_4_lut_42017.LUT_INIT = 16'he4aa;
    SB_LUT4 i13032_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n18316));
    defparam i13032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13033_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n18317));
    defparam i13033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49859_bdd_4_lut (.I0(n49859), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49862));
    defparam n49859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41948 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49853));
    defparam byte_transmit_counter_0__bdd_4_lut_41948.LUT_INIT = 16'he4aa;
    SB_LUT4 n49853_bdd_4_lut (.I0(n49853), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49856));
    defparam n49853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_1402 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[14] [5]), 
            .I2(n4), .I3(\data_in_frame[16] [7]), .O(n42311));
    defparam i2_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41943 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49847));
    defparam byte_transmit_counter_0__bdd_4_lut_41943.LUT_INIT = 16'he4aa;
    SB_LUT4 n49847_bdd_4_lut (.I0(n49847), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49850));
    defparam n49847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41938 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49841));
    defparam byte_transmit_counter_0__bdd_4_lut_41938.LUT_INIT = 16'he4aa;
    SB_LUT4 n49841_bdd_4_lut (.I0(n49841), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49844));
    defparam n49841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1403 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[14] [6]), .I3(GND_net), .O(n42103));
    defparam i2_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41933 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49835));
    defparam byte_transmit_counter_0__bdd_4_lut_41933.LUT_INIT = 16'he4aa;
    SB_LUT4 n49835_bdd_4_lut (.I0(n49835), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n49838));
    defparam n49835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_2_lut_adj_1404 (.I0(n42438), .I1(n41974), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4404));   // verilog/coms.v(73[16:43])
    defparam i3_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1405 (.I0(\data_in_frame[11] [0]), .I1(n42381), 
            .I2(n42462), .I3(n42103), .O(n22_adj_4405));   // verilog/coms.v(73[16:43])
    defparam i9_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41928 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49823));
    defparam byte_transmit_counter_0__bdd_4_lut_41928.LUT_INIT = 16'he4aa;
    SB_LUT4 i13034_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n18318));
    defparam i13034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1406 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(n6_adj_4130), .O(Kp_23__N_676));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1407 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n41891));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i13035_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n18319));
    defparam i13035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_809));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i13036_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n18320));
    defparam i13036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49823_bdd_4_lut (.I0(n49823), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n49826));
    defparam n49823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20048_2_lut (.I0(n31_adj_4140), .I1(n25297), .I2(GND_net), 
            .I3(GND_net), .O(n25307));
    defparam i20048_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1409 (.I0(n16680), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n44325), .O(n25611));
    defparam i2_3_lut_4_lut_adj_1409.LUT_INIT = 16'haa8a;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n16563), .I3(\FRAME_MATCHER.state [2]), .O(n16680));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'hfdff;
    SB_LUT4 i13037_3_lut_4_lut (.I0(n8_adj_4137), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n18321));
    defparam i13037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13129_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n18413));
    defparam i13129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13130_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n18414));
    defparam i13130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13131_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18415));
    defparam i13131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13132_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18416));
    defparam i13132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_adj_1411 (.I0(n16938), .I1(\data_in_frame[19] [4]), 
            .I2(n42268), .I3(GND_net), .O(n20_adj_4406));   // verilog/coms.v(73[16:43])
    defparam i7_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i13128_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n18412));
    defparam i13128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13133_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18417));
    defparam i13133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1412 (.I0(\data_in_frame[13] [1]), .I1(n22_adj_4405), 
            .I2(n16_adj_4404), .I3(n19), .O(n24_adj_4408));   // verilog/coms.v(73[16:43])
    defparam i11_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_41919 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49817));
    defparam byte_transmit_counter_0__bdd_4_lut_41919.LUT_INIT = 16'he4aa;
    SB_LUT4 n49817_bdd_4_lut (.I0(n49817), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n49820));
    defparam n49817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13126_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n18410));
    defparam i13126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13152_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n18436));
    defparam i13152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1413 (.I0(\data_in_frame[17] [3]), .I1(n24_adj_4408), 
            .I2(n20_adj_4406), .I3(n17185), .O(n42248));   // verilog/coms.v(73[16:43])
    defparam i12_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1414 (.I0(n42103), .I1(\data_in_frame[17] [1]), 
            .I2(n42393), .I3(n42311), .O(n10_adj_4409));   // verilog/coms.v(71[16:42])
    defparam i4_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i13127_3_lut_4_lut (.I0(n8_adj_4123), .I1(n41861), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n18411));
    defparam i13127_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13118_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n18402));
    defparam i13118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13119_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n18403));
    defparam i13119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13120_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n18404));
    defparam i13120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13121_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n18405));
    defparam i13121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13122_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n18406));
    defparam i13122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1415 (.I0(\data_in_frame[19] [3]), .I1(Kp_23__N_1213), 
            .I2(n10_adj_4409), .I3(Kp_23__N_1201), .O(n41959));
    defparam i1_4_lut_adj_1415.LUT_INIT = 16'h9669;
    SB_LUT4 i13153_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n18437));
    defparam i13153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1416 (.I0(n47), .I1(n26154), .I2(n4_adj_4329), 
            .I3(n13980), .O(n3735));
    defparam i1_4_lut_adj_1416.LUT_INIT = 16'h3032;
    SB_LUT4 i13123_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n18407));
    defparam i13123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13124_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n18408));
    defparam i13124_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1417 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [1]), .O(n14_adj_4410));
    defparam i6_4_lut_adj_1417.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1418 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[2] [2]), .O(n13_adj_4411));
    defparam i5_4_lut_adj_1418.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1419 (.I0(\data_in_frame[1] [5]), .I1(n13_adj_4411), 
            .I2(n14_adj_4410), .I3(GND_net), .O(n22_adj_4412));
    defparam i5_3_lut_adj_1419.LUT_INIT = 16'h0202;
    SB_LUT4 i10_4_lut_adj_1420 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [0]), .O(n27_adj_4413));
    defparam i10_4_lut_adj_1420.LUT_INIT = 16'h4000;
    SB_LUT4 i9_3_lut_adj_1421 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [7]), .I3(GND_net), .O(n26_adj_4414));
    defparam i9_3_lut_adj_1421.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_4_lut_adj_1422 (.I0(\data_in_frame[3] [2]), .I1(n15066), 
            .I2(\data_in_frame[5] [4]), .I3(n41891), .O(n17185));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i36340_2_lut (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44231));
    defparam i36340_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i36404_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[0] [2]), .O(n44302));
    defparam i36404_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1423 (.I0(n27_adj_4413), .I1(\data_in_frame[2] [1]), 
            .I2(n22_adj_4412), .I3(\data_in_frame[1] [4]), .O(n31_adj_4415));
    defparam i14_4_lut_adj_1423.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_1424 (.I0(n31_adj_4415), .I1(n44302), .I2(n44231), 
            .I3(n26_adj_4414), .O(\FRAME_MATCHER.state_31__N_2275 [3]));
    defparam i16_4_lut_adj_1424.LUT_INIT = 16'h0200;
    SB_LUT4 i13125_3_lut_4_lut (.I0(n8), .I1(n41861), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n18409));
    defparam i13125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [14]), 
            .I2(GND_net), .I3(GND_net), .O(n144));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1426 (.I0(\FRAME_MATCHER.state [12]), .I1(\FRAME_MATCHER.state [10]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [8]), 
            .O(n10));
    defparam i4_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\data_in_frame[3] [2]), .I1(n15066), 
            .I2(\data_in_frame[3] [1]), .I3(GND_net), .O(n4_adj_4131));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i13022_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n18306));
    defparam i13022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18425_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(\data_in_frame[5] [1]), 
            .I3(rx_data[1]), .O(n18307));
    defparam i18425_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13024_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n18308));
    defparam i13024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13025_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n18309));
    defparam i13025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13026_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n18310));
    defparam i13026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13029_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n18313));
    defparam i13029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13028_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n18312));
    defparam i13028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13027_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n18311));
    defparam i13027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13110_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18394));
    defparam i13110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13111_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18395));
    defparam i13111_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13112_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18396));
    defparam i13112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13113_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18397));
    defparam i13113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13114_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18398));
    defparam i13114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13115_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18399));
    defparam i13115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13116_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18400));
    defparam i13116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13117_3_lut_4_lut (.I0(n8_adj_4227), .I1(n41861), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18401));
    defparam i13117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13006_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n18290));
    defparam i13006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13007_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n18291));
    defparam i13007_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13008_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n18292));
    defparam i13008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13009_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n18293));
    defparam i13009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13010_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n18294));
    defparam i13010_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13011_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n18295));
    defparam i13011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13012_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n18296));
    defparam i13012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13154_3_lut_4_lut (.I0(n8_adj_4127), .I1(n41861), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n18438));
    defparam i13154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13013_3_lut_4_lut (.I0(n8_adj_4116), .I1(n41843), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n18297));
    defparam i13013_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.n41336(n41336), .clk32MHz(clk32MHz), .n41446(n41446), 
            .n41444(n41444), .n41442(n41442), .n41074(n41074), .\r_Clock_Count[8] (\r_Clock_Count[8] ), 
            .n41130(n41130), .\r_Clock_Count[7] (\r_Clock_Count[7] ), .n41224(n41224), 
            .\r_Clock_Count[6] (\r_Clock_Count[6] ), .r_SM_Main({Open_10, 
            r_SM_Main_c[1], Open_11}), .VCC_net(VCC_net), .n41348(n41348), 
            .tx_data({tx_data}), .tx_o(tx_o), .tx_enable(tx_enable), .GND_net(GND_net), 
            .n88(n88), .n118(n118), .\r_SM_Main[2] (\r_SM_Main[2] ), .n5(n5_adj_16), 
            .n44294(n44294), .n17955(n17955), .n17977(n17977), .n17980(n17980), 
            .n17863(n17863), .n17866(n17866), .n17869(n17869), .n17872(n17872), 
            .n18575(n18575), .n41424(n41424), .tx_active(tx_active), .n17974(n17974), 
            .\r_SM_Main_2__N_3106[0] (r_SM_Main_2__N_3106[0]), .n19921(n19921), 
            .n3(n3_adj_17), .n10142(n10142), .n4(n4_adj_4326)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.n17887(n17887), .r_Bit_Index({r_Bit_Index}), .clk32MHz(clk32MHz), 
            .n17890(n17890), .n18701(n18701), .VCC_net(VCC_net), .r_Clock_Count({Open_12, 
            Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, 
            \r_Clock_Count[0] }), .r_SM_Main({r_SM_Main}), .n18587(n18587), 
            .rx_data({rx_data}), .n41150(n41150), .rx_data_ready(rx_data_ready), 
            .n18583(n18583), .n18567(n18567), .\r_Clock_Count[5] (\r_Clock_Count[5] ), 
            .n18555(n18555), .\r_Clock_Count[1] (\r_Clock_Count[1] ), .\r_SM_Main_2__N_3032[2] (\r_SM_Main_2__N_3032[2] ), 
            .r_Rx_Data(r_Rx_Data), .PIN_13_N_50(PIN_13_N_50), .GND_net(GND_net), 
            .n27708(n27708), .n17657(n17657), .n17707(n17707), .n17849(n17849), 
            .n4694(n4694), .n221(n221), .n225(n225), .n226(n226), .n17897(n17897), 
            .n17896(n17896), .n17895(n17895), .n17894(n17894), .n17893(n17893), 
            .n17892(n17892), .n17891(n17891), .n16566(n16566), .n4(n4_adj_19), 
            .n25329(n25329), .n4_adj_13(n4_adj_20), .n4_adj_14(n4_adj_21), 
            .n16432(n16432)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n41336, clk32MHz, n41446, n41444, n41442, n41074, 
            \r_Clock_Count[8] , n41130, \r_Clock_Count[7] , n41224, 
            \r_Clock_Count[6] , r_SM_Main, VCC_net, n41348, tx_data, 
            tx_o, tx_enable, GND_net, n88, n118, \r_SM_Main[2] , 
            n5, n44294, n17955, n17977, n17980, n17863, n17866, 
            n17869, n17872, n18575, n41424, tx_active, n17974, \r_SM_Main_2__N_3106[0] , 
            n19921, n3, n10142, n4) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n41336;
    input clk32MHz;
    input n41446;
    input n41444;
    input n41442;
    input n41074;
    output \r_Clock_Count[8] ;
    input n41130;
    output \r_Clock_Count[7] ;
    input n41224;
    output \r_Clock_Count[6] ;
    output [2:0]r_SM_Main;
    input VCC_net;
    input n41348;
    input [7:0]tx_data;
    output tx_o;
    output tx_enable;
    input GND_net;
    output n88;
    output n118;
    output \r_SM_Main[2] ;
    input n5;
    output n44294;
    output n17955;
    output n17977;
    output n17980;
    output n17863;
    output n17866;
    output n17869;
    output n17872;
    output n18575;
    input n41424;
    output tx_active;
    input n17974;
    input \r_SM_Main_2__N_3106[0] ;
    output n19921;
    output n3;
    output n10142;
    output n4;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n41370, n17881;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n17884, n18621, n41368, n14181;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n27954, n17713, n41702, n27876, n109;
    wire [2:0]r_SM_Main_c;   // verilog/uart_tx.v(31[16:25])
    
    wire n36995, n37, n34599, n34598, n34597, n34596, n34595, 
        n34594, n34593, n34592, n17976, n50335, n49919, n49922, 
        n49814, o_Tx_Serial_N_3134, n12493, n49811;
    
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n41336));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n41446));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n41444));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n41442));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n41370));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17881));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17884));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(\r_Clock_Count[8] ), .C(clk32MHz), .D(n41074));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(\r_Clock_Count[7] ), .C(clk32MHz), .D(n41130));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(clk32MHz), .D(n41224));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n18621));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n41368));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n41348));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut (.I0(n27954), .I1(r_Bit_Index[1]), .I2(n17713), .I3(r_Bit_Index[0]), 
            .O(n17884));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut.LUT_INIT = 16'h2888;
    SB_LUT4 i2_3_lut (.I0(n88), .I1(n41702), .I2(n118), .I3(GND_net), 
            .O(n27876));   // verilog/uart_tx.v(32[16:29])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_879 (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n109));
    defparam i2_3_lut_adj_879.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_c[0]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(n27876), .O(n17713));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut (.I0(r_SM_Main[1]), .I1(n17713), .I2(n109), .I3(GND_net), 
            .O(n27954));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut.LUT_INIT = 16'h3b3b;
    SB_LUT4 i29122_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n36995));   // verilog/uart_tx.v(33[16:27])
    defparam i29122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_880 (.I0(n27954), .I1(r_Bit_Index[2]), .I2(n17713), 
            .I3(n36995), .O(n17881));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_880.LUT_INIT = 16'h2888;
    SB_LUT4 i1_2_lut (.I0(n37), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n41370));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_881 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), 
            .I2(GND_net), .I3(GND_net), .O(n118));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_881.LUT_INIT = 16'heeee;
    SB_LUT4 i36398_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44294));
    defparam i36398_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[2]), 
            .I3(r_Clock_Count[1]), .O(n88));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_adj_882 (.I0(\r_Clock_Count[7] ), .I1(\r_Clock_Count[6] ), 
            .I2(\r_Clock_Count[8] ), .I3(GND_net), .O(n41702));
    defparam i2_3_lut_adj_882.LUT_INIT = 16'hfefe;
    SB_LUT4 add_59_10_lut (.I0(\r_Clock_Count[8] ), .I1(\r_Clock_Count[8] ), 
            .I2(\r_SM_Main[2] ), .I3(n34599), .O(n17955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_59_9_lut (.I0(\r_Clock_Count[7] ), .I1(\r_Clock_Count[7] ), 
            .I2(\r_SM_Main[2] ), .I3(n34598), .O(n17977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_9 (.CI(n34598), .I0(\r_Clock_Count[7] ), .I1(\r_SM_Main[2] ), 
            .CO(n34599));
    SB_LUT4 add_59_8_lut (.I0(\r_Clock_Count[6] ), .I1(\r_Clock_Count[6] ), 
            .I2(\r_SM_Main[2] ), .I3(n34597), .O(n17980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_8 (.CI(n34597), .I0(\r_Clock_Count[6] ), .I1(\r_SM_Main[2] ), 
            .CO(n34598));
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n14181), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(\r_SM_Main[2] ), .I3(n34596), .O(n17863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n34596), .I0(r_Clock_Count[5]), .I1(\r_SM_Main[2] ), 
            .CO(n34597));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(\r_SM_Main[2] ), .I3(n34595), .O(n17866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n34595), .I0(r_Clock_Count[4]), .I1(\r_SM_Main[2] ), 
            .CO(n34596));
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(\r_SM_Main[2] ), .I3(n34594), .O(n17869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_5 (.CI(n34594), .I0(r_Clock_Count[3]), .I1(\r_SM_Main[2] ), 
            .CO(n34595));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(\r_SM_Main[2] ), .I3(n34593), .O(n17872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n34593), .I0(r_Clock_Count[2]), .I1(\r_SM_Main[2] ), 
            .CO(n34594));
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(\r_SM_Main[2] ), .I3(n34592), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n34592), .I0(r_Clock_Count[1]), .I1(\r_SM_Main[2] ), 
            .CO(n34593));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(\r_SM_Main[2] ), .I3(VCC_net), .O(n18575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(\r_SM_Main[2] ), 
            .CO(n34592));
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n17976));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n41424));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n17974));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(n50335));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n49919));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49919_bdd_4_lut (.I0(n49919), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n49922));
    defparam n49919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_883 (.I0(tx_active), .I1(\r_SM_Main_2__N_3106[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n19921));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_883.LUT_INIT = 16'heeee;
    SB_LUT4 i12_3_lut (.I0(n17713), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n41368));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i3_4_lut_adj_884 (.I0(r_SM_Main[1]), .I1(n27876), .I2(\r_SM_Main[2] ), 
            .I3(r_SM_Main_c[0]), .O(n50335));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_adj_884.LUT_INIT = 16'h0800;
    SB_LUT4 i20933221_i1_3_lut (.I0(n49922), .I1(n49814), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3134));
    defparam i20933221_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main_c[0]), .I1(o_Tx_Serial_N_3134), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i5126_2_lut (.I0(\r_SM_Main_2__N_3106[0] ), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n10142));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5126_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7361_4_lut (.I0(\r_SM_Main_2__N_3106[0] ), .I1(n109), .I2(r_SM_Main[1]), 
            .I3(n27876), .O(n12493));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7361_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_885 (.I0(\r_SM_Main[2] ), .I1(n12493), .I2(n27876), 
            .I3(r_SM_Main_c[0]), .O(n17976));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_885.LUT_INIT = 16'h0544;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(n27876), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main[2] ), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i1_3_lut_4_lut_adj_886 (.I0(r_SM_Main_c[0]), .I1(n27876), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main[2] ), .O(n18621));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut_adj_886.LUT_INIT = 16'h0078;
    SB_LUT4 i3_3_lut_4_lut (.I0(\r_SM_Main_2__N_3106[0] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main_c[0]), .I3(\r_SM_Main[2] ), .O(n14181));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_41997 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n49811));
    defparam r_Bit_Index_0__bdd_4_lut_41997.LUT_INIT = 16'he4aa;
    SB_LUT4 n49811_bdd_4_lut (.I0(n49811), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n49814));
    defparam n49811_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n17887, r_Bit_Index, clk32MHz, n17890, n18701, VCC_net, 
            r_Clock_Count, r_SM_Main, n18587, rx_data, n41150, rx_data_ready, 
            n18583, n18567, \r_Clock_Count[5] , n18555, \r_Clock_Count[1] , 
            \r_SM_Main_2__N_3032[2] , r_Rx_Data, PIN_13_N_50, GND_net, 
            n27708, n17657, n17707, n17849, n4694, n221, n225, 
            n226, n17897, n17896, n17895, n17894, n17893, n17892, 
            n17891, n16566, n4, n25329, n4_adj_13, n4_adj_14, n16432) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17887;
    output [2:0]r_Bit_Index;
    input clk32MHz;
    input n17890;
    input n18701;
    input VCC_net;
    output [7:0]r_Clock_Count;
    output [2:0]r_SM_Main;
    input n18587;
    output [7:0]rx_data;
    input n41150;
    output rx_data_ready;
    input n18583;
    input n18567;
    output \r_Clock_Count[5] ;
    input n18555;
    output \r_Clock_Count[1] ;
    output \r_SM_Main_2__N_3032[2] ;
    output r_Rx_Data;
    input PIN_13_N_50;
    input GND_net;
    output n27708;
    output n17657;
    output n17707;
    output n17849;
    output n4694;
    output n221;
    output n225;
    output n226;
    input n17897;
    input n17896;
    input n17895;
    input n17894;
    input n17893;
    input n17892;
    input n17891;
    output n16566;
    output n4;
    output n25329;
    output n4_adj_13;
    output n4_adj_14;
    output n16432;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n26084, n18573;
    wire [7:0]r_Clock_Count_c;   // verilog/uart_rx.v(32[17:30])
    
    wire n18570, n18564, n18561, n18558, n41870, r_Rx_Data_R, n144, 
        n6, n129, n81, n85, n76, n119, n131, n10, n44243, 
        n25923, n49979, n49982, n46622, n34591, n138;
    wire [31:0]n194;
    
    wire n34590, n34589, n46491, n34588, n46621, n34587, n34586, 
        n34585, n26082, n46619, n16437, n46620, n77, n43440;
    
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17887));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17890));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18701));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n26084));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18587));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n41150));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18583));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i7 (.Q(r_Clock_Count_c[7]), .C(clk32MHz), .E(VCC_net), 
            .D(n18573));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i6 (.Q(r_Clock_Count_c[6]), .C(clk32MHz), .E(VCC_net), 
            .D(n18570));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i5 (.Q(\r_Clock_Count[5] ), .C(clk32MHz), .E(VCC_net), 
            .D(n18567));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i4 (.Q(r_Clock_Count_c[4]), .C(clk32MHz), .E(VCC_net), 
            .D(n18564));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i3 (.Q(r_Clock_Count_c[3]), .C(clk32MHz), .E(VCC_net), 
            .D(n18561));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i2 (.Q(r_Clock_Count_c[2]), .C(clk32MHz), .E(VCC_net), 
            .D(n18558));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i1 (.Q(\r_Clock_Count[1] ), .C(clk32MHz), .E(VCC_net), 
            .D(n18555));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3032[2] ), 
            .R(n41870));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_50));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i147_2_lut (.I0(r_Clock_Count_c[4]), .I1(r_Clock_Count_c[7]), 
            .I2(GND_net), .I3(GND_net), .O(n144));
    defparam i147_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(\r_Clock_Count[1] ), .I1(r_Clock_Count_c[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut (.I0(n129), .I1(n81), .I2(n144), .I3(n6), .O(n85));
    defparam i4_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[0]), .I1(n85), .I2(r_Rx_Data), .I3(r_SM_Main[1]), 
            .O(n76));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut.LUT_INIT = 16'h22a2;
    SB_LUT4 i2_3_lut (.I0(r_Clock_Count_c[3]), .I1(r_SM_Main[0]), .I2(n119), 
            .I3(GND_net), .O(n131));
    defparam i2_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i4_4_lut_adj_868 (.I0(\r_Clock_Count[1] ), .I1(r_SM_Main[1]), 
            .I2(n131), .I3(r_Clock_Count_c[2]), .O(n10));
    defparam i4_4_lut_adj_868.LUT_INIT = 16'hfdff;
    SB_LUT4 i36352_2_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44243));
    defparam i36352_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_869 (.I0(r_SM_Main[2]), .I1(n27708), .I2(n44243), 
            .I3(n10), .O(n17657));
    defparam i1_4_lut_adj_869.LUT_INIT = 16'h7737;
    SB_LUT4 i1_4_lut_adj_870 (.I0(r_SM_Main[2]), .I1(n76), .I2(\r_SM_Main_2__N_3032[2] ), 
            .I3(r_SM_Main[1]), .O(n27708));   // verilog/uart_rx.v(36[17:26])
    defparam i1_4_lut_adj_870.LUT_INIT = 16'hafee;
    SB_LUT4 i1_2_lut_adj_871 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n81));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_872 (.I0(r_Clock_Count_c[6]), .I1(\r_Clock_Count[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n129));
    defparam i1_2_lut_adj_872.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_873 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n25923));
    defparam i2_3_lut_adj_873.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3032[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n17707));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i12565_3_lut (.I0(n17707), .I1(n25923), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17849));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12565_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1266_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4694));   // verilog/uart_rx.v(102[36:51])
    defparam i1266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n49979_bdd_4_lut (.I0(n49979), .I1(n85), .I2(r_Rx_Data), .I3(r_SM_Main[1]), 
            .O(n49982));
    defparam n49979_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_62_9_lut (.I0(n138), .I1(r_Clock_Count_c[7]), .I2(GND_net), 
            .I3(n34591), .O(n46622)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count_c[6]), .I2(GND_net), 
            .I3(n34590), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n34590), .I0(r_Clock_Count_c[6]), .I1(GND_net), 
            .CO(n34591));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(\r_Clock_Count[5] ), .I2(GND_net), 
            .I3(n34589), .O(n221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n34589), .I0(\r_Clock_Count[5] ), .I1(GND_net), 
            .CO(n34590));
    SB_LUT4 add_62_6_lut (.I0(n138), .I1(r_Clock_Count_c[4]), .I2(GND_net), 
            .I3(n34588), .O(n46491)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n34588), .I0(r_Clock_Count_c[4]), .I1(GND_net), 
            .CO(n34589));
    SB_LUT4 add_62_5_lut (.I0(n138), .I1(r_Clock_Count_c[3]), .I2(GND_net), 
            .I3(n34587), .O(n46621)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n34587), .I0(r_Clock_Count_c[3]), .I1(GND_net), 
            .CO(n34588));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count_c[2]), .I2(GND_net), 
            .I3(n34586), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n34586), .I0(r_Clock_Count_c[2]), .I1(GND_net), 
            .CO(n34587));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(\r_Clock_Count[1] ), .I2(GND_net), 
            .I3(n34585), .O(n225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n34585), .I0(\r_Clock_Count[1] ), .I1(GND_net), 
            .CO(n34586));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n34585));
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n26082));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17897));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17896));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17895));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17894));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17893));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17892));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17891));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i38930_3_lut_4_lut (.I0(\r_Clock_Count[1] ), .I1(n81), .I2(r_Rx_Data), 
            .I3(n131), .O(n46619));
    defparam i38930_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_4_lut_adj_874 (.I0(n27708), .I1(r_Clock_Count_c[2]), .I2(n194[2]), 
            .I3(n17657), .O(n18558));
    defparam i1_4_lut_adj_874.LUT_INIT = 16'ha088;
    SB_LUT4 i22525_3_lut (.I0(r_Clock_Count_c[3]), .I1(n46621), .I2(n17657), 
            .I3(GND_net), .O(n18561));
    defparam i22525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22579_3_lut (.I0(r_Clock_Count_c[4]), .I1(n46491), .I2(n17657), 
            .I3(GND_net), .O(n18564));
    defparam i22579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_875 (.I0(n27708), .I1(r_Clock_Count_c[6]), .I2(n194[6]), 
            .I3(n17657), .O(n18570));
    defparam i1_4_lut_adj_875.LUT_INIT = 16'ha088;
    SB_LUT4 i22552_3_lut (.I0(r_Clock_Count_c[7]), .I1(n46622), .I2(n17657), 
            .I3(GND_net), .O(n18573));
    defparam i22552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_876 (.I0(r_Bit_Index[0]), .I1(n16437), .I2(GND_net), 
            .I3(GND_net), .O(n16566));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_876.LUT_INIT = 16'heeee;
    SB_LUT4 equal_85_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_85_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i39441_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3032[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n46620));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i39441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i41193_4_lut (.I0(r_SM_Main[2]), .I1(n46619), .I2(n46620), 
            .I3(r_SM_Main[1]), .O(n26084));
    defparam i41193_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i20070_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n25329));
    defparam i20070_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_81_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_13));   // verilog/uart_rx.v(97[17:39])
    defparam equal_81_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_83_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_14));   // verilog/uart_rx.v(97[17:39])
    defparam equal_83_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_877 (.I0(r_Bit_Index[0]), .I1(n16437), .I2(GND_net), 
            .I3(GND_net), .O(n16432));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_877.LUT_INIT = 16'hdddd;
    SB_LUT4 i41190_2_lut (.I0(r_SM_Main[2]), .I1(n49982), .I2(GND_net), 
            .I3(GND_net), .O(n26082));
    defparam i41190_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(n25923), .I1(\r_SM_Main_2__N_3032[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n49979));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'hcf70;
    SB_LUT4 i3_4_lut (.I0(n77), .I1(\r_Clock_Count[5] ), .I2(r_Clock_Count_c[6]), 
            .I3(n144), .O(n43440));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i141_4_lut (.I0(r_SM_Main[2]), .I1(n76), .I2(n43440), .I3(r_SM_Main[1]), 
            .O(n138));   // verilog/uart_rx.v(36[17:26])
    defparam i141_4_lut.LUT_INIT = 16'hafee;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n41870));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3032[2] ), .O(n16437));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\r_Clock_Count[1] ), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count_c[2]), .I3(r_Clock_Count_c[3]), .O(n77));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut (.I0(\r_Clock_Count[1] ), .I1(n81), .I2(r_Clock_Count_c[3]), 
            .I3(n119), .O(\r_SM_Main_2__N_3032[2] ));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff80;
    SB_LUT4 i2_3_lut_4_lut_adj_878 (.I0(r_Clock_Count_c[7]), .I1(r_Clock_Count_c[4]), 
            .I2(r_Clock_Count_c[6]), .I3(\r_Clock_Count[5] ), .O(n119));
    defparam i2_3_lut_4_lut_adj_878.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n2592, encoder1_position, GND_net, 
            n18615, clk32MHz, n18614, n18613, n18612, n18611, n18610, 
            n18609, n18608, n18607, n18606, n18605, n18604, n18603, 
            n18602, n18601, n18600, n18599, n18598, n18597, n18596, 
            n18595, n18594, n18532, data_o, n17970, count_enable, 
            PIN_18_c_1, n18618, reg_B, PIN_19_c_0, n17973, n43352) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2592;
    output [23:0]encoder1_position;
    input GND_net;
    input n18615;
    input clk32MHz;
    input n18614;
    input n18613;
    input n18612;
    input n18611;
    input n18610;
    input n18609;
    input n18608;
    input n18607;
    input n18606;
    input n18605;
    input n18604;
    input n18603;
    input n18602;
    input n18601;
    input n18600;
    input n18599;
    input n18598;
    input n18597;
    input n18596;
    input n18595;
    input n18594;
    input n18532;
    output [1:0]data_o;
    input n17970;
    output count_enable;
    input PIN_18_c_1;
    input n18618;
    output [1:0]reg_B;
    input PIN_19_c_0;
    input n17973;
    output n43352;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2583, n34809, n34810, n34808, n34807, n34806, n34805, 
        n34804, n34803, n34802, n34801, n34800, n34799, n34798, 
        count_direction, n34797, B_delayed, A_delayed, n34820, n34819, 
        n34818, n34817, n34816, n34815, n34814, n34813, n34812, 
        n34811;
    
    SB_LUT4 add_599_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2583), 
            .I3(n34809), .O(n2592[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_14 (.CI(n34809), .I0(encoder1_position[12]), .I1(n2583), 
            .CO(n34810));
    SB_LUT4 add_599_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2583), 
            .I3(n34808), .O(n2592[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_13 (.CI(n34808), .I0(encoder1_position[11]), .I1(n2583), 
            .CO(n34809));
    SB_LUT4 add_599_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2583), 
            .I3(n34807), .O(n2592[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_12 (.CI(n34807), .I0(encoder1_position[10]), .I1(n2583), 
            .CO(n34808));
    SB_LUT4 add_599_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2583), 
            .I3(n34806), .O(n2592[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_11 (.CI(n34806), .I0(encoder1_position[9]), .I1(n2583), 
            .CO(n34807));
    SB_LUT4 add_599_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2583), 
            .I3(n34805), .O(n2592[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_10 (.CI(n34805), .I0(encoder1_position[8]), .I1(n2583), 
            .CO(n34806));
    SB_LUT4 add_599_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2583), 
            .I3(n34804), .O(n2592[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_9 (.CI(n34804), .I0(encoder1_position[7]), .I1(n2583), 
            .CO(n34805));
    SB_LUT4 add_599_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2583), 
            .I3(n34803), .O(n2592[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_8 (.CI(n34803), .I0(encoder1_position[6]), .I1(n2583), 
            .CO(n34804));
    SB_LUT4 add_599_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2583), 
            .I3(n34802), .O(n2592[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_7 (.CI(n34802), .I0(encoder1_position[5]), .I1(n2583), 
            .CO(n34803));
    SB_LUT4 add_599_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2583), 
            .I3(n34801), .O(n2592[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_6 (.CI(n34801), .I0(encoder1_position[4]), .I1(n2583), 
            .CO(n34802));
    SB_LUT4 add_599_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2583), 
            .I3(n34800), .O(n2592[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_5 (.CI(n34800), .I0(encoder1_position[3]), .I1(n2583), 
            .CO(n34801));
    SB_LUT4 add_599_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2583), 
            .I3(n34799), .O(n2592[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_4 (.CI(n34799), .I0(encoder1_position[2]), .I1(n2583), 
            .CO(n34800));
    SB_LUT4 add_599_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2583), 
            .I3(n34798), .O(n2592[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_3 (.CI(n34798), .I0(encoder1_position[1]), .I1(n2583), 
            .CO(n34799));
    SB_LUT4 add_599_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n34797), .O(n2592[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_2 (.CI(n34797), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n34798));
    SB_CARRY add_599_1 (.CI(GND_net), .I0(n2583), .I1(n2583), .CO(n34797));
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18615));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18614));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18613));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18612));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18611));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18610));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18609));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18608));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18607));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18606));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18605));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18604));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18603));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n18602));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n18601));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n18600));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n18599));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n18598));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n18597));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n18596));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n18595));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n18594));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n18532));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_599_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2583), 
            .I3(n34820), .O(n2592[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_599_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2583), 
            .I3(n34819), .O(n2592[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17970));   // quad.v(35[10] 41[6])
    SB_CARRY add_599_24 (.CI(n34819), .I0(encoder1_position[22]), .I1(n2583), 
            .CO(n34820));
    SB_LUT4 add_599_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2583), 
            .I3(n34818), .O(n2592[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_23 (.CI(n34818), .I0(encoder1_position[21]), .I1(n2583), 
            .CO(n34819));
    SB_LUT4 add_599_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2583), 
            .I3(n34817), .O(n2592[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_22 (.CI(n34817), .I0(encoder1_position[20]), .I1(n2583), 
            .CO(n34818));
    SB_LUT4 add_599_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2583), 
            .I3(n34816), .O(n2592[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_21 (.CI(n34816), .I0(encoder1_position[19]), .I1(n2583), 
            .CO(n34817));
    SB_LUT4 add_599_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2583), 
            .I3(n34815), .O(n2592[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_20 (.CI(n34815), .I0(encoder1_position[18]), .I1(n2583), 
            .CO(n34816));
    SB_LUT4 add_599_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2583), 
            .I3(n34814), .O(n2592[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_19 (.CI(n34814), .I0(encoder1_position[17]), .I1(n2583), 
            .CO(n34815));
    SB_LUT4 add_599_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2583), 
            .I3(n34813), .O(n2592[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_18 (.CI(n34813), .I0(encoder1_position[16]), .I1(n2583), 
            .CO(n34814));
    SB_LUT4 add_599_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2583), 
            .I3(n34812), .O(n2592[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_17 (.CI(n34812), .I0(encoder1_position[15]), .I1(n2583), 
            .CO(n34813));
    SB_LUT4 add_599_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2583), 
            .I3(n34811), .O(n2592[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_16 (.CI(n34811), .I0(encoder1_position[14]), .I1(n2583), 
            .CO(n34812));
    SB_LUT4 add_599_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2583), 
            .I3(n34810), .O(n2592[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_599_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_599_15 (.CI(n34810), .I0(encoder1_position[13]), .I1(n2583), 
            .CO(n34811));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(data_o[0]), .I2(B_delayed), 
            .I3(A_delayed), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i915_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2583));   // quad.v(37[5] 40[8])
    defparam i915_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.PIN_18_c_1(PIN_18_c_1), .clk32MHz(clk32MHz), 
            .n18618(n18618), .data_o({data_o}), .reg_B({reg_B}), .PIN_19_c_0(PIN_19_c_0), 
            .n17973(n17973), .n43352(n43352), .GND_net(GND_net)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (PIN_18_c_1, clk32MHz, n18618, data_o, reg_B, 
            PIN_19_c_0, n17973, n43352, GND_net) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input PIN_18_c_1;
    input clk32MHz;
    input n18618;
    output [1:0]data_o;
    output [1:0]reg_B;
    input PIN_19_c_0;
    input n17973;
    output n43352;
    input GND_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3463, n2;
    
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_18_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18618));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1194__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_19_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1194__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1194__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17973));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n43352));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i28903_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i28903_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i28896_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i28896_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n43352), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3463));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i28894_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i28894_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, deadband, \Kp[4] , \PID_CONTROLLER.err[21] , 
            \pwm_23__N_3310[10] , \pwm_23__N_3310[6] , \pwm_23__N_3310[4] , 
            PWMLimit, \PID_CONTROLLER.result[19] , n18644, pwm, clk32MHz, 
            n18643, n18642, n18641, n18639, n18637, n18636, n18635, 
            n18633, n18632, \PID_CONTROLLER.err[23] , n18630, n18629, 
            n18628, n18626, n18624, n18623, n18622, \PID_CONTROLLER.result[17] , 
            \Kp[5] , n18574, \Kp[6] , \Kp[7] , n21, n9, \PID_CONTROLLER.err[31] , 
            n27, n13, \Kp[1] , \PID_CONTROLLER.err[22] , \Kp[0] , 
            n18495, \PID_CONTROLLER.err_prev[31] , n18494, \PID_CONTROLLER.err_prev[23] , 
            n18493, \PID_CONTROLLER.err_prev[22] , n18492, \PID_CONTROLLER.err_prev[21] , 
            n18491, \PID_CONTROLLER.err_prev[20] , n18490, \PID_CONTROLLER.err_prev[19] , 
            n18489, \PID_CONTROLLER.err_prev[18] , n18488, \PID_CONTROLLER.err_prev[17] , 
            n18487, \PID_CONTROLLER.err_prev[16] , n18486, \PID_CONTROLLER.err_prev[15] , 
            n18485, \PID_CONTROLLER.err_prev[14] , n18484, \PID_CONTROLLER.err_prev[13] , 
            n18483, \PID_CONTROLLER.err_prev[12] , n18482, \PID_CONTROLLER.err_prev[11] , 
            n18481, \PID_CONTROLLER.err_prev[10] , n18480, \PID_CONTROLLER.err_prev[9] , 
            n18479, \PID_CONTROLLER.err_prev[8] , n18478, \PID_CONTROLLER.err_prev[7] , 
            n18477, \PID_CONTROLLER.err_prev[6] , n18476, \PID_CONTROLLER.err_prev[5] , 
            n18475, \PID_CONTROLLER.err_prev[4] , n18474, \PID_CONTROLLER.err_prev[3] , 
            n18473, \PID_CONTROLLER.err_prev[2] , n18472, \PID_CONTROLLER.err_prev[1] , 
            \Kp[2] , \Kp[3] , \PID_CONTROLLER.result[10] , \PID_CONTROLLER.result[13] , 
            n387, n21_adj_1, \Kd[1] , n9_adj_2, \Kd[0] , \Kd[2] , 
            \Ki[0] , n27_adj_3, n13_adj_4, \Kd[3] , \Ki[1] , n35, 
            \Kd[4] , n39, \Kd[5] , \Ki[2] , \PID_CONTROLLER.err[0] , 
            PIN_7_c_1, PIN_6_c_0, n22, \Kd[6] , \Ki[3] , \Kd[7] , 
            VCC_net, n853, GATES_5__N_3405, n44276, n855, n856, 
            \Ki[4] , n857, pwm_23__N_3307, n859, n860, n861, n862, 
            n863, n864, n865, n866, n867, n868, n869, n870, 
            n871, n872, n873, n874, n875, n46548, \Ki[5] , n448, 
            n449, n450, n451, n453, n455, n456, \PID_CONTROLLER.err[1] , 
            \PID_CONTROLLER.err[2] , \Ki[6] , n457, \PID_CONTROLLER.err[9] , 
            \Ki[7] , n459, n460, n462, n463, n464, \PID_CONTROLLER.err[5] , 
            \PID_CONTROLLER.result[6] , n466, \PID_CONTROLLER.result[4] , 
            n468, n469, n470, n471, n27_adj_5, n13_adj_6, n414, 
            n403, n35_adj_7, n9_adj_8, n21_adj_9, n410, n416, n401, 
            pwm_count, n407, n39_adj_10, \PID_CONTROLLER.err[6] , \PID_CONTROLLER.err[7] , 
            \PID_CONTROLLER.err[3] , \PID_CONTROLLER.err[8] , \PID_CONTROLLER.err[4] , 
            hall1, hall2, \GATES_5__N_3398[5] , hall3, n48474, \PID_CONTROLLER.err_prev[0] , 
            n25, n30, n26, PIN_8_c_2, PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, 
            \PID_CONTROLLER.err[10] , \PID_CONTROLLER.err[11] , \PID_CONTROLLER.err[12] , 
            \PID_CONTROLLER.err[13] , \PID_CONTROLLER.err[14] , \PID_CONTROLLER.err[15] , 
            \PID_CONTROLLER.err[16] , \PID_CONTROLLER.err[17] , \PID_CONTROLLER.err[18] , 
            \PID_CONTROLLER.err[19] , \PID_CONTROLLER.err[20] , \motor_state[23] , 
            \motor_state[22] , \motor_state[21] , \motor_state[20] , \motor_state[19] , 
            \motor_state[18] , \motor_state[17] , \motor_state[16] , \motor_state[15] , 
            \motor_state[14] , \motor_state[13] , \motor_state[12] , \motor_state[11] , 
            \motor_state[10] , \motor_state[9] , \motor_state[8] , \motor_state[7] , 
            \motor_state[6] , \motor_state[5] , \motor_state[4] , \motor_state[3] , 
            \motor_state[2] , \motor_state[1] , \motor_state[0] , n17967, 
            n43362, n13_adj_11, n9_adj_12, IntegralLimit, setpoint, 
            n16, n5, n29) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input [23:0]deadband;
    input \Kp[4] ;
    output \PID_CONTROLLER.err[21] ;
    output \pwm_23__N_3310[10] ;
    output \pwm_23__N_3310[6] ;
    output \pwm_23__N_3310[4] ;
    input [23:0]PWMLimit;
    output \PID_CONTROLLER.result[19] ;
    input n18644;
    output [23:0]pwm;
    input clk32MHz;
    input n18643;
    input n18642;
    input n18641;
    input n18639;
    input n18637;
    input n18636;
    input n18635;
    input n18633;
    input n18632;
    output \PID_CONTROLLER.err[23] ;
    input n18630;
    input n18629;
    input n18628;
    input n18626;
    input n18624;
    input n18623;
    input n18622;
    output \PID_CONTROLLER.result[17] ;
    input \Kp[5] ;
    input n18574;
    input \Kp[6] ;
    input \Kp[7] ;
    input n21;
    input n9;
    output \PID_CONTROLLER.err[31] ;
    input n27;
    input n13;
    input \Kp[1] ;
    output \PID_CONTROLLER.err[22] ;
    input \Kp[0] ;
    input n18495;
    output \PID_CONTROLLER.err_prev[31] ;
    input n18494;
    output \PID_CONTROLLER.err_prev[23] ;
    input n18493;
    output \PID_CONTROLLER.err_prev[22] ;
    input n18492;
    output \PID_CONTROLLER.err_prev[21] ;
    input n18491;
    output \PID_CONTROLLER.err_prev[20] ;
    input n18490;
    output \PID_CONTROLLER.err_prev[19] ;
    input n18489;
    output \PID_CONTROLLER.err_prev[18] ;
    input n18488;
    output \PID_CONTROLLER.err_prev[17] ;
    input n18487;
    output \PID_CONTROLLER.err_prev[16] ;
    input n18486;
    output \PID_CONTROLLER.err_prev[15] ;
    input n18485;
    output \PID_CONTROLLER.err_prev[14] ;
    input n18484;
    output \PID_CONTROLLER.err_prev[13] ;
    input n18483;
    output \PID_CONTROLLER.err_prev[12] ;
    input n18482;
    output \PID_CONTROLLER.err_prev[11] ;
    input n18481;
    output \PID_CONTROLLER.err_prev[10] ;
    input n18480;
    output \PID_CONTROLLER.err_prev[9] ;
    input n18479;
    output \PID_CONTROLLER.err_prev[8] ;
    input n18478;
    output \PID_CONTROLLER.err_prev[7] ;
    input n18477;
    output \PID_CONTROLLER.err_prev[6] ;
    input n18476;
    output \PID_CONTROLLER.err_prev[5] ;
    input n18475;
    output \PID_CONTROLLER.err_prev[4] ;
    input n18474;
    output \PID_CONTROLLER.err_prev[3] ;
    input n18473;
    output \PID_CONTROLLER.err_prev[2] ;
    input n18472;
    output \PID_CONTROLLER.err_prev[1] ;
    input \Kp[2] ;
    input \Kp[3] ;
    output \PID_CONTROLLER.result[10] ;
    output \PID_CONTROLLER.result[13] ;
    output n387;
    input n21_adj_1;
    input \Kd[1] ;
    input n9_adj_2;
    input \Kd[0] ;
    input \Kd[2] ;
    input \Ki[0] ;
    input n27_adj_3;
    input n13_adj_4;
    input \Kd[3] ;
    input \Ki[1] ;
    input n35;
    input \Kd[4] ;
    input n39;
    input \Kd[5] ;
    input \Ki[2] ;
    output \PID_CONTROLLER.err[0] ;
    output PIN_7_c_1;
    output PIN_6_c_0;
    input n22;
    input \Kd[6] ;
    input \Ki[3] ;
    input \Kd[7] ;
    input VCC_net;
    output n853;
    input GATES_5__N_3405;
    output n44276;
    output n855;
    output n856;
    input \Ki[4] ;
    output n857;
    output pwm_23__N_3307;
    output n859;
    output n860;
    output n861;
    output n862;
    output n863;
    output n864;
    output n865;
    output n866;
    output n867;
    output n868;
    output n869;
    output n870;
    output n871;
    output n872;
    output n873;
    output n874;
    output n875;
    output n46548;
    input \Ki[5] ;
    output n448;
    output n449;
    output n450;
    output n451;
    output n453;
    output n455;
    output n456;
    output \PID_CONTROLLER.err[1] ;
    output \PID_CONTROLLER.err[2] ;
    input \Ki[6] ;
    output n457;
    output \PID_CONTROLLER.err[9] ;
    input \Ki[7] ;
    output n459;
    output n460;
    output n462;
    output n463;
    output n464;
    output \PID_CONTROLLER.err[5] ;
    output \PID_CONTROLLER.result[6] ;
    output n466;
    output \PID_CONTROLLER.result[4] ;
    output n468;
    output n469;
    output n470;
    output n471;
    input n27_adj_5;
    input n13_adj_6;
    output n414;
    output n403;
    input n35_adj_7;
    input n9_adj_8;
    input n21_adj_9;
    output n410;
    output n416;
    output n401;
    output [8:0]pwm_count;
    output n407;
    input n39_adj_10;
    output \PID_CONTROLLER.err[6] ;
    output \PID_CONTROLLER.err[7] ;
    output \PID_CONTROLLER.err[3] ;
    output \PID_CONTROLLER.err[8] ;
    output \PID_CONTROLLER.err[4] ;
    input hall1;
    input hall2;
    output \GATES_5__N_3398[5] ;
    input hall3;
    input n48474;
    output \PID_CONTROLLER.err_prev[0] ;
    input n25;
    input n30;
    input n26;
    output PIN_8_c_2;
    output PIN_9_c_3;
    output PIN_10_c_4;
    output PIN_11_c_5;
    output \PID_CONTROLLER.err[10] ;
    output \PID_CONTROLLER.err[11] ;
    output \PID_CONTROLLER.err[12] ;
    output \PID_CONTROLLER.err[13] ;
    output \PID_CONTROLLER.err[14] ;
    output \PID_CONTROLLER.err[15] ;
    output \PID_CONTROLLER.err[16] ;
    output \PID_CONTROLLER.err[17] ;
    output \PID_CONTROLLER.err[18] ;
    output \PID_CONTROLLER.err[19] ;
    output \PID_CONTROLLER.err[20] ;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \motor_state[0] ;
    input n17967;
    output n43362;
    input n13_adj_11;
    input n9_adj_12;
    input [23:0]IntegralLimit;
    input [23:0]setpoint;
    input n16;
    input n5;
    output n29;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [28:0]n8741;
    wire [27:0]n8772;
    
    wire n36264, n47706, n8, n15, n47961, n48467, n35889;
    wire [20:0]n8469;
    
    wire n35890;
    wire [21:0]n8445;
    
    wire n35888, n36265, n35887, n35886;
    wire [22:0]n1801;
    wire [22:0]n1802;
    
    wire n36856, n36736;
    wire [22:0]n1797;
    
    wire n36737, n36544;
    wire [14:0]n9084;
    
    wire n36545;
    wire [31:0]pwm_23__N_3310;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    
    wire n18, n36263, n35885;
    wire [31:0]n57;
    
    wire n34665;
    wire [33:0]n282;
    
    wire n36735;
    wire [15:0]n9066;
    
    wire n725, n36543, n35884, n41, n36262, n707, n35883, n34666, 
        n36261, n628, n36542, n610, n35882, n513, n35881, n34664, 
        n416_c, n35880, n36260, n319, n35879, n222, n35878, n36259, 
        n32, n125, n531, n36541, n36857, n36734;
    wire [20:0]n9225;
    wire [19:0]n9555;
    
    wire n36943;
    wire [22:0]n8420;
    
    wire n35877, n36258, n36855, n35876, n37, n35875, n434, n36540, 
        n36733, n686, n36257, n512, n36732, n35874, n36944, n36942, 
        n337, n36539, n36854, n439, n36731, n35873, n36941, n589_adj_3465, 
        n36256, n35872, n240, n36538, n29_c, n35871, n36853, n31, 
        n50, n143, n7, n492, n36255, n35870, n35869, n366, n36730, 
        n36852;
    wire [16:0]n9047;
    
    wire n36537, n36536, n293, n36729, n395, n36254, n36535, n35868, 
        n298, n36253, n35867, n35866, n35865, n201, n36252, n35864, 
        n220, n36728, n36534, n11, n104, n35863;
    wire [0:0]n6817;
    wire [29:0]n8709;
    
    wire n36251;
    wire [31:0]n58;
    
    wire n35862;
    wire [55:0]n191;
    
    wire n36250, n704, n35861, n607, n35860, n36940, n510, n35859, 
        n36249, n36533, n413, n35858, n36851, n147, n36727, n36532, 
        n316, n35857, n36248, n33, n219_adj_3466, n35856, n11_adj_3467, 
        n36939, n29_adj_3468, n122, n36247;
    wire [23:0]n8394;
    
    wire n35855, n36850, n35854, n36531, n35853, n36246, n35852, 
        n35851, n36245, n35850, n5_c, n74, n35849, n36530, n36244, 
        n35848, n35847, n36243;
    wire [13:0]n9722;
    wire [12:0]n9738;
    
    wire n36726, n36529, n35846, n36242, n35845, n36725, n35844, 
        n36241, n35843, n36528, n35842, n36240, n35841, n35840, 
        n36239, n35839, n722, n36527, n701, n35838, n36238, n604, 
        n35837, n36849, n36724, n507, n35836, n36237, n410_c, 
        n35835, n625, n36526, n313_adj_3473, n35834, n36236, n216, 
        n35833, n26_c, n119, n36235;
    wire [24:0]n8367;
    
    wire n35832, n528, n36525, n35831, n36234, n35830, n545, n36938, 
        n36723, n35829, n36233, n35828, n431, n36524, n35827, 
        n36232, n35826, n35825, n36231, n35824, n34663, n334, 
        n36523, n35823, n36230, n35822, n36848, n36722, n35821, 
        n36229, n35820, n34662, n237_adj_3476, n36522, n35819, n36228, 
        n35818, n35817, n680, n36227, n35816, n34661, n47, n140, 
        n452, n35815, n583, n36226, n698, n35814, n36721, n601_adj_3478, 
        n35813, n486, n36225, n504, n35812, n34660;
    wire [17:0]n9027;
    
    wire n36521, n15_adj_3479, n407_c, n35811, n389, n36224, n310_adj_3480, 
        n35810, n34659, n36520, n213, n35809, n292, n36223, n23, 
        n116, n34658;
    wire [25:0]n8339;
    
    wire n35808, n195, n36222, n35807, n34657, n527, n36847, n36720, 
        n36519, n35806, n5_adj_3483, n98, n35805, n34656, n35804;
    wire [18:0]n9591;
    
    wire n36221, n35803, n34655, n36518, n36220, n35802, n34654, 
        n35801, n36219, n35800, n34653, n472, n36937, n36719, 
        n36517, n36218, n35799, n35798, n36217, n35797, n35796, 
        n36516, n36216, n35795, n45, n35794, n36215, n35793, n35792, 
        n34652, n454, n36846, n36718, n36515, n36214, n35791, 
        n35790, n17_adj_3486, n36213, n19_adj_3487, n43, n41_adj_3488, 
        n39_c, n36514, n695, n35789, n45_adj_3489, n43_adj_3490, 
        n37_adj_3491, n23_adj_3492, n25_adj_3493, n18640, n18638, 
        n18634;
    wire [31:0]n60;
    
    wire n18631, n18627, n18625, n29_adj_3494;
    wire [31:0]n61;
    
    wire n31_adj_3496, n35_c, n33_adj_3497, n549, n646, n36513, 
        n598, n35788, n36212, n501, n35787, n17_adj_3498, n19_adj_3499, 
        n11_adj_3500, n15_adj_3502, n743, n47150, n47144, n164, 
        n71, n404, n35786, n36211, n307_adj_3507, n35785, n36210, 
        n34651, n399, n36717, n12, n30_adj_3508, n261, n358, n47161, 
        n47934, n47930, n48795, n455_adj_3509, n48283, n48914, n210, 
        n35784, n6, n48419, n36209, n552, n48420, n16_adj_3510, 
        n24_adj_3511, n47123, n8_adj_3512, n47121, n48470, n47714, 
        n4, n649, n48417, n48418, n746, n47140, n10_adj_3514, 
        n47138, n48853, n47716, n49010, n49011, n48968, n47125, 
        n48734, n47722, n167, n48899, n264, n48, n43052, n43059, 
        n56, n361, n23_adj_3515, n25_adj_3516, n43083, n43089, n47999, 
        n47971, n458_adj_3519, n20_adj_3520, n113, n125_adj_3521, 
        n47272, n47250, n32_adj_3523, n48313, n555, n652, n48801, 
        n47973, n326, n36716, n47209, n47953, n50655, n222_adj_3526, 
        n28_adj_3527, n47215, n47957, n50650, n47955, n36512;
    wire [9:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(33[22:30])
    
    wire n72, n50612, n47207, n50624, n48297, n50616, n48797, 
        n749, n47266, n319_adj_3530, n145, n12_adj_3531, n30_adj_3533, 
        n98_adj_3534, n48011, n48329, n48327, n47268, n416_adj_3536, 
        n48600, n48994, n47983, n48596, n48918, n49036, n36511, 
        n6_adj_3538, n48427, n47965, n54, n47233, n50608, n18_adj_3539, 
        n48465, n47704, n16_adj_3540, n24_adj_3541, n8_adj_3542, n47248, 
        n48849, n48850, n48592, n48893, n47702, n26_adj_3543, n47205, 
        n719, n36510, n36208;
    wire [26:0]n8310;
    
    wire n35783, n35782, n36207, n513_adj_3544, n35781, n34650, 
        n381, n36845, n24_adj_3547, n35780, n35779, n36206, n35778, 
        n622, n36509, n35777, n36205, n35776, n35775, n253, n36204, 
        n35774, n218_adj_3548;
    wire [31:0]\PID_CONTROLLER.result_31__N_3353 ;
    
    wire n36715, n525, n36508, n35773, n180_adj_3549, n36203, n752, 
        n34, n35772, n48851;
    wire [24:0]\PID_CONTROLLER.err_31__N_3175 ;
    
    wire n171, n35771;
    wire [5:0]GATES_5__N_3138;
    
    wire n428, n36507, n35_adj_3550, n107, n35770, n35769, n48852, 
        n101, n48711, n35768, n36714;
    wire [17:0]n9624;
    
    wire n36202, n36201, n35767, n8_adj_3551, n48421, n48422, n331, 
        n36506, n36200, n35766, n35765, n36936, n308_adj_3555, n36844, 
        n36199, n35764, n692, n35763, n234_adj_3556, n36505, n36198, 
        n595, n35762, n498, n35761, n610_adj_3557, n36197, n47940, 
        n401_c, n35760, n30_adj_3558, n198, n304, n35759, n44, 
        n137, n36196, n207, n35758, n43813, n47712, n47943, n17_adj_3559, 
        n110, n48301;
    wire [27:0]n8280;
    
    wire n35757, n47710, n48469, n36195, n4_adj_3560, n34649, n48437;
    wire [18:0]n9006;
    
    wire n36504, n36194, n48438, n35756, n35755, n36503, n36193, 
        n35754, n35753, n291;
    wire [11:0]n9753;
    
    wire n36713, n36192, n35752, n35751, n47262, n36502, n36191, 
        n35750, n707_adj_3562, n35749, n10_adj_3563, n47260, n48847, 
        n36935, n295, n235_adj_3565, n36843, n36712, n36190, n35748, 
        n35747, n36501, n36189, n35746, n35745, n36188, n35744, 
        n35743, n36500, n36187, n35742, n35741, n36711, n36186, 
        n35740, n35739, n36499, n36185, n35738, n35737, n689, 
        n35736, n592, n35735, n36498;
    wire [16:0]n9654;
    
    wire n36184, n36183, n495, n35734, n47692, n398, n35733, n162, 
        n36842, n36710, n301, n35732, n392, n36182, n204, n35731, 
        n36497, n36181, n14, n107_adj_3567, n46520, n25957, n36934, 
        n36709, n36496;
    wire [28:0]n8249;
    
    wire n35730, n36180, n34765, n35729, n36179;
    wire [23:0]n63;
    
    wire n34764;
    wire [23:0]n852;
    
    wire n49008, n49009, n489, n34763, n35728, n48972, n49072, 
        n36933, n34762, n36708, n35727, n48895, n36495, n36178, 
        n20_adj_3571, n89, n47698, pwm_23__N_3309, n36177, n35726, 
        n48897, n364, n36494, n36707, n36493, n35725, n34761, 
        n716, n36492, n35724, n36176, n35723, n34760, n36706, 
        n619, n36491, n36175, n35722, n34759, n36174, n34758, 
        n36173;
    wire [22:0]n1800;
    
    wire n36840, n522, n36490, n35721, n35720, n35719, n36172, 
        n35718, n34757, n1699, n34756, n36171, n425, n36489, n35717, 
        n35716, n34755, n36705, n36170, n35715, n328, n36488, 
        n35714, n34754, n36704, n36169, n36168, n231_adj_3581, n36487, 
        n35713, n35712, n36703, n35711;
    wire [15:0]n9681;
    
    wire n36167, n35710, n34753, n35709, n41_adj_3583, n134, n686_adj_3584, 
        n35708;
    wire [19:0]n8984;
    
    wire n36486, n36166, n589_adj_3585, n35707, n36485, n34752, 
        n36165, n492_adj_3587, n35706, n36839, n395_adj_3588, n35705, 
        n36164, n36702, n298_adj_3589, n35704, n36163, n36838, n34751, 
        n36837, n201_adj_3591, n35703, n36484, n11_adj_3592, n104_adj_3593, 
        n36162;
    wire [22:0]n1804;
    wire [21:0]n9201;
    
    wire n36932, n36931;
    wire [0:0]n6807;
    wire [29:0]n8217;
    
    wire n35702, n34750, n36836;
    wire [55:0]n64;
    
    wire n35701, n34749;
    wire [10:0]n9767;
    
    wire n36701, n36483, n36161, n36700, n36835, n35700, n34748, 
        n36834, n36699, n36482, n36930, n36160, n36833, n36698, 
        n35699, n36929, n36697, n35698, n36159, n34747, n36928, 
        n36481, n36832, n36158, n36696, n34746, n35697, n36831, 
        n36695, n36157, n35696, n35695, n36927, n36830, n35694, 
        n36694, n36926, n36829, n36480, n36925, n36693, n36156, 
        n36828, n36692, n36479, n35693, n34745, n36155, n36478, 
        n36691, n36154, n35692, n35691, n36477, n36153, n35690, 
        n36152, n36827, n36476, n34744, n35689, n34743, n35688, 
        n36475, n35687, n36924, n36474;
    wire [14:0]n9705;
    
    wire n36151;
    wire [9:0]n9780;
    
    wire n36690, n35686, n36150, n36826, n713, n36473, n25958, 
        n36923, n36149, n36689, n616, n36472, n586, n176, n36688, 
        n36825, n683, n36922, n244_adj_3607, n36148, n35685, n519, 
        n36471, n524, n36824, n36687, n422, n36470, n35684, n36147, 
        n437, n35683, n467, n36686, n564, n6_adj_3612;
    wire [3:0]n9612;
    wire [4:0]n9577;
    
    wire n325, n36469, n35682, n36921, n36920, n228_adj_3613, n36468, 
        n36146, n451_c, n36823, n49785, n34742, n34741, n35681, 
        n36145, n38, n131_adj_3617, n35680, n36685, n36144;
    wire [20:0]n8961;
    
    wire n36467, n36143, n36142, n378, n36822, n36466, n35679, 
        n36141, n36465, n680_adj_3618, n35678, n36684, n36464, n36140, 
        n583_adj_3620, n35677, n36139, n486_adj_3621, n35676, n273, 
        n36683, n36463, n389_adj_3622, n35675, n36138, n80, n34740, 
        n292_adj_3624, n35674, n36137, n36462, n36136, n195_adj_3625, 
        n35673, n36135, n36919, n305, n36821, n36682, n34739, 
        n36461, n23926, n34738, n36460, n36681, n36134, n5_adj_3630, 
        n98_adj_3631, n36918, n36459;
    wire [5:0]n9547;
    
    wire n44039, n658, n35672;
    wire [4:0]n9584;
    
    wire n561, n35671, n370_adj_3633, n232_adj_3635, n36820, n36458, 
        n34094, n34487, n34737, n36133, n159, n36819;
    wire [8:0]n9792;
    
    wire n36680, n36679, n36457, n36132, n23686, n34736, n36456, 
        n36131, n36130;
    wire [3:0]n9618;
    
    wire n470_c, n35670, n373, n35669, n36455, n36129, n36678, 
        n276, n35668, n34735, n36128, n36454, n36677, n83, n179, 
        n36127, n35667, n655, n35666, n710, n36453, n35665, n8_adj_3640, 
        n36917, n17_adj_3642, n86, n36676, n36126, n34734, n613, 
        n36452, n35664, n36125, n36124;
    wire [22:0]n1799;
    
    wire n36817, n35663, n4_adj_3644, n6_adj_3645, n35662, n1695, 
        n36675, n44310, n36123, n4_adj_3646, n14_adj_3647, n516_adj_3648, 
        n36451, n43598, n419, n36450, n36122, n36121, n35661, 
        n36120, n35660, n35659, n35658, n322, n36449, n36119, 
        n35657, n536, n36916, n36816, n101_adj_3650;
    wire [31:0]n66;
    
    wire n34898, n35656, n8_adj_3651, n198_adj_3652, n463_c, n36915, 
        n36674, n295_adj_3653, n225_adj_3654, n36448, n36118, n35_adj_3655, 
        n128_adj_3656, n35655, n36117, n392_adj_3657, n510_adj_3658, 
        n36815, n34733, n35654;
    wire [21:0]n8937;
    
    wire n36447, n36673, n35653, n36446, n489_adj_3660, n35652, 
        n317, n586_adj_3661, n34897, n583_adj_3662, n683_adj_3663, 
        n36445, n390, n36914, n36116, n36814, n23155, n34732, 
        n35651, n36444, n35650, n36115, n36114, n36672, n36113, 
        n35649, n35648, n36443, n36112, n35647, n36111, n35646, 
        n35645, n36110, n34731, n35644, n36671, n36442, n36109, 
        n36441, n36670, n35643, n36108, n36913, n36440, n36107, 
        n35642, n36669, n36106, n36105, n36439, n35641, n36104, 
        n35640, n35639, n36438, n34896, n34730;
    wire [5:0]n9539;
    
    wire n35638, n36437, n36103, n36436, n35637, n36813, n36102, 
        n36101, n36668, n35636, n1, n34729, n35635, n34895, n36435, 
        n35634, n36100, n36912, n36812, n36099, n36098, n34728, 
        n36667, n4_adj_3668, n36097, n34377, n34352, n36434, n36433, 
        n36096, n36811, n34894, n34727, n36095, n7_adj_3670, n8_adj_3671, 
        n8_adj_3672, n36432, n36666, n36094, n36431, n36911;
    wire [6:0]n8700;
    
    wire n36093, n36092, n36665, n36091, n36430, n36810, n36090, 
        n36089, n36429, n34893, n34726, n36088, n36809, n36664, 
        n36428;
    wire [7:0]n8690;
    
    wire n36087, n36086, n36427, n1_adj_3674, n34725, n34892, n34724, 
        n36085, n36663, n36084;
    wire [22:0]n1803;
    
    wire n36909, n36808, n36083, n36662, n1_adj_3675, n34723;
    wire [22:0]n8912;
    
    wire n36426, n36082, n36425, n36081, n36424;
    wire [31:0]n67;
    
    wire n41_adj_3676;
    wire [8:0]n8679;
    
    wire n36080, n34891, n45_adj_3678, n43_adj_3680, n36079, n36661, 
        n36423, n36078, n36077, n34722;
    wire [8:0]n6821;
    
    wire n36991, n36807, n37_adj_3681, n1711, n36660, n36659, n36422, 
        n36421, n36076, n36075, n29_adj_3682, n31_adj_3683, n36990, 
        n36074, n36073, n23_adj_3684, n34890, n36658, n36420, n34721, 
        n34889, n34624, n34623, n36806, n36657, n36419;
    wire [9:0]n8667;
    
    wire n36072, n36071, n36070, n36418, n36069, n25_adj_3686, n34720, 
        n36417, n36989, n36908, n36068, n34888, n36656, n36067, 
        n17_adj_3688, n34622, n36416, n36805, n19_adj_3690, n34887, 
        n36066, n36415, n36988, n355, n36065, n36414, n258, n36064, 
        n36655, n36413, n33_adj_3692, n11_adj_3693, n34886, n36987, 
        n36907, n36654, n15_adj_3695, n36804, n36412, n34719, n68, 
        n161, n34885, n36986, n47101, n36411;
    wire [10:0]n8654;
    
    wire n36063, n36906, n36062, n12_adj_3698, n34621, n34718, n34884, 
        n34620, n34717, n10_adj_3701, n30_adj_3703, n36905, n704_adj_3704, 
        n36410;
    wire [6:0]n69;
    wire [6:0]Kd_delay_counter;   // verilog/motorControl.v(27[13:29])
    
    wire n36803, n36061, n36985, n36060, n36653, n36904, n34883, 
        n36802, n740, n36059, n36652, n47118, n47902, n47898, 
        n643, n36058, n34716, n48789, n607_adj_3708, n36409, n34619, 
        n546, n36057, n48267, n36651, n34882, n36650, n510_adj_3710, 
        n36408, n36984, n521, n36801, n48912, n413_adj_3712, n36407, 
        n34715, n449_adj_3713, n36056, n36649, n352, n36055, n316_adj_3714, 
        n36406, n6_adj_3715, n48411, n48412, n255, n36054, n16_adj_3717, 
        n65, n158, n219_adj_3718, n36405;
    wire [11:0]n8640;
    
    wire n36053, n36052, n8_adj_3720, n36051, n34881, n24_adj_3721, 
        n47107, n47087, n47085, n48928, n36983, n34714, n47728, 
        n10_adj_3723, n36050, n29_adj_3724, n122_adj_3725, n36648, 
        n34618, n8_adj_3728;
    wire [23:0]n8886;
    
    wire n36404, n36049, n737, n36048, n34880, n36403;
    wire [8:0]n70;
    
    wire n12_adj_3730, n46522, n4_adj_3732, n48409, n640, n36047, 
        n34713, n36402, n448_adj_3735, n36800, n48410, n36647, n36982, 
        n47097, n543, n36046, n47095, n48855;
    wire [9:0]n73;
    
    wire n55_adj_3736, n47730, n34879, n49012, n49013, n375, n36799, 
        n36981, n36903, n446, n36045, n34617, n48966, n302, n36798, 
        n34712, n36401, n349, n36044, n47089, n34878, n49050, 
        n47736, n49068, n36400, n36646, n43824, n49069, n252, 
        n36043, n36645, n62, n155_adj_3741, n36399, n36398, n36902, 
        n229_adj_3743, n36797, n34877, n36397, n34616, n34876, n34711;
    wire [12:0]n8625;
    
    wire n36042, n34875, n34710, n36644, n36396, n36041, n34874, 
        n34709, n36040, n34873, n34872, n34615, n34708, n34871, 
        n36643, n36395, n156_adj_3746, n36796, n36394, n34870, n36393, 
        n36980, n36039, n14_adj_3747, n83_adj_3748, n36038, n36901, 
        n34707, n34706, n34869, n36037, n36979, n34868, n734, 
        n36036, n36392, n36978, n36900, n637, n36035;
    wire [6:0]n9192;
    
    wire n752_adj_3752, n36642, n36391, n540, n36034, n34705, n34614;
    wire [22:0]n1798;
    
    wire n36794, n655_adj_3754, n36641, n34704, n443_adj_3755, n36033, 
        n34703, n35519, n35518, n36390, n36977, n346, n36032, 
        n35517, n35516, n36976, n36899, n249, n36031, n35515, 
        n35514, n36898, n1691, n36793, n35513, n558, n36640, n36389, 
        n59, n152_adj_3759, n36975, n34613, n35512, n36388, n36792;
    wire [13:0]n8609;
    
    wire n36030, n461, n36639, n36897, n364_adj_3762, n36638, n34612, 
        n36791, n267, n36637, n36029, n701_adj_3764, n36387, n35511, 
        n604_adj_3766, n36386, n36790, n36028, n170_adj_3767, n36896, 
        n34611, n507_adj_3769, n36385, n36027;
    wire [7:0]n9182;
    
    wire n36636, n749_adj_3770, n36635, n410_adj_3771, n36384, n36026, 
        n36789, n36025, n34610, n36024, n313_adj_3773, n36383, n731, 
        n36023, n36974, n36895, n652_adj_3776, n36634, n634, n36022, 
        n34702, n216_adj_3777, n36382, n34609, n537_adj_3779, n36021, 
        n34608, n26_adj_3781, n119_adj_3782, n36973, n36894, n440, 
        n36020;
    wire [24:0]n8859;
    
    wire n36381, n343, n36019, n555_adj_3785, n36633, n36380, n246_adj_3786, 
        n36018, n56_adj_3787, n149_adj_3788, n36788, n36379;
    wire [14:0]n8592;
    
    wire n36017, n36016, n35497, n35496, n35495, n36015, n35494, 
        n458_adj_3792, n36632, n36378, n35493, n36014, n35492, n35491, 
        n36013, n35490, n36377, n36012, n35489, n35488, n36011, 
        n35487, n361_adj_3799, n36631, n36376, n35486, n36010, n35485, 
        n35484, n728, n36009, n36787, n36375, n631, n36008, n534, 
        n36007, n264_adj_3803, n36630, n36374, n437_adj_3804, n36006, 
        n340, n36005, n533, n36893, n36373, n243_adj_3806, n36004, 
        n53_adj_3807, n146_adj_3808, n74_adj_3809, n167_adj_3810, n36372;
    wire [15:0]n8574;
    
    wire n36003, n36002, n36786, n36371, n36001, n36000;
    wire [8:0]n9171;
    
    wire n36629, n36370, n35999, n35998, n36628, n36369, n35997, 
        n35996, n36368, n35995, n725_adj_3811, n35994, n36785, n746_adj_3812, 
        n36627, n36367, n628_adj_3813, n35993, n531_adj_3814, n35992, 
        n36366, n434_adj_3815, n35991, n337_adj_3816, n35990, n36972, 
        n460_adj_3819, n36892, n649_adj_3820, n36626, n36365, n240_adj_3821, 
        n35989, n50_adj_3822, n143_adj_3823, n36364;
    wire [16:0]n8555;
    
    wire n35988, n35987, n35986, n36784, n552_adj_3824, n36625, 
        n698_adj_3825, n36363, n35985, n34607, n455_adj_3827, n36624, 
        n35984, n34606, n36783, n34605, n34701, n358_adj_3830, n36623, 
        n601_adj_3831, n36362, n36782, n35983, n34700, n36971, n387_adj_3833, 
        n36891, n34604, n261_adj_3835, n36622, n35982, n504_adj_3836, 
        n36361, n34699, n407_adj_3837, n36360, n35981, n35980, n71_adj_3838, 
        n164_adj_3839, n310_adj_3840, n36359, n35979, n34603, n34698;
    wire [9:0]n9159;
    
    wire n36621, n41825, n722_adj_3842, n35978, n34602, n36970, 
        n314_adj_3845, n36890, n36781, n36620, n36780, n213_adj_3846, 
        n36358, n625_adj_3847, n35977, n34697, n36969, n34601, n528_adj_3849, 
        n35976, n241_adj_3851, n36889, n34600, n36968, n20_adj_3853, 
        n26_adj_3854, n24_adj_3855, n28_adj_3856, n23_adj_3857, n168_adj_3859, 
        n36888, n17_adj_3860, n34696, n23_adj_3861, n116_adj_3862, 
        n26_adj_3863, n95, n431_adj_3864, n35975, n36779, n36886, 
        n36967, n334_adj_3867, n35974, n36966, n1707, n518, n36778, 
        n445, n36777, n36619, n36965;
    wire [23:0]n75;
    wire [23:0]n76;
    
    wire n34695, n237_adj_3872, n35973, n743_adj_3873, n36618, n47_adj_3874, 
        n140_adj_3875, n36885, n372, n36776;
    wire [25:0]n8831;
    
    wire n36357, n45_adj_3877, n34694, n36356, n646_adj_3879, n36617, 
        n878, n36355, n41830;
    wire [17:0]n8535;
    
    wire n35972, n42569, n46668, n35971, n18_adj_3883, n36964, n549_adj_3884, 
        n36616, n299_adj_3886, n36775, n452_adj_3887, n36615, n226_adj_3889, 
        n36774, n36354, n35970, n36884, n36963, n43_adj_3890, n34693, 
        n36883, n153_adj_3893, n36773, n355_adj_3894, n36614, n36353, 
        n36352, n11_adj_3895, n80_adj_3896, n258_adj_3897, n36613, 
        n36351, n36350, n36882, n68_adj_3898, n161_adj_3899, n36349, 
        n36348, n36771, n1687, n35969, n36962;
    wire [10:0]n9146;
    
    wire n36612, n36347, n36611, n36881, n36770, n36610, n36609, 
        n36961, n36880, n36769, n740_adj_3900, n36608, n643_adj_3901, 
        n36607, n36879, n36768, n35968, n546_adj_3902, n36606, n36346, 
        n449_adj_3903, n36605, n36345, n36767, n352_adj_3904, n36604, 
        n36344, n41_adj_3905, n34692, n35967, n36343, n35966, n36878, 
        n36342, n35965, n255_adj_3909, n36603, n35964, n35963, n36766, 
        n36877, n36341, n65_adj_3910, n158_adj_3911, n36340, n36339, 
        n35962, n36960, n719_adj_3912, n35961;
    wire [11:0]n9132;
    
    wire n36602, n695_adj_3913, n36338, n622_adj_3914, n35960, n598_adj_3915, 
        n36337, n525_adj_3916, n35959, n36959, n36876, n36765, n36601, 
        n501_adj_3917, n36336, n404_adj_3918, n36335, n36600, n307_adj_3919, 
        n36334, n428_adj_3920, n35958, n210_adj_3921, n36333, n331_adj_3922, 
        n35957, n234_adj_3923, n35956, n36764, n1703, n36958, n20_adj_3924, 
        n113_adj_3925, n44_adj_3926, n137_adj_3927;
    wire [18:0]n8514;
    
    wire n35955, n35954, n36763, n36599;
    wire [26:0]n8802;
    
    wire n36332, n36331, n36330, n36598, n35953, n36329, n35952, 
        n35951, n36328, n36875, n36762, n737_adj_3928, n36597, n36957, 
        n36327, n640_adj_3929, n36596, n543_adj_3930, n36595, n35950, 
        n36326, n36325, n39_adj_3931, n34691, n446_adj_3933, n36594, 
        n36761, n35949, n349_adj_3934, n36593, n36324, n36323, n252_adj_3935, 
        n36592, n36322, n35948;
    wire [24:0]n79;
    
    wire n34844, n37_adj_3937, n34690, n34843, n36321, n35_adj_3939, 
        n34689, n33_adj_3941, n34688, n34842, n35947, n36956, n36874, 
        n36760, n62_adj_3944, n155_adj_3945, n35946, n36320, n34841, 
        n34840;
    wire [12:0]n9117;
    
    wire n36591, n31_adj_3948, n34687, n36319, n34839, n29_adj_3951, 
        n34686, n36590, n34838, n34837, n35945, n36759, n27_adj_3955, 
        n34685, n36589, n34836, n36318, n36873, n36758, n36588, 
        n35944, n36317, n34835, n716_adj_3959, n35943, n25_adj_3960, 
        n34684, n34834, n36587, n36316, n34833, n36315, n619_adj_3964, 
        n35942, n23_adj_3965, n34683, n34832, n522_adj_3968, n35941, 
        n21_adj_3969, n34682, n34831, n19_adj_3972, n34681, n34830, 
        n36872, n36314, n425_adj_3975, n35940, n36757, n36871, n36586, 
        n34829, n36313, n17_adj_3977, n34680, n328_adj_3979, n35939, 
        n36756, n734_adj_3980, n36585, n637_adj_3981, n36584, n231_adj_3982, 
        n35938, n41_adj_3983, n134_adj_3984, n692_adj_3985, n36312, 
        n34828, n15_adj_3987, n34679, n595_adj_3989, n36311;
    wire [19:0]n8492;
    
    wire n35937, n36955, n540_adj_3990, n36583, n34827, n35936, 
        n13_adj_3992, n34678, n530, n36870, n498_adj_3994, n36310, 
        n515, n36755, n35935, n401_adj_3995, n36309, n35934, n443_adj_3996, 
        n36582, n35933, n34826, n35932, n11_adj_3998, n34677, n304_adj_4000, 
        n36308, n442, n36754, n346_adj_4001, n36581, n35931, n369, 
        n36753, n249_adj_4002, n36580, n34825, n35930, n35929, n9_adj_4004, 
        n34676, n34824, n207_adj_4007, n36307, n17_adj_4008, n110_adj_4009, 
        n59_adj_4010, n152_adj_4011, n35928, n36306, n35927, n36305;
    wire [13:0]n9101;
    
    wire n36579, n34823, n36304, n35926, n36578, n7_adj_4013, n34675, 
        n34822, n35925, n713_adj_4016, n35924, n457_adj_4017, n36869, 
        n36303, n36577, n36302, n296_adj_4018, n36752, n36576, n36301, 
        n36954, n36575, n34821, n36300, n223_adj_4020, n36751, n36574, 
        n384, n36868, n36573, n5_adj_4021, n34674, n150_adj_4023, 
        n36750, n1683, n36953, n616_adj_4024, n35923, n731_adj_4026, 
        n36572, n519_adj_4027, n35922, n634_adj_4028, n36571;
    wire [22:0]n1796;
    
    wire n311_adj_4029, n36867, n3_adj_4030, n34673, n36299, n537_adj_4032, 
        n36570, n36298, n36952, n36297, n8_adj_4033, n77, n36296, 
        n422_adj_4034, n35921, n440_adj_4035, n36569, n36295, n36294, 
        n325_adj_4036, n35920, n343_adj_4037, n36568, n36951, n36293, 
        n228_adj_4038, n35919, n36748, n246_adj_4039, n36567, n36292, 
        n36291, n38_adj_4040, n131_adj_4041, n238_adj_4042, n36866, 
        n56_adj_4043, n149_adj_4044, n36290, n36289, n36747, n36566, 
        n36565, n36288, n36287, n36950, n36564, n36286, n689_adj_4045, 
        n36285, n36563, n592_adj_4046, n36284, n36746, n495_adj_4047, 
        n36283, n36562, n398_adj_4048, n36282, n165_adj_4049, n36865, 
        n36745, n35918, n36561, n35917, n36560, n35916, n23_adj_4052, 
        n92, n36744, n301_adj_4053, n36281, n36949, n36559, n35915, 
        n728_adj_4054, n36558, n35914, n36743, n631_adj_4055, n36557, 
        n35913, n35912, n534_adj_4056, n36556, n36863, n36742, n35911, 
        n437_adj_4057, n36555, n35910, n340_adj_4058, n36554, n35909, 
        n36948, n36741, n204_adj_4059, n36280, n35908, n14_adj_4060, 
        n107_adj_4061, n36862, n35907, n243_adj_4062, n36553, n36279, 
        n35906, n36740, n36278, n35905, n53_adj_4063, n146_adj_4064, 
        n36277, n710_adj_4065, n35904, n36276, n36552, n36551, n613_adj_4066, 
        n35903, n36275, n516_adj_4067, n35902, n36274, n419_adj_4068, 
        n35901, n48426, n34672, n34671, n322_adj_4070, n35900, n36861, 
        n36739, n36550, n36273, n225_adj_4071, n35899, n36272, n35_adj_4072, 
        n128_adj_4073, n36271, n36549, n36947, n34670, n36738, n35898, 
        n36270, n35897, n36860, n36946, n34669, n36859, n35896, 
        n34668, n36548, n36269, n35895, n34667, n35894, n36268, 
        n36547, n35893, n36267, n36945, n35892, n36858, n35891, 
        n36546, n36266, n12_adj_4079, n43808, n8_adj_4080, n11_adj_4081, 
        n4_adj_4082, n48425, n47225, n6_adj_4085, n8_adj_4086;
    wire [5:0]GATES_5__N_3398;
    
    wire n19_adj_4088, n44318, n44314, n44316, n29_adj_4089, n6_adj_4090, 
        n46595, n6_adj_4093, n18_adj_4094, n24_adj_4095, n22_adj_4096, 
        n26_adj_4097, n43573, n11_adj_4098, n9_adj_4099, n17_adj_4100, 
        n48045, n48043, n47292, n50913, n48049, n48037, n47306, 
        n50901, n10_adj_4101, n30_adj_4102, n5_adj_4103, n48053, n48051, 
        n47324, n48347, n48815, n48039, n48606, n48922, n49040, 
        n6_adj_4104, n47368, n24_adj_4105, n48447, n47298, n50866, 
        n48463, n47680, n4_adj_4106, n48439, n48440, n8_adj_4107, 
        n47286, n6_adj_4108, n16_adj_4109, n47288, n48590, n47690, 
        n48891, n4_adj_4110, n48443, n47309, n48845, n47682, n49006, 
        n49007, n48025, n48732, n47688, n48892, n48889;
    
    SB_LUT4 add_4449_15_lut (.I0(GND_net), .I1(n8772[12]), .I2(GND_net), 
            .I3(n36264), .O(n8741[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40564_4_lut (.I0(n47706), .I1(n8), .I2(n15), .I3(n47961), 
            .O(n48467));   // verilog/motorControl.v(44[31:51])
    defparam i40564_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4432_14 (.CI(n35889), .I0(n8469[11]), .I1(GND_net), .CO(n35890));
    SB_LUT4 add_4432_13_lut (.I0(GND_net), .I1(n8469[10]), .I2(GND_net), 
            .I3(n35888), .O(n8445[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_13 (.CI(n35888), .I0(n8469[10]), .I1(GND_net), .CO(n35889));
    SB_CARRY add_4449_15 (.CI(n36264), .I0(n8772[12]), .I1(GND_net), .CO(n36265));
    SB_LUT4 add_4432_12_lut (.I0(GND_net), .I1(n8469[9]), .I2(GND_net), 
            .I3(n35887), .O(n8445[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_12 (.CI(n35887), .I0(n8469[9]), .I1(GND_net), .CO(n35888));
    SB_LUT4 add_4432_11_lut (.I0(GND_net), .I1(n8469[8]), .I2(GND_net), 
            .I3(n35886), .O(n8445[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_17_lut (.I0(GND_net), .I1(n1802[14]), .I2(GND_net), 
            .I3(n36856), .O(n1801[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_12 (.CI(n36736), .I0(n1797[9]), .I1(GND_net), 
            .CO(n36737));
    SB_CARRY add_4462_9 (.CI(n36544), .I0(n9084[6]), .I1(GND_net), .CO(n36545));
    SB_LUT4 i40565_3_lut (.I0(n48467), .I1(pwm_23__N_3310[8]), .I2(\PID_CONTROLLER.result [8]), 
            .I3(GND_net), .O(n18));   // verilog/motorControl.v(44[31:51])
    defparam i40565_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4449_14_lut (.I0(GND_net), .I1(n8772[11]), .I2(GND_net), 
            .I3(n36263), .O(n8741[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_11 (.CI(n35886), .I0(n8469[8]), .I1(GND_net), .CO(n35887));
    SB_LUT4 add_4432_10_lut (.I0(GND_net), .I1(n8469[7]), .I2(GND_net), 
            .I3(n35885), .O(n8445[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_10 (.CI(n35885), .I0(n8469[7]), .I1(GND_net), .CO(n35886));
    SB_LUT4 unary_minus_17_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n57[17]), 
            .I3(n34665), .O(pwm_23__N_3310[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_11_lut (.I0(GND_net), .I1(n1797[8]), .I2(GND_net), 
            .I3(n36735), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_8_lut (.I0(GND_net), .I1(n9084[5]), .I2(n725), .I3(n36543), 
            .O(n9066[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_9_lut (.I0(GND_net), .I1(n8469[6]), .I2(GND_net), 
            .I3(n35884), .O(n8445[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_14 (.CI(n36263), .I0(n8772[11]), .I1(GND_net), .CO(n36264));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i41_2_lut  (.I0(deadband[20]), 
            .I1(\PID_CONTROLLER.result [20]), .I2(GND_net), .I3(GND_net), 
            .O(n41));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i41_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 add_4449_13_lut (.I0(GND_net), .I1(n8772[10]), .I2(GND_net), 
            .I3(n36262), .O(n8741[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_9 (.CI(n35884), .I0(n8469[6]), .I1(GND_net), .CO(n35885));
    SB_CARRY add_4462_8 (.CI(n36543), .I0(n9084[5]), .I1(n725), .CO(n36544));
    SB_LUT4 add_4432_8_lut (.I0(GND_net), .I1(n8469[5]), .I2(n707), .I3(n35883), 
            .O(n8445[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_19 (.CI(n34665), .I0(GND_net), .I1(n57[17]), 
            .CO(n34666));
    SB_CARRY add_4432_8 (.CI(n35883), .I0(n8469[5]), .I1(n707), .CO(n35884));
    SB_CARRY add_4449_13 (.CI(n36262), .I0(n8772[10]), .I1(GND_net), .CO(n36263));
    SB_LUT4 add_4449_12_lut (.I0(GND_net), .I1(n8772[9]), .I2(GND_net), 
            .I3(n36261), .O(n8741[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_7_lut (.I0(GND_net), .I1(n9084[4]), .I2(n628), .I3(n36542), 
            .O(n9066[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_7_lut (.I0(GND_net), .I1(n8469[4]), .I2(n610), .I3(n35882), 
            .O(n8445[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_12 (.CI(n36261), .I0(n8772[9]), .I1(GND_net), .CO(n36262));
    SB_CARRY add_4432_7 (.CI(n35882), .I0(n8469[4]), .I1(n610), .CO(n35883));
    SB_LUT4 add_4432_6_lut (.I0(GND_net), .I1(n8469[3]), .I2(n513), .I3(n35881), 
            .O(n8445[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_6 (.CI(n35881), .I0(n8469[3]), .I1(n513), .CO(n35882));
    SB_LUT4 unary_minus_17_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n57[16]), 
            .I3(n34664), .O(pwm_23__N_3310[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_5_lut (.I0(GND_net), .I1(n8469[2]), .I2(n416_c), 
            .I3(n35880), .O(n8445[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_11_lut (.I0(GND_net), .I1(n8772[8]), .I2(GND_net), 
            .I3(n36260), .O(n8741[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_5 (.CI(n35880), .I0(n8469[2]), .I1(n416_c), .CO(n35881));
    SB_LUT4 add_4432_4_lut (.I0(GND_net), .I1(n8469[1]), .I2(n319), .I3(n35879), 
            .O(n8445[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_11 (.CI(n36735), .I0(n1797[8]), .I1(GND_net), 
            .CO(n36736));
    SB_CARRY add_4462_7 (.CI(n36542), .I0(n9084[4]), .I1(n628), .CO(n36543));
    SB_CARRY add_4449_11 (.CI(n36260), .I0(n8772[8]), .I1(GND_net), .CO(n36261));
    SB_CARRY add_4432_4 (.CI(n35879), .I0(n8469[1]), .I1(n319), .CO(n35880));
    SB_LUT4 add_4432_3_lut (.I0(GND_net), .I1(n8469[0]), .I2(n222), .I3(n35878), 
            .O(n8445[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_10_lut (.I0(GND_net), .I1(n8772[7]), .I2(GND_net), 
            .I3(n36259), .O(n8741[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_3 (.CI(n35878), .I0(n8469[0]), .I1(n222), .CO(n35879));
    SB_LUT4 add_4432_2_lut (.I0(GND_net), .I1(n32), .I2(n125), .I3(GND_net), 
            .O(n8445[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_6_lut (.I0(GND_net), .I1(n9084[3]), .I2(n531), .I3(n36541), 
            .O(n9066[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_10 (.CI(n36259), .I0(n8772[7]), .I1(GND_net), .CO(n36260));
    SB_CARRY add_4432_2 (.CI(GND_net), .I0(n32), .I1(n125), .CO(n35878));
    SB_CARRY mult_14_add_1216_17 (.CI(n36856), .I0(n1802[14]), .I1(GND_net), 
            .CO(n36857));
    SB_LUT4 mult_14_add_1211_10_lut (.I0(GND_net), .I1(n1797[7]), .I2(GND_net), 
            .I3(n36734), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_13_lut (.I0(GND_net), .I1(n9555[10]), .I2(GND_net), 
            .I3(n36943), .O(n9225[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_24_lut (.I0(GND_net), .I1(n8445[21]), .I2(GND_net), 
            .I3(n35877), .O(n8420[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_9_lut (.I0(GND_net), .I1(n8772[6]), .I2(GND_net), 
            .I3(n36258), .O(n8741[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_16_lut (.I0(GND_net), .I1(n1802[13]), .I2(GND_net), 
            .I3(n36855), .O(n1801[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_23_lut (.I0(GND_net), .I1(n8445[20]), .I2(GND_net), 
            .I3(n35876), .O(n8420[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_6 (.CI(n36541), .I0(n9084[3]), .I1(n531), .CO(n36542));
    SB_CARRY mult_14_add_1211_10 (.CI(n36734), .I0(n1797[7]), .I1(GND_net), 
            .CO(n36735));
    SB_CARRY add_4431_23 (.CI(n35876), .I0(n8445[20]), .I1(GND_net), .CO(n35877));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i37_2_lut  (.I0(deadband[18]), 
            .I1(\PID_CONTROLLER.result [18]), .I2(GND_net), .I3(GND_net), 
            .O(n37));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i37_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY mult_14_add_1216_16 (.CI(n36855), .I0(n1802[13]), .I1(GND_net), 
            .CO(n36856));
    SB_LUT4 add_4431_22_lut (.I0(GND_net), .I1(n8445[19]), .I2(GND_net), 
            .I3(n35875), .O(n8420[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_5_lut (.I0(GND_net), .I1(n9084[2]), .I2(n434), .I3(n36540), 
            .O(n9066[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_22 (.CI(n35875), .I0(n8445[19]), .I1(GND_net), .CO(n35876));
    SB_LUT4 mult_14_add_1211_9_lut (.I0(GND_net), .I1(n1797[6]), .I2(GND_net), 
            .I3(n36733), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_9 (.CI(n36258), .I0(n8772[6]), .I1(GND_net), .CO(n36259));
    SB_CARRY mult_14_add_1211_9 (.CI(n36733), .I0(n1797[6]), .I1(GND_net), 
            .CO(n36734));
    SB_CARRY add_4462_5 (.CI(n36540), .I0(n9084[2]), .I1(n434), .CO(n36541));
    SB_LUT4 add_4449_8_lut (.I0(GND_net), .I1(n8772[5]), .I2(n686), .I3(n36257), 
            .O(n8741[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_8_lut (.I0(GND_net), .I1(n1797[5]), .I2(n512), 
            .I3(n36732), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_21_lut (.I0(GND_net), .I1(n8445[18]), .I2(GND_net), 
            .I3(n35874), .O(n8420[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_13 (.CI(n36943), .I0(n9555[10]), .I1(GND_net), .CO(n36944));
    SB_LUT4 add_4473_12_lut (.I0(GND_net), .I1(n9555[9]), .I2(GND_net), 
            .I3(n36942), .O(n9225[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_4_lut (.I0(GND_net), .I1(n9084[1]), .I2(n337), .I3(n36539), 
            .O(n9066[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_8 (.CI(n36732), .I0(n1797[5]), .I1(n512), 
            .CO(n36733));
    SB_LUT4 mult_14_add_1216_15_lut (.I0(GND_net), .I1(n1802[12]), .I2(GND_net), 
            .I3(n36854), .O(n1801[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_12 (.CI(n36942), .I0(n9555[9]), .I1(GND_net), .CO(n36943));
    SB_LUT4 mult_14_add_1211_7_lut (.I0(GND_net), .I1(n1797[4]), .I2(n439), 
            .I3(n36731), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_4 (.CI(n36539), .I0(n9084[1]), .I1(n337), .CO(n36540));
    SB_CARRY add_4431_21 (.CI(n35874), .I0(n8445[18]), .I1(GND_net), .CO(n35875));
    SB_CARRY add_4449_8 (.CI(n36257), .I0(n8772[5]), .I1(n686), .CO(n36258));
    SB_LUT4 add_4431_20_lut (.I0(GND_net), .I1(n8445[17]), .I2(GND_net), 
            .I3(n35873), .O(n8420[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_20 (.CI(n35873), .I0(n8445[17]), .I1(GND_net), .CO(n35874));
    SB_LUT4 add_4473_11_lut (.I0(GND_net), .I1(n9555[8]), .I2(GND_net), 
            .I3(n36941), .O(n9225[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_7_lut (.I0(GND_net), .I1(n8772[4]), .I2(n589_adj_3465), 
            .I3(n36256), .O(n8741[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_19_lut (.I0(GND_net), .I1(n8445[16]), .I2(GND_net), 
            .I3(n35872), .O(n8420[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_19 (.CI(n35872), .I0(n8445[16]), .I1(GND_net), .CO(n35873));
    SB_LUT4 add_4462_3_lut (.I0(GND_net), .I1(n9084[0]), .I2(n240), .I3(n36538), 
            .O(n9066[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_11 (.CI(n36941), .I0(n9555[8]), .I1(GND_net), .CO(n36942));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i29_2_lut  (.I0(deadband[14]), 
            .I1(\PID_CONTROLLER.result [14]), .I2(GND_net), .I3(GND_net), 
            .O(n29_c));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i29_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY mult_14_add_1216_15 (.CI(n36854), .I0(n1802[12]), .I1(GND_net), 
            .CO(n36855));
    SB_CARRY add_4462_3 (.CI(n36538), .I0(n9084[0]), .I1(n240), .CO(n36539));
    SB_LUT4 add_4431_18_lut (.I0(GND_net), .I1(n8445[15]), .I2(GND_net), 
            .I3(n35871), .O(n8420[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_14_lut (.I0(GND_net), .I1(n1802[11]), .I2(GND_net), 
            .I3(n36853), .O(n1801[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i31_2_lut  (.I0(deadband[15]), 
            .I1(\PID_CONTROLLER.result [15]), .I2(GND_net), .I3(GND_net), 
            .O(n31));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i31_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY mult_14_add_1211_7 (.CI(n36731), .I0(n1797[4]), .I1(n439), 
            .CO(n36732));
    SB_CARRY add_4431_18 (.CI(n35871), .I0(n8445[15]), .I1(GND_net), .CO(n35872));
    SB_LUT4 add_4462_2_lut (.I0(GND_net), .I1(n50), .I2(n143), .I3(GND_net), 
            .O(n9066[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_7 (.CI(n36256), .I0(n8772[4]), .I1(n589_adj_3465), 
            .CO(n36257));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i7_2_lut  (.I0(deadband[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i7_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 add_4449_6_lut (.I0(GND_net), .I1(n8772[3]), .I2(n492), .I3(n36255), 
            .O(n8741[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_17_lut (.I0(GND_net), .I1(n8445[14]), .I2(GND_net), 
            .I3(n35870), .O(n8420[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_17 (.CI(n35870), .I0(n8445[14]), .I1(GND_net), .CO(n35871));
    SB_CARRY add_4449_6 (.CI(n36255), .I0(n8772[3]), .I1(n492), .CO(n36256));
    SB_CARRY mult_14_add_1216_14 (.CI(n36853), .I0(n1802[11]), .I1(GND_net), 
            .CO(n36854));
    SB_LUT4 add_4431_16_lut (.I0(GND_net), .I1(n8445[13]), .I2(GND_net), 
            .I3(n35869), .O(n8420[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_6_lut (.I0(GND_net), .I1(n1797[3]), .I2(n366), 
            .I3(n36730), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_13_lut (.I0(GND_net), .I1(n1802[10]), .I2(GND_net), 
            .I3(n36852), .O(n1801[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_2 (.CI(GND_net), .I0(n50), .I1(n143), .CO(n36538));
    SB_CARRY add_4431_16 (.CI(n35869), .I0(n8445[13]), .I1(GND_net), .CO(n35870));
    SB_CARRY mult_14_add_1211_6 (.CI(n36730), .I0(n1797[3]), .I1(n366), 
            .CO(n36731));
    SB_LUT4 add_4461_18_lut (.I0(GND_net), .I1(n9066[15]), .I2(GND_net), 
            .I3(n36537), .O(n9047[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_17_lut (.I0(GND_net), .I1(n9066[14]), .I2(GND_net), 
            .I3(n36536), .O(n9047[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_5_lut (.I0(GND_net), .I1(n1797[2]), .I2(n293), 
            .I3(n36729), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_17 (.CI(n36536), .I0(n9066[14]), .I1(GND_net), .CO(n36537));
    SB_LUT4 add_4449_5_lut (.I0(GND_net), .I1(n8772[2]), .I2(n395), .I3(n36254), 
            .O(n8741[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_5 (.CI(n36729), .I0(n1797[2]), .I1(n293), 
            .CO(n36730));
    SB_LUT4 add_4461_16_lut (.I0(GND_net), .I1(n9066[13]), .I2(GND_net), 
            .I3(n36535), .O(n9047[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_16 (.CI(n36535), .I0(n9066[13]), .I1(GND_net), .CO(n36536));
    SB_LUT4 add_4431_15_lut (.I0(GND_net), .I1(n8445[12]), .I2(GND_net), 
            .I3(n35868), .O(n8420[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_5 (.CI(n36254), .I0(n8772[2]), .I1(n395), .CO(n36255));
    SB_CARRY unary_minus_17_add_3_18 (.CI(n34664), .I0(GND_net), .I1(n57[16]), 
            .CO(n34665));
    SB_CARRY mult_14_add_1216_13 (.CI(n36852), .I0(n1802[10]), .I1(GND_net), 
            .CO(n36853));
    SB_CARRY add_4431_15 (.CI(n35868), .I0(n8445[12]), .I1(GND_net), .CO(n35869));
    SB_LUT4 add_4449_4_lut (.I0(GND_net), .I1(n8772[1]), .I2(n298), .I3(n36253), 
            .O(n8741[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_14_lut (.I0(GND_net), .I1(n8445[11]), .I2(GND_net), 
            .I3(n35867), .O(n8420[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_14 (.CI(n35867), .I0(n8445[11]), .I1(GND_net), .CO(n35868));
    SB_LUT4 add_4431_13_lut (.I0(GND_net), .I1(n8445[10]), .I2(GND_net), 
            .I3(n35866), .O(n8420[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_13 (.CI(n35866), .I0(n8445[10]), .I1(GND_net), .CO(n35867));
    SB_CARRY add_4449_4 (.CI(n36253), .I0(n8772[1]), .I1(n298), .CO(n36254));
    SB_LUT4 add_4431_12_lut (.I0(GND_net), .I1(n8445[9]), .I2(GND_net), 
            .I3(n35865), .O(n8420[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_12 (.CI(n35865), .I0(n8445[9]), .I1(GND_net), .CO(n35866));
    SB_LUT4 add_4449_3_lut (.I0(GND_net), .I1(n8772[0]), .I2(n201), .I3(n36252), 
            .O(n8741[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_11_lut (.I0(GND_net), .I1(n8445[8]), .I2(GND_net), 
            .I3(n35864), .O(n8420[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_4_lut (.I0(GND_net), .I1(n1797[1]), .I2(n220), 
            .I3(n36728), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_15_lut (.I0(GND_net), .I1(n9066[12]), .I2(GND_net), 
            .I3(n36534), .O(n9047[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_3 (.CI(n36252), .I0(n8772[0]), .I1(n201), .CO(n36253));
    SB_LUT4 add_4449_2_lut (.I0(GND_net), .I1(n11), .I2(n104), .I3(GND_net), 
            .O(n8741[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_11 (.CI(n35864), .I0(n8445[8]), .I1(GND_net), .CO(n35865));
    SB_LUT4 add_4431_10_lut (.I0(GND_net), .I1(n8445[7]), .I2(GND_net), 
            .I3(n35863), .O(n8420[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_2 (.CI(GND_net), .I0(n11), .I1(n104), .CO(n36252));
    SB_CARRY mult_14_add_1211_4 (.CI(n36728), .I0(n1797[1]), .I1(n220), 
            .CO(n36729));
    SB_LUT4 mult_12_add_2137_32_lut (.I0(n58[25]), .I1(n8709[29]), .I2(GND_net), 
            .I3(n36251), .O(n6817[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4431_10 (.CI(n35863), .I0(n8445[7]), .I1(GND_net), .CO(n35864));
    SB_LUT4 add_4431_9_lut (.I0(GND_net), .I1(n8445[6]), .I2(GND_net), 
            .I3(n35862), .O(n8420[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_15 (.CI(n36534), .I0(n9066[12]), .I1(GND_net), .CO(n36535));
    SB_LUT4 mult_12_add_2137_31_lut (.I0(GND_net), .I1(n8709[28]), .I2(GND_net), 
            .I3(n36250), .O(n191[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_9 (.CI(n35862), .I0(n8445[6]), .I1(GND_net), .CO(n35863));
    SB_LUT4 add_4431_8_lut (.I0(GND_net), .I1(n8445[5]), .I2(n704), .I3(n35861), 
            .O(n8420[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_8 (.CI(n35861), .I0(n8445[5]), .I1(n704), .CO(n35862));
    SB_LUT4 add_4431_7_lut (.I0(GND_net), .I1(n8445[4]), .I2(n607), .I3(n35860), 
            .O(n8420[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_7 (.CI(n35860), .I0(n8445[4]), .I1(n607), .CO(n35861));
    SB_CARRY mult_12_add_2137_31 (.CI(n36250), .I0(n8709[28]), .I1(GND_net), 
            .CO(n36251));
    SB_LUT4 add_4473_10_lut (.I0(GND_net), .I1(n9555[7]), .I2(GND_net), 
            .I3(n36940), .O(n9225[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_6_lut (.I0(GND_net), .I1(n8445[3]), .I2(n510), .I3(n35859), 
            .O(n8420[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_6 (.CI(n35859), .I0(n8445[3]), .I1(n510), .CO(n35860));
    SB_LUT4 mult_12_add_2137_30_lut (.I0(GND_net), .I1(n8709[27]), .I2(GND_net), 
            .I3(n36249), .O(n191[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_14_lut (.I0(GND_net), .I1(n9066[11]), .I2(GND_net), 
            .I3(n36533), .O(n9047[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_10 (.CI(n36940), .I0(n9555[7]), .I1(GND_net), .CO(n36941));
    SB_LUT4 add_4431_5_lut (.I0(GND_net), .I1(n8445[2]), .I2(n413), .I3(n35858), 
            .O(n8420[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_5 (.CI(n35858), .I0(n8445[2]), .I1(n413), .CO(n35859));
    SB_LUT4 mult_14_add_1216_12_lut (.I0(GND_net), .I1(n1802[9]), .I2(GND_net), 
            .I3(n36851), .O(n1801[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_3_lut (.I0(GND_net), .I1(n1797[0]), .I2(n147), 
            .I3(n36727), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_14 (.CI(n36533), .I0(n9066[11]), .I1(GND_net), .CO(n36534));
    SB_CARRY mult_12_add_2137_30 (.CI(n36249), .I0(n8709[27]), .I1(GND_net), 
            .CO(n36250));
    SB_LUT4 add_4461_13_lut (.I0(GND_net), .I1(n9066[10]), .I2(GND_net), 
            .I3(n36532), .O(n9047[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4431_4_lut (.I0(GND_net), .I1(n8445[1]), .I2(n316), .I3(n35857), 
            .O(n8420[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_12 (.CI(n36851), .I0(n1802[9]), .I1(GND_net), 
            .CO(n36852));
    SB_LUT4 mult_12_add_2137_29_lut (.I0(GND_net), .I1(n8709[26]), .I2(GND_net), 
            .I3(n36248), .O(n191[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_4 (.CI(n35857), .I0(n8445[1]), .I1(n316), .CO(n35858));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i33_2_lut  (.I0(deadband[16]), 
            .I1(\PID_CONTROLLER.result [16]), .I2(GND_net), .I3(GND_net), 
            .O(n33));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i33_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 add_4431_3_lut (.I0(GND_net), .I1(n8445[0]), .I2(n219_adj_3466), 
            .I3(n35856), .O(n8420[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_29 (.CI(n36248), .I0(n8709[26]), .I1(GND_net), 
            .CO(n36249));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i11_2_lut  (.I0(deadband[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3467));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i11_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY add_4431_3 (.CI(n35856), .I0(n8445[0]), .I1(n219_adj_3466), 
            .CO(n35857));
    SB_CARRY mult_14_add_1211_3 (.CI(n36727), .I0(n1797[0]), .I1(n147), 
            .CO(n36728));
    SB_LUT4 add_4473_9_lut (.I0(GND_net), .I1(n9555[6]), .I2(GND_net), 
            .I3(n36939), .O(n9225[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_13 (.CI(n36532), .I0(n9066[10]), .I1(GND_net), .CO(n36533));
    SB_LUT4 add_4431_2_lut (.I0(GND_net), .I1(n29_adj_3468), .I2(n122), 
            .I3(GND_net), .O(n8420[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4431_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_28_lut (.I0(GND_net), .I1(n8709[25]), .I2(GND_net), 
            .I3(n36247), .O(n191[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4431_2 (.CI(GND_net), .I0(n29_adj_3468), .I1(n122), .CO(n35856));
    SB_LUT4 add_4430_25_lut (.I0(GND_net), .I1(n8420[22]), .I2(GND_net), 
            .I3(n35855), .O(n8394[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_11_lut (.I0(GND_net), .I1(n1802[8]), .I2(GND_net), 
            .I3(n36850), .O(n1801[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_24_lut (.I0(GND_net), .I1(n8420[21]), .I2(GND_net), 
            .I3(n35854), .O(n8394[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_12_lut (.I0(GND_net), .I1(n9066[9]), .I2(GND_net), 
            .I3(n36531), .O(n9047[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_12 (.CI(n36531), .I0(n9066[9]), .I1(GND_net), .CO(n36532));
    SB_CARRY add_4430_24 (.CI(n35854), .I0(n8420[21]), .I1(GND_net), .CO(n35855));
    SB_CARRY mult_12_add_2137_28 (.CI(n36247), .I0(n8709[25]), .I1(GND_net), 
            .CO(n36248));
    SB_LUT4 add_4430_23_lut (.I0(GND_net), .I1(n8420[20]), .I2(GND_net), 
            .I3(n35853), .O(n8394[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_23 (.CI(n35853), .I0(n8420[20]), .I1(GND_net), .CO(n35854));
    SB_LUT4 mult_12_add_2137_27_lut (.I0(GND_net), .I1(n8709[24]), .I2(GND_net), 
            .I3(n36246), .O(n191[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_22_lut (.I0(GND_net), .I1(n8420[19]), .I2(GND_net), 
            .I3(n35852), .O(n8394[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_22 (.CI(n35852), .I0(n8420[19]), .I1(GND_net), .CO(n35853));
    SB_CARRY mult_12_add_2137_27 (.CI(n36246), .I0(n8709[24]), .I1(GND_net), 
            .CO(n36247));
    SB_LUT4 add_4430_21_lut (.I0(GND_net), .I1(n8420[18]), .I2(GND_net), 
            .I3(n35851), .O(n8394[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_26_lut (.I0(GND_net), .I1(n8709[23]), .I2(GND_net), 
            .I3(n36245), .O(n191[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_21 (.CI(n35851), .I0(n8420[18]), .I1(GND_net), .CO(n35852));
    SB_LUT4 add_4430_20_lut (.I0(GND_net), .I1(n8420[17]), .I2(GND_net), 
            .I3(n35850), .O(n8394[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_20 (.CI(n35850), .I0(n8420[17]), .I1(GND_net), .CO(n35851));
    SB_LUT4 mult_14_add_1211_2_lut (.I0(GND_net), .I1(n5_c), .I2(n74), 
            .I3(GND_net), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_19_lut (.I0(GND_net), .I1(n8420[16]), .I2(GND_net), 
            .I3(n35849), .O(n8394[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_11_lut (.I0(GND_net), .I1(n9066[8]), .I2(GND_net), 
            .I3(n36530), .O(n9047[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_2 (.CI(GND_net), .I0(n5_c), .I1(n74), .CO(n36727));
    SB_CARRY add_4461_11 (.CI(n36530), .I0(n9066[8]), .I1(GND_net), .CO(n36531));
    SB_CARRY mult_12_add_2137_26 (.CI(n36245), .I0(n8709[23]), .I1(GND_net), 
            .CO(n36246));
    SB_CARRY add_4430_19 (.CI(n35849), .I0(n8420[16]), .I1(GND_net), .CO(n35850));
    SB_LUT4 mult_12_add_2137_25_lut (.I0(GND_net), .I1(n8709[22]), .I2(GND_net), 
            .I3(n36244), .O(n191[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_18_lut (.I0(GND_net), .I1(n8420[15]), .I2(GND_net), 
            .I3(n35848), .O(n8394[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_18 (.CI(n35848), .I0(n8420[15]), .I1(GND_net), .CO(n35849));
    SB_CARRY mult_12_add_2137_25 (.CI(n36244), .I0(n8709[22]), .I1(GND_net), 
            .CO(n36245));
    SB_LUT4 add_4430_17_lut (.I0(GND_net), .I1(n8420[14]), .I2(GND_net), 
            .I3(n35847), .O(n8394[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_17 (.CI(n35847), .I0(n8420[14]), .I1(GND_net), .CO(n35848));
    SB_LUT4 mult_12_add_2137_24_lut (.I0(GND_net), .I1(n8709[21]), .I2(GND_net), 
            .I3(n36243), .O(n191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_15_lut (.I0(GND_net), .I1(n9738[12]), .I2(GND_net), 
            .I3(n36726), .O(n9722[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_10_lut (.I0(GND_net), .I1(n9066[7]), .I2(GND_net), 
            .I3(n36529), .O(n9047[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_24 (.CI(n36243), .I0(n8709[21]), .I1(GND_net), 
            .CO(n36244));
    SB_LUT4 add_4430_16_lut (.I0(GND_net), .I1(n8420[13]), .I2(GND_net), 
            .I3(n35846), .O(n8394[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_16 (.CI(n35846), .I0(n8420[13]), .I1(GND_net), .CO(n35847));
    SB_LUT4 mult_12_add_2137_23_lut (.I0(GND_net), .I1(n8709[20]), .I2(GND_net), 
            .I3(n36242), .O(n191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_15_lut (.I0(GND_net), .I1(n8420[12]), .I2(GND_net), 
            .I3(n35845), .O(n8394[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_15 (.CI(n35845), .I0(n8420[12]), .I1(GND_net), .CO(n35846));
    SB_CARRY add_4473_9 (.CI(n36939), .I0(n9555[6]), .I1(GND_net), .CO(n36940));
    SB_CARRY mult_14_add_1216_11 (.CI(n36850), .I0(n1802[8]), .I1(GND_net), 
            .CO(n36851));
    SB_LUT4 add_4783_14_lut (.I0(GND_net), .I1(n9738[11]), .I2(GND_net), 
            .I3(n36725), .O(n9722[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_10 (.CI(n36529), .I0(n9066[7]), .I1(GND_net), .CO(n36530));
    SB_CARRY mult_12_add_2137_23 (.CI(n36242), .I0(n8709[20]), .I1(GND_net), 
            .CO(n36243));
    SB_LUT4 add_4430_14_lut (.I0(GND_net), .I1(n8420[11]), .I2(GND_net), 
            .I3(n35844), .O(n8394[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_14 (.CI(n35844), .I0(n8420[11]), .I1(GND_net), .CO(n35845));
    SB_LUT4 mult_12_add_2137_22_lut (.I0(GND_net), .I1(n8709[19]), .I2(GND_net), 
            .I3(n36241), .O(n191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_13_lut (.I0(GND_net), .I1(n8420[10]), .I2(GND_net), 
            .I3(n35843), .O(n8394[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_13 (.CI(n35843), .I0(n8420[10]), .I1(GND_net), .CO(n35844));
    SB_LUT4 add_4461_9_lut (.I0(GND_net), .I1(n9066[6]), .I2(GND_net), 
            .I3(n36528), .O(n9047[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_22 (.CI(n36241), .I0(n8709[19]), .I1(GND_net), 
            .CO(n36242));
    SB_LUT4 add_4430_12_lut (.I0(GND_net), .I1(n8420[9]), .I2(GND_net), 
            .I3(n35842), .O(n8394[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_12 (.CI(n35842), .I0(n8420[9]), .I1(GND_net), .CO(n35843));
    SB_LUT4 mult_12_add_2137_21_lut (.I0(GND_net), .I1(n8709[18]), .I2(GND_net), 
            .I3(n36240), .O(n191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_11_lut (.I0(GND_net), .I1(n8420[8]), .I2(GND_net), 
            .I3(n35841), .O(n8394[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_11 (.CI(n35841), .I0(n8420[8]), .I1(GND_net), .CO(n35842));
    SB_CARRY add_4783_14 (.CI(n36725), .I0(n9738[11]), .I1(GND_net), .CO(n36726));
    SB_CARRY add_4461_9 (.CI(n36528), .I0(n9066[6]), .I1(GND_net), .CO(n36529));
    SB_CARRY mult_12_add_2137_21 (.CI(n36240), .I0(n8709[18]), .I1(GND_net), 
            .CO(n36241));
    SB_LUT4 add_4430_10_lut (.I0(GND_net), .I1(n8420[7]), .I2(GND_net), 
            .I3(n35840), .O(n8394[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_10 (.CI(n35840), .I0(n8420[7]), .I1(GND_net), .CO(n35841));
    SB_LUT4 mult_12_add_2137_20_lut (.I0(GND_net), .I1(n8709[17]), .I2(GND_net), 
            .I3(n36239), .O(n191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_9_lut (.I0(GND_net), .I1(n8420[6]), .I2(GND_net), 
            .I3(n35839), .O(n8394[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_9 (.CI(n35839), .I0(n8420[6]), .I1(GND_net), .CO(n35840));
    SB_LUT4 add_4461_8_lut (.I0(GND_net), .I1(n9066[5]), .I2(n722), .I3(n36527), 
            .O(n9047[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_20 (.CI(n36239), .I0(n8709[17]), .I1(GND_net), 
            .CO(n36240));
    SB_LUT4 add_4430_8_lut (.I0(GND_net), .I1(n8420[5]), .I2(n701), .I3(n35838), 
            .O(n8394[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_8 (.CI(n35838), .I0(n8420[5]), .I1(n701), .CO(n35839));
    SB_LUT4 mult_12_add_2137_19_lut (.I0(GND_net), .I1(n8709[16]), .I2(GND_net), 
            .I3(n36238), .O(n191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_7_lut (.I0(GND_net), .I1(n8420[4]), .I2(n604), .I3(n35837), 
            .O(n8394[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_7 (.CI(n35837), .I0(n8420[4]), .I1(n604), .CO(n35838));
    SB_LUT4 mult_14_add_1216_10_lut (.I0(GND_net), .I1(n1802[7]), .I2(GND_net), 
            .I3(n36849), .O(n1801[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_13_lut (.I0(GND_net), .I1(n9738[10]), .I2(GND_net), 
            .I3(n36724), .O(n9722[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_8 (.CI(n36527), .I0(n9066[5]), .I1(n722), .CO(n36528));
    SB_CARRY mult_12_add_2137_19 (.CI(n36238), .I0(n8709[16]), .I1(GND_net), 
            .CO(n36239));
    SB_LUT4 add_4430_6_lut (.I0(GND_net), .I1(n8420[3]), .I2(n507), .I3(n35836), 
            .O(n8394[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_6 (.CI(n35836), .I0(n8420[3]), .I1(n507), .CO(n35837));
    SB_LUT4 mult_12_add_2137_18_lut (.I0(GND_net), .I1(n8709[15]), .I2(GND_net), 
            .I3(n36237), .O(n191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_5_lut (.I0(GND_net), .I1(n8420[2]), .I2(n410_c), 
            .I3(n35835), .O(n8394[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_5 (.CI(n35835), .I0(n8420[2]), .I1(n410_c), .CO(n35836));
    SB_LUT4 add_4461_7_lut (.I0(GND_net), .I1(n9066[4]), .I2(n625), .I3(n36526), 
            .O(n9047[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_18 (.CI(n36237), .I0(n8709[15]), .I1(GND_net), 
            .CO(n36238));
    SB_LUT4 add_4430_4_lut (.I0(GND_net), .I1(n8420[1]), .I2(n313_adj_3473), 
            .I3(n35834), .O(n8394[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_4 (.CI(n35834), .I0(n8420[1]), .I1(n313_adj_3473), 
            .CO(n35835));
    SB_LUT4 mult_12_add_2137_17_lut (.I0(GND_net), .I1(n8709[14]), .I2(GND_net), 
            .I3(n36236), .O(n191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4430_3_lut (.I0(GND_net), .I1(n8420[0]), .I2(n216), .I3(n35833), 
            .O(n8394[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_3 (.CI(n35833), .I0(n8420[0]), .I1(n216), .CO(n35834));
    SB_CARRY add_4783_13 (.CI(n36724), .I0(n9738[10]), .I1(GND_net), .CO(n36725));
    SB_CARRY add_4461_7 (.CI(n36526), .I0(n9066[4]), .I1(n625), .CO(n36527));
    SB_CARRY mult_12_add_2137_17 (.CI(n36236), .I0(n8709[14]), .I1(GND_net), 
            .CO(n36237));
    SB_LUT4 add_4430_2_lut (.I0(GND_net), .I1(n26_c), .I2(n119), .I3(GND_net), 
            .O(n8394[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4430_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_16_lut (.I0(GND_net), .I1(n8709[13]), .I2(GND_net), 
            .I3(n36235), .O(n191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4430_2 (.CI(GND_net), .I0(n26_c), .I1(n119), .CO(n35833));
    SB_LUT4 add_4429_26_lut (.I0(GND_net), .I1(n8394[23]), .I2(GND_net), 
            .I3(n35832), .O(n8367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_6_lut (.I0(GND_net), .I1(n9066[3]), .I2(n528), .I3(n36525), 
            .O(n9047[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_16 (.CI(n36235), .I0(n8709[13]), .I1(GND_net), 
            .CO(n36236));
    SB_LUT4 add_4429_25_lut (.I0(GND_net), .I1(n8394[22]), .I2(GND_net), 
            .I3(n35831), .O(n8367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_15_lut (.I0(GND_net), .I1(n8709[12]), .I2(GND_net), 
            .I3(n36234), .O(n191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_25 (.CI(n35831), .I0(n8394[22]), .I1(GND_net), .CO(n35832));
    SB_LUT4 add_4429_24_lut (.I0(GND_net), .I1(n8394[21]), .I2(GND_net), 
            .I3(n35830), .O(n8367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_8_lut (.I0(GND_net), .I1(n9555[5]), .I2(n545), .I3(n36938), 
            .O(n9225[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_10 (.CI(n36849), .I0(n1802[7]), .I1(GND_net), 
            .CO(n36850));
    SB_LUT4 add_4783_12_lut (.I0(GND_net), .I1(n9738[9]), .I2(GND_net), 
            .I3(n36723), .O(n9722[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_6 (.CI(n36525), .I0(n9066[3]), .I1(n528), .CO(n36526));
    SB_CARRY mult_12_add_2137_15 (.CI(n36234), .I0(n8709[12]), .I1(GND_net), 
            .CO(n36235));
    SB_CARRY add_4429_24 (.CI(n35830), .I0(n8394[21]), .I1(GND_net), .CO(n35831));
    SB_LUT4 add_4429_23_lut (.I0(GND_net), .I1(n8394[20]), .I2(GND_net), 
            .I3(n35829), .O(n8367[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_14_lut (.I0(GND_net), .I1(n8709[11]), .I2(GND_net), 
            .I3(n36233), .O(n191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_23 (.CI(n35829), .I0(n8394[20]), .I1(GND_net), .CO(n35830));
    SB_LUT4 add_4429_22_lut (.I0(GND_net), .I1(n8394[19]), .I2(GND_net), 
            .I3(n35828), .O(n8367[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_5_lut (.I0(GND_net), .I1(n9066[2]), .I2(n431), .I3(n36524), 
            .O(n9047[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_14 (.CI(n36233), .I0(n8709[11]), .I1(GND_net), 
            .CO(n36234));
    SB_CARRY add_4429_22 (.CI(n35828), .I0(n8394[19]), .I1(GND_net), .CO(n35829));
    SB_LUT4 add_4429_21_lut (.I0(GND_net), .I1(n8394[18]), .I2(GND_net), 
            .I3(n35827), .O(n8367[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_13_lut (.I0(GND_net), .I1(n8709[10]), .I2(GND_net), 
            .I3(n36232), .O(n191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_21 (.CI(n35827), .I0(n8394[18]), .I1(GND_net), .CO(n35828));
    SB_LUT4 add_4429_20_lut (.I0(GND_net), .I1(n8394[17]), .I2(GND_net), 
            .I3(n35826), .O(n8367[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4783_12 (.CI(n36723), .I0(n9738[9]), .I1(GND_net), .CO(n36724));
    SB_CARRY add_4461_5 (.CI(n36524), .I0(n9066[2]), .I1(n431), .CO(n36525));
    SB_CARRY mult_12_add_2137_13 (.CI(n36232), .I0(n8709[10]), .I1(GND_net), 
            .CO(n36233));
    SB_CARRY add_4429_20 (.CI(n35826), .I0(n8394[17]), .I1(GND_net), .CO(n35827));
    SB_LUT4 add_4429_19_lut (.I0(GND_net), .I1(n8394[16]), .I2(GND_net), 
            .I3(n35825), .O(n8367[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_12_lut (.I0(GND_net), .I1(n8709[9]), .I2(GND_net), 
            .I3(n36231), .O(n191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_19 (.CI(n35825), .I0(n8394[16]), .I1(GND_net), .CO(n35826));
    SB_LUT4 add_4429_18_lut (.I0(GND_net), .I1(n8394[15]), .I2(GND_net), 
            .I3(n35824), .O(n8367[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n57[15]), 
            .I3(n34663), .O(pwm_23__N_3310[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_4_lut (.I0(GND_net), .I1(n9066[1]), .I2(n334), .I3(n36523), 
            .O(n9047[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_12 (.CI(n36231), .I0(n8709[9]), .I1(GND_net), 
            .CO(n36232));
    SB_CARRY add_4429_18 (.CI(n35824), .I0(n8394[15]), .I1(GND_net), .CO(n35825));
    SB_LUT4 add_4429_17_lut (.I0(GND_net), .I1(n8394[14]), .I2(GND_net), 
            .I3(n35823), .O(n8367[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_11_lut (.I0(GND_net), .I1(n8709[8]), .I2(GND_net), 
            .I3(n36230), .O(n191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_17 (.CI(n35823), .I0(n8394[14]), .I1(GND_net), .CO(n35824));
    SB_LUT4 add_4429_16_lut (.I0(GND_net), .I1(n8394[13]), .I2(GND_net), 
            .I3(n35822), .O(n8367[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_17 (.CI(n34663), .I0(GND_net), .I1(n57[15]), 
            .CO(n34664));
    SB_LUT4 mult_14_add_1216_9_lut (.I0(GND_net), .I1(n1802[6]), .I2(GND_net), 
            .I3(n36848), .O(n1801[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_11_lut (.I0(GND_net), .I1(n9738[8]), .I2(GND_net), 
            .I3(n36722), .O(n9722[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_4 (.CI(n36523), .I0(n9066[1]), .I1(n334), .CO(n36524));
    SB_CARRY mult_12_add_2137_11 (.CI(n36230), .I0(n8709[8]), .I1(GND_net), 
            .CO(n36231));
    SB_CARRY add_4429_16 (.CI(n35822), .I0(n8394[13]), .I1(GND_net), .CO(n35823));
    SB_LUT4 add_4429_15_lut (.I0(GND_net), .I1(n8394[12]), .I2(GND_net), 
            .I3(n35821), .O(n8367[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_10_lut (.I0(GND_net), .I1(n8709[7]), .I2(GND_net), 
            .I3(n36229), .O(n191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_15 (.CI(n35821), .I0(n8394[12]), .I1(GND_net), .CO(n35822));
    SB_LUT4 add_4429_14_lut (.I0(GND_net), .I1(n8394[11]), .I2(GND_net), 
            .I3(n35820), .O(n8367[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n57[14]), 
            .I3(n34662), .O(pwm_23__N_3310[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_3_lut (.I0(GND_net), .I1(n9066[0]), .I2(n237_adj_3476), 
            .I3(n36522), .O(n9047[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_10 (.CI(n36229), .I0(n8709[7]), .I1(GND_net), 
            .CO(n36230));
    SB_CARRY add_4429_14 (.CI(n35820), .I0(n8394[11]), .I1(GND_net), .CO(n35821));
    SB_LUT4 add_4429_13_lut (.I0(GND_net), .I1(n8394[10]), .I2(GND_net), 
            .I3(n35819), .O(n8367[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_9_lut (.I0(GND_net), .I1(n8709[6]), .I2(GND_net), 
            .I3(n36228), .O(n191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_13 (.CI(n35819), .I0(n8394[10]), .I1(GND_net), .CO(n35820));
    SB_LUT4 add_4429_12_lut (.I0(GND_net), .I1(n8394[9]), .I2(GND_net), 
            .I3(n35818), .O(n8367[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_16 (.CI(n34662), .I0(GND_net), .I1(n57[14]), 
            .CO(n34663));
    SB_CARRY add_4783_11 (.CI(n36722), .I0(n9738[8]), .I1(GND_net), .CO(n36723));
    SB_CARRY add_4461_3 (.CI(n36522), .I0(n9066[0]), .I1(n237_adj_3476), 
            .CO(n36523));
    SB_CARRY mult_12_add_2137_9 (.CI(n36228), .I0(n8709[6]), .I1(GND_net), 
            .CO(n36229));
    SB_CARRY add_4429_12 (.CI(n35818), .I0(n8394[9]), .I1(GND_net), .CO(n35819));
    SB_LUT4 add_4429_11_lut (.I0(GND_net), .I1(n8394[8]), .I2(GND_net), 
            .I3(n35817), .O(n8367[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_8_lut (.I0(GND_net), .I1(n8709[5]), .I2(n680), 
            .I3(n36227), .O(n191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_11 (.CI(n35817), .I0(n8394[8]), .I1(GND_net), .CO(n35818));
    SB_LUT4 add_4429_10_lut (.I0(GND_net), .I1(n8394[7]), .I2(GND_net), 
            .I3(n35816), .O(n8367[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n57[13]), 
            .I3(n34661), .O(pwm_23__N_3310[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4461_2_lut (.I0(GND_net), .I1(n47), .I2(n140), .I3(GND_net), 
            .O(n9047[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4461_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n452));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_12_add_2137_8 (.CI(n36227), .I0(n8709[5]), .I1(n680), 
            .CO(n36228));
    SB_CARRY add_4429_10 (.CI(n35816), .I0(n8394[7]), .I1(GND_net), .CO(n35817));
    SB_LUT4 add_4429_9_lut (.I0(GND_net), .I1(n8394[6]), .I2(GND_net), 
            .I3(n35815), .O(n8367[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_7_lut (.I0(GND_net), .I1(n8709[4]), .I2(n583), 
            .I3(n36226), .O(n191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_9 (.CI(n35815), .I0(n8394[6]), .I1(GND_net), .CO(n35816));
    SB_LUT4 add_4429_8_lut (.I0(GND_net), .I1(n8394[5]), .I2(n698), .I3(n35814), 
            .O(n8367[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_15 (.CI(n34661), .I0(GND_net), .I1(n57[13]), 
            .CO(n34662));
    SB_CARRY add_4473_8 (.CI(n36938), .I0(n9555[5]), .I1(n545), .CO(n36939));
    SB_CARRY mult_14_add_1216_9 (.CI(n36848), .I0(n1802[6]), .I1(GND_net), 
            .CO(n36849));
    SB_LUT4 add_4783_10_lut (.I0(GND_net), .I1(n9738[7]), .I2(GND_net), 
            .I3(n36721), .O(n9722[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4461_2 (.CI(GND_net), .I0(n47), .I1(n140), .CO(n36522));
    SB_CARRY mult_12_add_2137_7 (.CI(n36226), .I0(n8709[4]), .I1(n583), 
            .CO(n36227));
    SB_CARRY add_4429_8 (.CI(n35814), .I0(n8394[5]), .I1(n698), .CO(n35815));
    SB_LUT4 add_4429_7_lut (.I0(GND_net), .I1(n8394[4]), .I2(n601_adj_3478), 
            .I3(n35813), .O(n8367[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_6_lut (.I0(GND_net), .I1(n8709[3]), .I2(n486), 
            .I3(n36225), .O(n191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_7 (.CI(n35813), .I0(n8394[4]), .I1(n601_adj_3478), 
            .CO(n35814));
    SB_LUT4 add_4429_6_lut (.I0(GND_net), .I1(n8394[3]), .I2(n504), .I3(n35812), 
            .O(n8367[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n57[12]), 
            .I3(n34660), .O(pwm_23__N_3310[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_14 (.CI(n34660), .I0(GND_net), .I1(n57[12]), 
            .CO(n34661));
    SB_LUT4 add_4460_19_lut (.I0(GND_net), .I1(n9047[16]), .I2(GND_net), 
            .I3(n36521), .O(n9027[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_6 (.CI(n36225), .I0(n8709[3]), .I1(n486), 
            .CO(n36226));
    SB_CARRY add_4429_6 (.CI(n35812), .I0(n8394[3]), .I1(n504), .CO(n35813));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i15_2_lut  (.I0(deadband[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3479));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i15_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 add_4429_5_lut (.I0(GND_net), .I1(n8394[2]), .I2(n407_c), 
            .I3(n35811), .O(n8367[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_5_lut (.I0(GND_net), .I1(n8709[2]), .I2(n389), 
            .I3(n36224), .O(n191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_5 (.CI(n35811), .I0(n8394[2]), .I1(n407_c), .CO(n35812));
    SB_LUT4 add_4429_4_lut (.I0(GND_net), .I1(n8394[1]), .I2(n310_adj_3480), 
            .I3(n35810), .O(n8367[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n57[11]), 
            .I3(n34659), .O(pwm_23__N_3310[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_13 (.CI(n34659), .I0(GND_net), .I1(n57[11]), 
            .CO(n34660));
    SB_CARRY add_4783_10 (.CI(n36721), .I0(n9738[7]), .I1(GND_net), .CO(n36722));
    SB_LUT4 add_4460_18_lut (.I0(GND_net), .I1(n9047[15]), .I2(GND_net), 
            .I3(n36520), .O(n9027[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_5 (.CI(n36224), .I0(n8709[2]), .I1(n389), 
            .CO(n36225));
    SB_CARRY add_4429_4 (.CI(n35810), .I0(n8394[1]), .I1(n310_adj_3480), 
            .CO(n35811));
    SB_LUT4 add_4429_3_lut (.I0(GND_net), .I1(n8394[0]), .I2(n213), .I3(n35809), 
            .O(n8367[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_4_lut (.I0(GND_net), .I1(n8709[1]), .I2(n292), 
            .I3(n36223), .O(n191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_3 (.CI(n35809), .I0(n8394[0]), .I1(n213), .CO(n35810));
    SB_LUT4 add_4429_2_lut (.I0(GND_net), .I1(n23), .I2(n116), .I3(GND_net), 
            .O(n8367[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n57[10]), 
            .I3(n34658), .O(\pwm_23__N_3310[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_12 (.CI(n34658), .I0(GND_net), .I1(n57[10]), 
            .CO(n34659));
    SB_CARRY add_4460_18 (.CI(n36520), .I0(n9047[15]), .I1(GND_net), .CO(n36521));
    SB_CARRY mult_12_add_2137_4 (.CI(n36223), .I0(n8709[1]), .I1(n292), 
            .CO(n36224));
    SB_CARRY add_4429_2 (.CI(GND_net), .I0(n23), .I1(n116), .CO(n35809));
    SB_LUT4 add_4428_27_lut (.I0(GND_net), .I1(n8367[24]), .I2(GND_net), 
            .I3(n35808), .O(n8339[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_3_lut (.I0(GND_net), .I1(n8709[0]), .I2(n195), 
            .I3(n36222), .O(n191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_26_lut (.I0(GND_net), .I1(n8367[23]), .I2(GND_net), 
            .I3(n35807), .O(n8339[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_26 (.CI(n35807), .I0(n8367[23]), .I1(GND_net), .CO(n35808));
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n57[9]), 
            .I3(n34657), .O(pwm_23__N_3310[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_11 (.CI(n34657), .I0(GND_net), .I1(n57[9]), 
            .CO(n34658));
    SB_LUT4 mult_14_add_1216_8_lut (.I0(GND_net), .I1(n1802[5]), .I2(n527), 
            .I3(n36847), .O(n1801[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_9_lut (.I0(GND_net), .I1(n9738[6]), .I2(GND_net), 
            .I3(n36720), .O(n9722[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_17_lut (.I0(GND_net), .I1(n9047[14]), .I2(GND_net), 
            .I3(n36519), .O(n9027[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_3 (.CI(n36222), .I0(n8709[0]), .I1(n195), 
            .CO(n36223));
    SB_LUT4 add_4428_25_lut (.I0(GND_net), .I1(n8367[22]), .I2(GND_net), 
            .I3(n35806), .O(n8339[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_25 (.CI(n35806), .I0(n8367[22]), .I1(GND_net), .CO(n35807));
    SB_LUT4 mult_12_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3483), .I2(n98), 
            .I3(GND_net), .O(n191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_24_lut (.I0(GND_net), .I1(n8367[21]), .I2(GND_net), 
            .I3(n35805), .O(n8339[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_24 (.CI(n35805), .I0(n8367[21]), .I1(GND_net), .CO(n35806));
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n57[8]), 
            .I3(n34656), .O(pwm_23__N_3310[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_10 (.CI(n34656), .I0(GND_net), .I1(n57[8]), 
            .CO(n34657));
    SB_CARRY add_4460_17 (.CI(n36519), .I0(n9047[14]), .I1(GND_net), .CO(n36520));
    SB_CARRY mult_12_add_2137_2 (.CI(GND_net), .I0(n5_adj_3483), .I1(n98), 
            .CO(n36222));
    SB_LUT4 add_4428_23_lut (.I0(GND_net), .I1(n8367[20]), .I2(GND_net), 
            .I3(n35804), .O(n8339[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_23 (.CI(n35804), .I0(n8367[20]), .I1(GND_net), .CO(n35805));
    SB_LUT4 add_4767_21_lut (.I0(GND_net), .I1(n9591[18]), .I2(GND_net), 
            .I3(n36221), .O(n9555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_22_lut (.I0(GND_net), .I1(n8367[19]), .I2(GND_net), 
            .I3(n35803), .O(n8339[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_22 (.CI(n35803), .I0(n8367[19]), .I1(GND_net), .CO(n35804));
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n57[7]), 
            .I3(n34655), .O(pwm_23__N_3310[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_9 (.CI(n34655), .I0(GND_net), .I1(n57[7]), 
            .CO(n34656));
    SB_CARRY add_4783_9 (.CI(n36720), .I0(n9738[6]), .I1(GND_net), .CO(n36721));
    SB_LUT4 add_4460_16_lut (.I0(GND_net), .I1(n9047[13]), .I2(GND_net), 
            .I3(n36518), .O(n9027[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_20_lut (.I0(GND_net), .I1(n9591[17]), .I2(GND_net), 
            .I3(n36220), .O(n9555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_21_lut (.I0(GND_net), .I1(n8367[18]), .I2(GND_net), 
            .I3(n35802), .O(n8339[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_20 (.CI(n36220), .I0(n9591[17]), .I1(GND_net), .CO(n36221));
    SB_CARRY add_4428_21 (.CI(n35802), .I0(n8367[18]), .I1(GND_net), .CO(n35803));
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n57[6]), 
            .I3(n34654), .O(\pwm_23__N_3310[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_20_lut (.I0(GND_net), .I1(n8367[17]), .I2(GND_net), 
            .I3(n35801), .O(n8339[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_8 (.CI(n34654), .I0(GND_net), .I1(n57[6]), 
            .CO(n34655));
    SB_CARRY add_4460_16 (.CI(n36518), .I0(n9047[13]), .I1(GND_net), .CO(n36519));
    SB_LUT4 add_4767_19_lut (.I0(GND_net), .I1(n9591[16]), .I2(GND_net), 
            .I3(n36219), .O(n9555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_20 (.CI(n35801), .I0(n8367[17]), .I1(GND_net), .CO(n35802));
    SB_CARRY add_4767_19 (.CI(n36219), .I0(n9591[16]), .I1(GND_net), .CO(n36220));
    SB_LUT4 add_4428_19_lut (.I0(GND_net), .I1(n8367[16]), .I2(GND_net), 
            .I3(n35800), .O(n8339[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_19 (.CI(n35800), .I0(n8367[16]), .I1(GND_net), .CO(n35801));
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n57[5]), 
            .I3(n34653), .O(pwm_23__N_3310[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_7_lut (.I0(GND_net), .I1(n9555[4]), .I2(n472), .I3(n36937), 
            .O(n9225[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_8 (.CI(n36847), .I0(n1802[5]), .I1(n527), 
            .CO(n36848));
    SB_LUT4 add_4783_8_lut (.I0(GND_net), .I1(n9738[5]), .I2(n545), .I3(n36719), 
            .O(n9722[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_15_lut (.I0(GND_net), .I1(n9047[12]), .I2(GND_net), 
            .I3(n36517), .O(n9027[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_18_lut (.I0(GND_net), .I1(n9591[15]), .I2(GND_net), 
            .I3(n36218), .O(n9555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_18_lut (.I0(GND_net), .I1(n8367[15]), .I2(GND_net), 
            .I3(n35799), .O(n8339[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_18 (.CI(n35799), .I0(n8367[15]), .I1(GND_net), .CO(n35800));
    SB_CARRY add_4767_18 (.CI(n36218), .I0(n9591[15]), .I1(GND_net), .CO(n36219));
    SB_LUT4 add_4428_17_lut (.I0(GND_net), .I1(n8367[14]), .I2(GND_net), 
            .I3(n35798), .O(n8339[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_17 (.CI(n35798), .I0(n8367[14]), .I1(GND_net), .CO(n35799));
    SB_CARRY add_4460_15 (.CI(n36517), .I0(n9047[12]), .I1(GND_net), .CO(n36518));
    SB_LUT4 add_4767_17_lut (.I0(GND_net), .I1(n9591[14]), .I2(GND_net), 
            .I3(n36217), .O(n9555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_16_lut (.I0(GND_net), .I1(n8367[13]), .I2(GND_net), 
            .I3(n35797), .O(n8339[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_16 (.CI(n35797), .I0(n8367[13]), .I1(GND_net), .CO(n35798));
    SB_CARRY add_4767_17 (.CI(n36217), .I0(n9591[14]), .I1(GND_net), .CO(n36218));
    SB_LUT4 add_4428_15_lut (.I0(GND_net), .I1(n8367[12]), .I2(GND_net), 
            .I3(n35796), .O(n8339[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_15 (.CI(n35796), .I0(n8367[12]), .I1(GND_net), .CO(n35797));
    SB_CARRY add_4783_8 (.CI(n36719), .I0(n9738[5]), .I1(n545), .CO(n36720));
    SB_LUT4 add_4460_14_lut (.I0(GND_net), .I1(n9047[11]), .I2(GND_net), 
            .I3(n36516), .O(n9027[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_16_lut (.I0(GND_net), .I1(n9591[13]), .I2(GND_net), 
            .I3(n36216), .O(n9555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_14_lut (.I0(GND_net), .I1(n8367[11]), .I2(GND_net), 
            .I3(n35795), .O(n8339[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i45_2_lut  (.I0(deadband[22]), 
            .I1(\PID_CONTROLLER.result [22]), .I2(GND_net), .I3(GND_net), 
            .O(n45));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i45_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY add_4428_14 (.CI(n35795), .I0(n8367[11]), .I1(GND_net), .CO(n35796));
    SB_CARRY add_4767_16 (.CI(n36216), .I0(n9591[13]), .I1(GND_net), .CO(n36217));
    SB_LUT4 add_4428_13_lut (.I0(GND_net), .I1(n8367[10]), .I2(GND_net), 
            .I3(n35794), .O(n8339[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_13 (.CI(n35794), .I0(n8367[10]), .I1(GND_net), .CO(n35795));
    SB_CARRY unary_minus_17_add_3_7 (.CI(n34653), .I0(GND_net), .I1(n57[5]), 
            .CO(n34654));
    SB_CARRY add_4460_14 (.CI(n36516), .I0(n9047[11]), .I1(GND_net), .CO(n36517));
    SB_LUT4 add_4767_15_lut (.I0(GND_net), .I1(n9591[12]), .I2(GND_net), 
            .I3(n36215), .O(n9555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_12_lut (.I0(GND_net), .I1(n8367[9]), .I2(GND_net), 
            .I3(n35793), .O(n8339[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_12 (.CI(n35793), .I0(n8367[9]), .I1(GND_net), .CO(n35794));
    SB_CARRY add_4767_15 (.CI(n36215), .I0(n9591[12]), .I1(GND_net), .CO(n36216));
    SB_LUT4 add_4428_11_lut (.I0(GND_net), .I1(n8367[8]), .I2(GND_net), 
            .I3(n35792), .O(n8339[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_11 (.CI(n35792), .I0(n8367[8]), .I1(GND_net), .CO(n35793));
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n57[4]), 
            .I3(n34652), .O(\pwm_23__N_3310[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_7_lut (.I0(GND_net), .I1(n1802[4]), .I2(n454), 
            .I3(n36846), .O(n1801[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_7_lut (.I0(GND_net), .I1(n9738[4]), .I2(n472), .I3(n36718), 
            .O(n9722[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_13_lut (.I0(GND_net), .I1(n9047[10]), .I2(GND_net), 
            .I3(n36515), .O(n9027[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_14_lut (.I0(GND_net), .I1(n9591[11]), .I2(GND_net), 
            .I3(n36214), .O(n9555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_10_lut (.I0(GND_net), .I1(n8367[7]), .I2(GND_net), 
            .I3(n35791), .O(n8339[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_10 (.CI(n35791), .I0(n8367[7]), .I1(GND_net), .CO(n35792));
    SB_CARRY add_4767_14 (.CI(n36214), .I0(n9591[11]), .I1(GND_net), .CO(n36215));
    SB_LUT4 add_4428_9_lut (.I0(GND_net), .I1(n8367[6]), .I2(GND_net), 
            .I3(n35790), .O(n8339[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_9 (.CI(n35790), .I0(n8367[6]), .I1(GND_net), .CO(n35791));
    SB_CARRY unary_minus_17_add_3_6 (.CI(n34652), .I0(GND_net), .I1(n57[4]), 
            .CO(n34653));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i17_2_lut  (.I0(deadband[8]), .I1(\PID_CONTROLLER.result [8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3486));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i17_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY add_4783_7 (.CI(n36718), .I0(n9738[4]), .I1(n472), .CO(n36719));
    SB_LUT4 add_4767_13_lut (.I0(GND_net), .I1(n9591[10]), .I2(GND_net), 
            .I3(n36213), .O(n9555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4460_13 (.CI(n36515), .I0(n9047[10]), .I1(GND_net), .CO(n36516));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i19_2_lut  (.I0(deadband[9]), .I1(\PID_CONTROLLER.result [9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3487));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i19_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i43_2_lut  (.I0(deadband[21]), 
            .I1(\PID_CONTROLLER.result [21]), .I2(GND_net), .I3(GND_net), 
            .O(n43));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i43_2_lut .LUT_INIT = 16'h6666;
    SB_CARRY add_4767_13 (.CI(n36213), .I0(n9591[10]), .I1(GND_net), .CO(n36214));
    SB_LUT4 LessThan_20_i41_2_lut (.I0(PWMLimit[20]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3488));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i39_2_lut (.I0(PWMLimit[19]), .I1(\PID_CONTROLLER.result[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n39_c));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4460_12_lut (.I0(GND_net), .I1(n9047[9]), .I2(GND_net), 
            .I3(n36514), .O(n9027[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_8_lut (.I0(GND_net), .I1(n8367[5]), .I2(n695), .I3(n35789), 
            .O(n8339[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i45_2_lut (.I0(PWMLimit[22]), .I1(\PID_CONTROLLER.result [22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_3489));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4428_8 (.CI(n35789), .I0(n8367[5]), .I1(n695), .CO(n35790));
    SB_LUT4 LessThan_20_i43_2_lut (.I0(PWMLimit[21]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_3490));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i37_2_lut (.I0(PWMLimit[18]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3491));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i23_2_lut (.I0(PWMLimit[11]), .I1(\PID_CONTROLLER.result [11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3492));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i25_2_lut (.I0(PWMLimit[12]), .I1(\PID_CONTROLLER.result [12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3493));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i25_2_lut.LUT_INIT = 16'h6666;
    SB_DFF pwm__i23 (.Q(pwm[23]), .C(clk32MHz), .D(n18644));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i22 (.Q(pwm[22]), .C(clk32MHz), .D(n18643));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i21 (.Q(pwm[21]), .C(clk32MHz), .D(n18642));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i20 (.Q(pwm[20]), .C(clk32MHz), .D(n18641));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i19 (.Q(pwm[19]), .C(clk32MHz), .D(n18640));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i18 (.Q(pwm[18]), .C(clk32MHz), .D(n18639));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i17 (.Q(pwm[17]), .C(clk32MHz), .D(n18638));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i16 (.Q(pwm[16]), .C(clk32MHz), .D(n18637));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i15 (.Q(pwm[15]), .C(clk32MHz), .D(n18636));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i14 (.Q(pwm[14]), .C(clk32MHz), .D(n18635));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i13 (.Q(pwm[13]), .C(clk32MHz), .D(n18634));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i12 (.Q(pwm[12]), .C(clk32MHz), .D(n18633));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i11 (.Q(pwm[11]), .C(clk32MHz), .D(n18632));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 sub_11_inv_0_i24_1_lut (.I0(\PID_CONTROLLER.err[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[23]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm__i10 (.Q(pwm[10]), .C(clk32MHz), .D(n18631));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i9 (.Q(pwm[9]), .C(clk32MHz), .D(n18630));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i8 (.Q(pwm[8]), .C(clk32MHz), .D(n18629));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i7 (.Q(pwm[7]), .C(clk32MHz), .D(n18628));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i6 (.Q(pwm[6]), .C(clk32MHz), .D(n18627));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i5 (.Q(pwm[5]), .C(clk32MHz), .D(n18626));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i4 (.Q(pwm[4]), .C(clk32MHz), .D(n18625));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i3 (.Q(pwm[3]), .C(clk32MHz), .D(n18624));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i2 (.Q(pwm[2]), .C(clk32MHz), .D(n18623));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 LessThan_20_i29_2_lut (.I0(PWMLimit[14]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3494));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[0]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm__i1 (.Q(pwm[1]), .C(clk32MHz), .D(n18622));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 LessThan_20_i31_2_lut (.I0(PWMLimit[15]), .I1(\PID_CONTROLLER.result [15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_3496));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i35_2_lut (.I0(PWMLimit[17]), .I1(\PID_CONTROLLER.result[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_c));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i33_2_lut (.I0(PWMLimit[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_3497));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4460_12 (.CI(n36514), .I0(n9047[9]), .I1(GND_net), .CO(n36515));
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n549));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_DFF pwm__i0 (.Q(pwm[0]), .C(clk32MHz), .D(n18574));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_10_i434_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n646));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4460_11_lut (.I0(GND_net), .I1(n9047[8]), .I2(GND_net), 
            .I3(n36513), .O(n9027[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4428_7_lut (.I0(GND_net), .I1(n8367[4]), .I2(n598), .I3(n35788), 
            .O(n8339[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_12_lut (.I0(GND_net), .I1(n9591[9]), .I2(GND_net), 
            .I3(n36212), .O(n9555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_7 (.CI(n35788), .I0(n8367[4]), .I1(n598), .CO(n35789));
    SB_LUT4 add_4428_6_lut (.I0(GND_net), .I1(n8367[3]), .I2(n501), .I3(n35787), 
            .O(n8339[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(PWMLimit[8]), .I1(\PID_CONTROLLER.result [8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3498));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(PWMLimit[9]), .I1(\PID_CONTROLLER.result [9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3499));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(PWMLimit[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3500));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[1]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(PWMLimit[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3502));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i499_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39248_4_lut (.I0(n21), .I1(n19_adj_3499), .I2(n17_adj_3498), 
            .I3(n9), .O(n47150));
    defparam i39248_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_11_inv_0_i32_1_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[26]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39242_4_lut (.I0(n27), .I1(n15_adj_3502), .I2(n13), .I3(n11_adj_3500), 
            .O(n47144));
    defparam i39242_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4767_12 (.CI(n36212), .I0(n9591[9]), .I1(GND_net), .CO(n36213));
    SB_LUT4 mult_10_i111_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4428_6 (.CI(n35787), .I0(n8367[3]), .I1(n501), .CO(n35788));
    SB_LUT4 mult_10_i48_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n71));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i48_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.err_prev__i25  (.Q(\PID_CONTROLLER.err_prev[31] ), 
           .C(clk32MHz), .D(n18495));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i24  (.Q(\PID_CONTROLLER.err_prev[23] ), 
           .C(clk32MHz), .D(n18494));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i23  (.Q(\PID_CONTROLLER.err_prev[22] ), 
           .C(clk32MHz), .D(n18493));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[2]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.err_prev__i22  (.Q(\PID_CONTROLLER.err_prev[21] ), 
           .C(clk32MHz), .D(n18492));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i21  (.Q(\PID_CONTROLLER.err_prev[20] ), 
           .C(clk32MHz), .D(n18491));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i20  (.Q(\PID_CONTROLLER.err_prev[19] ), 
           .C(clk32MHz), .D(n18490));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i19  (.Q(\PID_CONTROLLER.err_prev[18] ), 
           .C(clk32MHz), .D(n18489));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i18  (.Q(\PID_CONTROLLER.err_prev[17] ), 
           .C(clk32MHz), .D(n18488));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i17  (.Q(\PID_CONTROLLER.err_prev[16] ), 
           .C(clk32MHz), .D(n18487));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i16  (.Q(\PID_CONTROLLER.err_prev[15] ), 
           .C(clk32MHz), .D(n18486));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i15  (.Q(\PID_CONTROLLER.err_prev[14] ), 
           .C(clk32MHz), .D(n18485));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i14  (.Q(\PID_CONTROLLER.err_prev[13] ), 
           .C(clk32MHz), .D(n18484));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i13  (.Q(\PID_CONTROLLER.err_prev[12] ), 
           .C(clk32MHz), .D(n18483));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i12  (.Q(\PID_CONTROLLER.err_prev[11] ), 
           .C(clk32MHz), .D(n18482));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i11  (.Q(\PID_CONTROLLER.err_prev[10] ), 
           .C(clk32MHz), .D(n18481));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i10  (.Q(\PID_CONTROLLER.err_prev[9] ), 
           .C(clk32MHz), .D(n18480));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i9  (.Q(\PID_CONTROLLER.err_prev[8] ), 
           .C(clk32MHz), .D(n18479));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i8  (.Q(\PID_CONTROLLER.err_prev[7] ), 
           .C(clk32MHz), .D(n18478));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i7  (.Q(\PID_CONTROLLER.err_prev[6] ), 
           .C(clk32MHz), .D(n18477));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i6  (.Q(\PID_CONTROLLER.err_prev[5] ), 
           .C(clk32MHz), .D(n18476));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1216_7 (.CI(n36846), .I0(n1802[4]), .I1(n454), 
            .CO(n36847));
    SB_DFF \PID_CONTROLLER.err_prev__i5  (.Q(\PID_CONTROLLER.err_prev[4] ), 
           .C(clk32MHz), .D(n18475));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i4  (.Q(\PID_CONTROLLER.err_prev[3] ), 
           .C(clk32MHz), .D(n18474));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i3  (.Q(\PID_CONTROLLER.err_prev[2] ), 
           .C(clk32MHz), .D(n18473));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i2  (.Q(\PID_CONTROLLER.err_prev[1] ), 
           .C(clk32MHz), .D(n18472));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_4428_5_lut (.I0(GND_net), .I1(n8367[2]), .I2(n404), .I3(n35786), 
            .O(n8339[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_11_lut (.I0(GND_net), .I1(n9591[8]), .I2(GND_net), 
            .I3(n36211), .O(n9555[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_5 (.CI(n35786), .I0(n8367[2]), .I1(n404), .CO(n35787));
    SB_LUT4 add_4428_4_lut (.I0(GND_net), .I1(n8367[1]), .I2(n307_adj_3507), 
            .I3(n35785), .O(n8339[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_11 (.CI(n36211), .I0(n9591[8]), .I1(GND_net), .CO(n36212));
    SB_LUT4 add_4767_10_lut (.I0(GND_net), .I1(n9591[7]), .I2(GND_net), 
            .I3(n36210), .O(n9555[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n57[3]), 
            .I3(n34651), .O(pwm_23__N_3310[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_6_lut (.I0(GND_net), .I1(n9738[3]), .I2(n399), .I3(n36717), 
            .O(n9722[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i30_3_lut (.I0(n12), .I1(\PID_CONTROLLER.result[17] ), 
            .I2(n35_c), .I3(GND_net), .O(n30_adj_3508));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i176_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n261));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i241_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n358));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40031_4_lut (.I0(n13), .I1(n11_adj_3500), .I2(n9), .I3(n47161), 
            .O(n47934));
    defparam i40031_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40027_4_lut (.I0(n19_adj_3499), .I1(n17_adj_3498), .I2(n15_adj_3502), 
            .I3(n47934), .O(n47930));
    defparam i40027_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40892_4_lut (.I0(n25_adj_3493), .I1(n23_adj_3492), .I2(n21), 
            .I3(n47930), .O(n48795));
    defparam i40892_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n455_adj_3509));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4460_11 (.CI(n36513), .I0(n9047[8]), .I1(GND_net), .CO(n36514));
    SB_LUT4 i40380_4_lut (.I0(n31_adj_3496), .I1(n29_adj_3494), .I2(n27), 
            .I3(n48795), .O(n48283));
    defparam i40380_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i41011_4_lut (.I0(n37_adj_3491), .I1(n35_c), .I2(n33_adj_3497), 
            .I3(n48283), .O(n48914));
    defparam i41011_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_4767_10 (.CI(n36210), .I0(n9591[7]), .I1(GND_net), .CO(n36211));
    SB_CARRY add_4428_4 (.CI(n35785), .I0(n8367[1]), .I1(n307_adj_3507), 
            .CO(n35786));
    SB_LUT4 add_4428_3_lut (.I0(GND_net), .I1(n8367[0]), .I2(n210), .I3(n35784), 
            .O(n8339[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40516_3_lut (.I0(n6), .I1(\PID_CONTROLLER.result[10] ), .I2(n21), 
            .I3(GND_net), .O(n48419));   // verilog/motorControl.v(45[12:27])
    defparam i40516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4767_9_lut (.I0(GND_net), .I1(n9591[6]), .I2(GND_net), 
            .I3(n36209), .O(n9555[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n552));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40517_3_lut (.I0(n48419), .I1(\PID_CONTROLLER.result [11]), 
            .I2(n23_adj_3492), .I3(GND_net), .O(n48420));   // verilog/motorControl.v(45[12:27])
    defparam i40517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i24_3_lut (.I0(n16_adj_3510), .I1(\PID_CONTROLLER.result [22]), 
            .I2(n45_adj_3489), .I3(GND_net), .O(n24_adj_3511));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39221_4_lut (.I0(n43_adj_3490), .I1(n25_adj_3493), .I2(n23_adj_3492), 
            .I3(n47150), .O(n47123));
    defparam i39221_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40567_4_lut (.I0(n24_adj_3511), .I1(n8_adj_3512), .I2(n45_adj_3489), 
            .I3(n47121), .O(n48470));   // verilog/motorControl.v(45[12:27])
    defparam i40567_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39811_3_lut (.I0(n48420), .I1(\PID_CONTROLLER.result [12]), 
            .I2(n25_adj_3493), .I3(GND_net), .O(n47714));   // verilog/motorControl.v(45[12:27])
    defparam i39811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i4_4_lut (.I0(\PID_CONTROLLER.result [0]), .I1(\PID_CONTROLLER.result [1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[3]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i436_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n649));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40514_3_lut (.I0(n4), .I1(\PID_CONTROLLER.result[13] ), .I2(n27), 
            .I3(GND_net), .O(n48417));   // verilog/motorControl.v(45[12:27])
    defparam i40514_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4428_3 (.CI(n35784), .I0(n8367[0]), .I1(n210), .CO(n35785));
    SB_LUT4 i40515_3_lut (.I0(n48417), .I1(\PID_CONTROLLER.result [14]), 
            .I2(n29_adj_3494), .I3(GND_net), .O(n48418));   // verilog/motorControl.v(45[12:27])
    defparam i40515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i501_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39238_4_lut (.I0(n33_adj_3497), .I1(n31_adj_3496), .I2(n29_adj_3494), 
            .I3(n47144), .O(n47140));
    defparam i39238_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40950_4_lut (.I0(n30_adj_3508), .I1(n10_adj_3514), .I2(n35_c), 
            .I3(n47138), .O(n48853));   // verilog/motorControl.v(45[12:27])
    defparam i40950_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39813_3_lut (.I0(n48418), .I1(\PID_CONTROLLER.result [15]), 
            .I2(n31_adj_3496), .I3(GND_net), .O(n47716));   // verilog/motorControl.v(45[12:27])
    defparam i39813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41107_4_lut (.I0(n47716), .I1(n48853), .I2(n35_c), .I3(n47140), 
            .O(n49010));   // verilog/motorControl.v(45[12:27])
    defparam i41107_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41108_3_lut (.I0(n49010), .I1(\PID_CONTROLLER.result [18]), 
            .I2(n37_adj_3491), .I3(GND_net), .O(n49011));   // verilog/motorControl.v(45[12:27])
    defparam i41108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41065_3_lut (.I0(n49011), .I1(\PID_CONTROLLER.result[19] ), 
            .I2(n39_c), .I3(GND_net), .O(n48968));   // verilog/motorControl.v(45[12:27])
    defparam i41065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39223_4_lut (.I0(n43_adj_3490), .I1(n41_adj_3488), .I2(n39_c), 
            .I3(n48914), .O(n47125));
    defparam i39223_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40831_4_lut (.I0(n47714), .I1(n48470), .I2(n45_adj_3489), 
            .I3(n47123), .O(n48734));   // verilog/motorControl.v(45[12:27])
    defparam i40831_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39819_3_lut (.I0(n48968), .I1(\PID_CONTROLLER.result [20]), 
            .I2(n41_adj_3488), .I3(GND_net), .O(n47722));   // verilog/motorControl.v(45[12:27])
    defparam i39819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i113_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n167));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40996_4_lut (.I0(n47722), .I1(n48734), .I2(n45_adj_3489), 
            .I3(n47125), .O(n48899));   // verilog/motorControl.v(45[12:27])
    defparam i40996_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i178_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n264));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40997_3_lut (.I0(n48899), .I1(\PID_CONTROLLER.result [23]), 
            .I2(PWMLimit[23]), .I3(GND_net), .O(n48));   // verilog/motorControl.v(45[12:27])
    defparam i40997_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut (.I0(\PID_CONTROLLER.result [26]), .I1(n48), .I2(\PID_CONTROLLER.result [24]), 
            .I3(\PID_CONTROLLER.result [25]), .O(n43052));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_838 (.I0(\PID_CONTROLLER.result [26]), .I1(n48), 
            .I2(\PID_CONTROLLER.result [24]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n43059));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_838.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut (.I0(\PID_CONTROLLER.result [27]), .I1(PWMLimit[23]), 
            .I2(n43059), .I3(n43052), .O(n56));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut.LUT_INIT = 16'hb3a2;
    SB_LUT4 mult_10_i243_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n361));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i23_2_lut  (.I0(deadband[11]), 
            .I1(\PID_CONTROLLER.result [11]), .I2(GND_net), .I3(GND_net), 
            .O(n23_adj_3515));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i23_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i25_2_lut  (.I0(deadband[12]), 
            .I1(\PID_CONTROLLER.result [12]), .I2(GND_net), .I3(GND_net), 
            .O(n25_adj_3516));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i25_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_839 (.I0(\PID_CONTROLLER.result [30]), .I1(n56), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n43083));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_839.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_840 (.I0(\PID_CONTROLLER.result [30]), .I1(n56), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n43089));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_840.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_841 (.I0(PWMLimit[23]), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n43089), .I3(n43083), .O(n387));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_841.LUT_INIT = 16'hb3a2;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[4]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40096_3_lut (.I0(n25_adj_3516), .I1(n23_adj_3515), .I2(n21_adj_1), 
            .I3(GND_net), .O(n47999));
    defparam i40096_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i40068_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\PID_CONTROLLER.result [27]), .I3(n47999), .O(n47971));
    defparam i40068_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n458_adj_3519));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4428_2_lut (.I0(GND_net), .I1(n20_adj_3520), .I2(n113), 
            .I3(GND_net), .O(n8339[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4428_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4428_2 (.CI(GND_net), .I0(n20_adj_3520), .I1(n113), .CO(n35784));
    SB_LUT4 mult_12_i85_2_lut (.I0(\Kd[1] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_3521));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i85_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4783_6 (.CI(n36717), .I0(n9738[3]), .I1(n399), .CO(n36718));
    SB_LUT4 i39369_4_lut (.I0(n21_adj_1), .I1(n19_adj_3487), .I2(n17_adj_3486), 
            .I3(n9_adj_2), .O(n47272));
    defparam i39369_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39347_4_lut (.I0(n43), .I1(n25_adj_3516), .I2(n23_adj_3515), 
            .I3(n47272), .O(n47250));
    defparam i39347_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_12_i22_2_lut (.I0(\Kd[0] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_3523));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40410_4_lut (.I0(deadband[23]), .I1(n45), .I2(\PID_CONTROLLER.result [23]), 
            .I3(n47250), .O(n48313));
    defparam i40410_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n555));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i438_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n652));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40898_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\PID_CONTROLLER.result [25]), .I3(n48313), .O(n48801));
    defparam i40898_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i40070_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\PID_CONTROLLER.result [27]), .I3(n48801), .O(n47973));
    defparam i40070_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[5]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4783_5_lut (.I0(GND_net), .I1(n9738[2]), .I2(n326), .I3(n36716), 
            .O(n9722[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39306_4_lut (.I0(\PID_CONTROLLER.result [15]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(pwm_23__N_3310[15]), .I3(pwm_23__N_3310[14]), .O(n47209));
    defparam i39306_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i40050_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n47209), 
            .I2(pwm_23__N_3310[16]), .I3(GND_net), .O(n47953));
    defparam i40050_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 pwm_23__I_833_i45_rep_313_2_lut (.I0(\PID_CONTROLLER.result [22]), 
            .I1(pwm_23__N_3310[22]), .I2(GND_net), .I3(GND_net), .O(n50655));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i45_rep_313_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[6]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i150_2_lut (.I0(\Kd[2] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n222_adj_3526));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_833_i28_3_lut (.I0(pwm_23__N_3310[14]), .I1(pwm_23__N_3310[15]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(GND_net), .O(n28_adj_3527));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39312_4_lut (.I0(\PID_CONTROLLER.result [12]), .I1(\PID_CONTROLLER.result [11]), 
            .I2(pwm_23__N_3310[12]), .I3(pwm_23__N_3310[11]), .O(n47215));
    defparam i39312_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i40054_3_lut (.I0(pwm_23__N_3310[13]), .I1(n47215), .I2(\PID_CONTROLLER.result[13] ), 
            .I3(GND_net), .O(n47957));
    defparam i40054_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 pwm_23__I_833_i29_rep_308_2_lut (.I0(\PID_CONTROLLER.result [14]), 
            .I1(pwm_23__N_3310[14]), .I2(GND_net), .I3(GND_net), .O(n50650));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i29_rep_308_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40052_4_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n50650), 
            .I2(pwm_23__N_3310[15]), .I3(n47957), .O(n47955));
    defparam i40052_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_4460_10_lut (.I0(GND_net), .I1(n9047[7]), .I2(GND_net), 
            .I3(n36512), .O(n9027[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i49_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n72));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i49_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 pwm_23__I_833_i33_rep_270_2_lut (.I0(\PID_CONTROLLER.result [16]), 
            .I1(pwm_23__N_3310[16]), .I2(GND_net), .I3(GND_net), .O(n50612));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i33_rep_270_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39304_4_lut (.I0(pwm_23__N_3310[17]), .I1(n50612), .I2(\PID_CONTROLLER.result[17] ), 
            .I3(n47955), .O(n47207));
    defparam i39304_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 pwm_23__I_833_i37_rep_282_2_lut (.I0(\PID_CONTROLLER.result [18]), 
            .I1(pwm_23__N_3310[18]), .I2(GND_net), .I3(GND_net), .O(n50624));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i37_rep_282_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40394_4_lut (.I0(pwm_23__N_3310[19]), .I1(n50624), .I2(\PID_CONTROLLER.result[19] ), 
            .I3(n47207), .O(n48297));
    defparam i40394_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 pwm_23__I_833_i41_rep_274_2_lut (.I0(\PID_CONTROLLER.result [20]), 
            .I1(pwm_23__N_3310[20]), .I2(GND_net), .I3(GND_net), .O(n50616));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i41_rep_274_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40894_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(n50616), 
            .I2(pwm_23__N_3310[21]), .I3(n48297), .O(n48797));
    defparam i40894_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i503_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39363_4_lut (.I0(n27_adj_3), .I1(n15_adj_3479), .I2(n13_adj_4), 
            .I3(n11_adj_3467), .O(n47266));
    defparam i39363_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_12_i215_2_lut (.I0(\Kd[3] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n319_adj_3530));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i98_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n145));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i98_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i30_3_lut  (.I0(n12_adj_3531), 
            .I1(\PID_CONTROLLER.result[17] ), .I2(n35), .I3(GND_net), 
            .O(n30_adj_3533));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3534));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4767_9 (.CI(n36209), .I0(n9591[6]), .I1(GND_net), .CO(n36210));
    SB_LUT4 i40108_4_lut (.I0(n9_adj_2), .I1(n7), .I2(deadband[2]), .I3(\PID_CONTROLLER.result [2]), 
            .O(n48011));
    defparam i40108_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i40426_4_lut (.I0(n15_adj_3479), .I1(n13_adj_4), .I2(n11_adj_3467), 
            .I3(n48011), .O(n48329));
    defparam i40426_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i40424_4_lut (.I0(n21_adj_1), .I1(n19_adj_3487), .I2(n17_adj_3486), 
            .I3(n48329), .O(n48327));
    defparam i40424_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[7]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39365_4_lut (.I0(n27_adj_3), .I1(n25_adj_3516), .I2(n23_adj_3515), 
            .I3(n48327), .O(n47268));
    defparam i39365_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_12_i280_2_lut (.I0(\Kd[4] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n416_adj_3536));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40697_4_lut (.I0(n33), .I1(n31), .I2(n29_c), .I3(n47268), 
            .O(n48600));
    defparam i40697_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i41091_4_lut (.I0(n39), .I1(n37), .I2(n35), .I3(n48600), 
            .O(n48994));
    defparam i41091_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i40080_4_lut (.I0(n45), .I1(n43), .I2(n41), .I3(n48994), 
            .O(n47983));
    defparam i40080_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i40693_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [23]), 
            .I2(\PID_CONTROLLER.result [24]), .I3(n47983), .O(n48596));
    defparam i40693_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i41015_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [25]), 
            .I2(\PID_CONTROLLER.result [26]), .I3(n48596), .O(n48918));
    defparam i41015_4_lut.LUT_INIT = 16'hff7e;
    SB_CARRY add_4460_10 (.CI(n36512), .I0(n9047[7]), .I1(GND_net), .CO(n36513));
    SB_LUT4 i41133_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\PID_CONTROLLER.result [28]), .I3(n48918), .O(n49036));
    defparam i41133_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 add_4460_9_lut (.I0(GND_net), .I1(n9047[6]), .I2(GND_net), 
            .I3(n36511), .O(n9027[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40524_3_lut (.I0(n6_adj_3538), .I1(\PID_CONTROLLER.result [26]), 
            .I2(deadband[23]), .I3(GND_net), .O(n48427));   // verilog/motorControl.v(44[10:27])
    defparam i40524_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40062_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(n25_adj_3516), .O(n47965));
    defparam i40062_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i54_4_lut  (.I0(\PID_CONTROLLER.result [12]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(deadband[23]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n54));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i54_4_lut .LUT_INIT = 16'h8f0e;
    SB_CARRY unary_minus_17_add_3_5 (.CI(n34651), .I0(GND_net), .I1(n57[3]), 
            .CO(n34652));
    SB_LUT4 i39330_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n47971), .O(n47233));
    defparam i39330_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i61_rep_266_2_lut  (.I0(deadband[23]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(GND_net), .I3(GND_net), 
            .O(n50608));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i61_rep_266_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 i40562_3_lut (.I0(n54), .I1(n18_adj_3539), .I2(n47965), .I3(GND_net), 
            .O(n48465));   // verilog/motorControl.v(44[10:27])
    defparam i40562_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39801_4_lut (.I0(n48427), .I1(\PID_CONTROLLER.result [28]), 
            .I2(deadband[23]), .I3(\PID_CONTROLLER.result [27]), .O(n47704));   // verilog/motorControl.v(44[10:27])
    defparam i39801_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i24_3_lut  (.I0(n16_adj_3540), 
            .I1(\PID_CONTROLLER.result [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_3541));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i40946_4_lut (.I0(n24_adj_3541), .I1(n8_adj_3542), .I2(n45), 
            .I3(n47248), .O(n48849));   // verilog/motorControl.v(44[10:27])
    defparam i40946_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i40947_3_lut (.I0(n48849), .I1(\PID_CONTROLLER.result [23]), 
            .I2(deadband[23]), .I3(GND_net), .O(n48850));   // verilog/motorControl.v(44[10:27])
    defparam i40947_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40689_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n47973), .O(n48592));
    defparam i40689_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i40990_4_lut (.I0(n47704), .I1(n48465), .I2(n50608), .I3(n47233), 
            .O(n48893));   // verilog/motorControl.v(44[10:27])
    defparam i40990_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39799_4_lut (.I0(n48850), .I1(\PID_CONTROLLER.result [25]), 
            .I2(deadband[23]), .I3(\PID_CONTROLLER.result [24]), .O(n47702));   // verilog/motorControl.v(44[10:27])
    defparam i39799_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 pwm_23__I_833_i26_3_lut (.I0(pwm_23__N_3310[13]), .I1(pwm_23__N_3310[17]), 
            .I2(\PID_CONTROLLER.result[17] ), .I3(GND_net), .O(n26_adj_3543));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39302_4_lut (.I0(pwm_23__N_3310[17]), .I1(pwm_23__N_3310[13]), 
            .I2(\PID_CONTROLLER.result[17] ), .I3(\PID_CONTROLLER.result[13] ), 
            .O(n47205));
    defparam i39302_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_4460_9 (.CI(n36511), .I0(n9047[6]), .I1(GND_net), .CO(n36512));
    SB_LUT4 add_4460_8_lut (.I0(GND_net), .I1(n9047[5]), .I2(n719), .I3(n36510), 
            .O(n9027[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_8_lut (.I0(GND_net), .I1(n9591[5]), .I2(n545), .I3(n36208), 
            .O(n9555[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4427_28_lut (.I0(GND_net), .I1(n8339[25]), .I2(GND_net), 
            .I3(n35783), .O(n8310[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4427_27_lut (.I0(GND_net), .I1(n8339[24]), .I2(GND_net), 
            .I3(n35782), .O(n8310[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_8 (.CI(n36208), .I0(n9591[5]), .I1(n545), .CO(n36209));
    SB_LUT4 add_4767_7_lut (.I0(GND_net), .I1(n9591[4]), .I2(n472), .I3(n36207), 
            .O(n9555[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i345_2_lut (.I0(\Kd[5] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n513_adj_3544));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i345_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4427_27 (.CI(n35782), .I0(n8339[24]), .I1(GND_net), .CO(n35783));
    SB_LUT4 add_4427_26_lut (.I0(GND_net), .I1(n8339[23]), .I2(GND_net), 
            .I3(n35781), .O(n8310[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n57[2]), 
            .I3(n34650), .O(pwm_23__N_3310[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_7 (.CI(n36937), .I0(n9555[4]), .I1(n472), .CO(n36938));
    SB_CARRY add_4427_26 (.CI(n35781), .I0(n8339[23]), .I1(GND_net), .CO(n35782));
    SB_LUT4 mult_14_add_1216_6_lut (.I0(GND_net), .I1(n1802[3]), .I2(n381), 
            .I3(n36845), .O(n1801[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_23__I_833_i24_3_lut (.I0(pwm_23__N_3310[11]), .I1(pwm_23__N_3310[12]), 
            .I2(\PID_CONTROLLER.result [12]), .I3(GND_net), .O(n24_adj_3547));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4427_25_lut (.I0(GND_net), .I1(n8339[22]), .I2(GND_net), 
            .I3(n35780), .O(n8310[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4460_8 (.CI(n36510), .I0(n9047[5]), .I1(n719), .CO(n36511));
    SB_CARRY add_4767_7 (.CI(n36207), .I0(n9591[4]), .I1(n472), .CO(n36208));
    SB_CARRY add_4427_25 (.CI(n35780), .I0(n8339[22]), .I1(GND_net), .CO(n35781));
    SB_LUT4 add_4427_24_lut (.I0(GND_net), .I1(n8339[21]), .I2(GND_net), 
            .I3(n35779), .O(n8310[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_6_lut (.I0(GND_net), .I1(n9591[3]), .I2(n399), .I3(n36206), 
            .O(n9555[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_24 (.CI(n35779), .I0(n8339[21]), .I1(GND_net), .CO(n35780));
    SB_LUT4 add_4427_23_lut (.I0(GND_net), .I1(n8339[20]), .I2(GND_net), 
            .I3(n35778), .O(n8310[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4783_5 (.CI(n36716), .I0(n9738[2]), .I1(n326), .CO(n36717));
    SB_LUT4 add_4460_7_lut (.I0(GND_net), .I1(n9047[4]), .I2(n622), .I3(n36509), 
            .O(n9027[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_6 (.CI(n36206), .I0(n9591[3]), .I1(n399), .CO(n36207));
    SB_CARRY add_4427_23 (.CI(n35778), .I0(n8339[20]), .I1(GND_net), .CO(n35779));
    SB_LUT4 add_4427_22_lut (.I0(GND_net), .I1(n8339[19]), .I2(GND_net), 
            .I3(n35777), .O(n8310[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_5_lut (.I0(GND_net), .I1(n9591[2]), .I2(n326), .I3(n36205), 
            .O(n9555[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_22 (.CI(n35777), .I0(n8339[19]), .I1(GND_net), .CO(n35778));
    SB_LUT4 add_4427_21_lut (.I0(GND_net), .I1(n8339[18]), .I2(GND_net), 
            .I3(n35776), .O(n8310[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4460_7 (.CI(n36509), .I0(n9047[4]), .I1(n622), .CO(n36510));
    SB_CARRY add_4767_5 (.CI(n36205), .I0(n9591[2]), .I1(n326), .CO(n36206));
    SB_CARRY add_4427_21 (.CI(n35776), .I0(n8339[18]), .I1(GND_net), .CO(n35777));
    SB_LUT4 add_4427_20_lut (.I0(GND_net), .I1(n8339[17]), .I2(GND_net), 
            .I3(n35775), .O(n8310[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_4_lut (.I0(GND_net), .I1(n9591[1]), .I2(n253), .I3(n36204), 
            .O(n9555[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_20 (.CI(n35775), .I0(n8339[17]), .I1(GND_net), .CO(n35776));
    SB_LUT4 add_4427_19_lut (.I0(GND_net), .I1(n8339[16]), .I2(GND_net), 
            .I3(n35774), .O(n8310[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i147_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n218_adj_3548));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i147_2_lut.LUT_INIT = 16'h4444;
    SB_DFF \PID_CONTROLLER.result_i0  (.Q(\PID_CONTROLLER.result [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1216_6 (.CI(n36845), .I0(n1802[3]), .I1(n381), 
            .CO(n36846));
    SB_LUT4 add_4783_4_lut (.I0(GND_net), .I1(n9738[1]), .I2(n253), .I3(n36715), 
            .O(n9722[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_6_lut (.I0(GND_net), .I1(n9047[3]), .I2(n525), .I3(n36508), 
            .O(n9027[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_4 (.CI(n36204), .I0(n9591[1]), .I1(n253), .CO(n36205));
    SB_CARRY add_4427_19 (.CI(n35774), .I0(n8339[16]), .I1(GND_net), .CO(n35775));
    SB_LUT4 add_4427_18_lut (.I0(GND_net), .I1(n8339[15]), .I2(GND_net), 
            .I3(n35773), .O(n8310[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_3_lut (.I0(GND_net), .I1(n9591[0]), .I2(n180_adj_3549), 
            .I3(n36203), .O(n9555[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_18 (.CI(n35773), .I0(n8339[15]), .I1(GND_net), .CO(n35774));
    SB_CARRY add_4783_4 (.CI(n36715), .I0(n9738[1]), .I1(n253), .CO(n36716));
    SB_LUT4 mult_10_i505_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_833_i34_3_lut (.I0(n26_adj_3543), .I1(pwm_23__N_3310[18]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(GND_net), .O(n34));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4427_17_lut (.I0(GND_net), .I1(n8339[14]), .I2(GND_net), 
            .I3(n35772), .O(n8310[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40948_4_lut (.I0(n34), .I1(n24_adj_3547), .I2(n50624), .I3(n47205), 
            .O(n48851));   // verilog/motorControl.v(44[31:51])
    defparam i40948_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4427_17 (.CI(n35772), .I0(n8339[14]), .I1(GND_net), .CO(n35773));
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err[0] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4460_6 (.CI(n36508), .I0(n9047[3]), .I1(n525), .CO(n36509));
    SB_LUT4 add_4427_16_lut (.I0(GND_net), .I1(n8339[13]), .I2(GND_net), 
            .I3(n35771), .O(n8310[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF GATES_i2 (.Q(PIN_7_c_1), .C(clk32MHz), .D(GATES_5__N_3138[1]));   // verilog/motorControl.v(64[10] 111[6])
    SB_CARRY add_4767_3 (.CI(n36203), .I0(n9591[0]), .I1(n180_adj_3549), 
            .CO(n36204));
    SB_LUT4 add_4460_5_lut (.I0(GND_net), .I1(n9047[2]), .I2(n428), .I3(n36507), 
            .O(n9027[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4767_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9555[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4767_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_16 (.CI(n35771), .I0(n8339[13]), .I1(GND_net), .CO(n35772));
    SB_LUT4 add_4427_15_lut (.I0(GND_net), .I1(n8339[12]), .I2(GND_net), 
            .I3(n35770), .O(n8310[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_15 (.CI(n35770), .I0(n8339[12]), .I1(GND_net), .CO(n35771));
    SB_LUT4 add_4427_14_lut (.I0(GND_net), .I1(n8339[11]), .I2(GND_net), 
            .I3(n35769), .O(n8310[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4767_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36203));
    SB_CARRY add_4427_14 (.CI(n35769), .I0(n8339[11]), .I1(GND_net), .CO(n35770));
    SB_LUT4 i40949_3_lut (.I0(n48851), .I1(pwm_23__N_3310[19]), .I2(\PID_CONTROLLER.result[19] ), 
            .I3(GND_net), .O(n48852));   // verilog/motorControl.v(44[31:51])
    defparam i40949_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i69_2_lut (.I0(\Kd[1] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i40808_3_lut (.I0(n48852), .I1(pwm_23__N_3310[20]), .I2(\PID_CONTROLLER.result [20]), 
            .I3(GND_net), .O(n48711));   // verilog/motorControl.v(44[31:51])
    defparam i40808_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_17_add_3_4 (.CI(n34650), .I0(GND_net), .I1(n57[2]), 
            .CO(n34651));
    SB_LUT4 add_4427_13_lut (.I0(GND_net), .I1(n8339[10]), .I2(GND_net), 
            .I3(n35768), .O(n8310[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4783_3_lut (.I0(GND_net), .I1(n9738[0]), .I2(n180_adj_3549), 
            .I3(n36714), .O(n9722[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4460_5 (.CI(n36507), .I0(n9047[2]), .I1(n428), .CO(n36508));
    SB_LUT4 add_4770_20_lut (.I0(GND_net), .I1(n9624[17]), .I2(GND_net), 
            .I3(n36202), .O(n9591[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_13 (.CI(n35768), .I0(n8339[10]), .I1(GND_net), .CO(n35769));
    SB_LUT4 add_4770_19_lut (.I0(GND_net), .I1(n9624[16]), .I2(GND_net), 
            .I3(n36201), .O(n9591[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4427_12_lut (.I0(GND_net), .I1(n8339[9]), .I2(GND_net), 
            .I3(n35767), .O(n8310[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i6_2_lut (.I0(\Kd[0] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3551));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4427_12 (.CI(n35767), .I0(n8339[9]), .I1(GND_net), .CO(n35768));
    SB_DFF GATES_i1 (.Q(PIN_6_c_0), .C(clk32MHz), .D(GATES_5__N_3138[0]));   // verilog/motorControl.v(64[10] 111[6])
    SB_CARRY add_4770_19 (.CI(n36201), .I0(n9624[16]), .I1(GND_net), .CO(n36202));
    SB_LUT4 i40518_3_lut (.I0(n22), .I1(pwm_23__N_3310[22]), .I2(\PID_CONTROLLER.result [22]), 
            .I3(GND_net), .O(n48421));   // verilog/motorControl.v(44[31:51])
    defparam i40518_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40519_3_lut (.I0(n48421), .I1(pwm_23__N_3310[23]), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n48422));   // verilog/motorControl.v(44[31:51])
    defparam i40519_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4460_4_lut (.I0(GND_net), .I1(n9047[1]), .I2(n331), .I3(n36506), 
            .O(n9027[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_18_lut (.I0(GND_net), .I1(n9624[15]), .I2(GND_net), 
            .I3(n36200), .O(n9591[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4427_11_lut (.I0(GND_net), .I1(n8339[8]), .I2(GND_net), 
            .I3(n35766), .O(n8310[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4770_18 (.CI(n36200), .I0(n9624[15]), .I1(GND_net), .CO(n36201));
    SB_CARRY add_4427_11 (.CI(n35766), .I0(n8339[8]), .I1(GND_net), .CO(n35767));
    SB_LUT4 add_4427_10_lut (.I0(GND_net), .I1(n8339[7]), .I2(GND_net), 
            .I3(n35765), .O(n8310[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_6_lut (.I0(GND_net), .I1(n9555[3]), .I2(n399), .I3(n36936), 
            .O(n9225[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_5_lut (.I0(GND_net), .I1(n1802[2]), .I2(n308_adj_3555), 
            .I3(n36844), .O(n1801[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4783_3 (.CI(n36714), .I0(n9738[0]), .I1(n180_adj_3549), 
            .CO(n36715));
    SB_CARRY add_4460_4 (.CI(n36506), .I0(n9047[1]), .I1(n331), .CO(n36507));
    SB_LUT4 add_4770_17_lut (.I0(GND_net), .I1(n9624[14]), .I2(GND_net), 
            .I3(n36199), .O(n9591[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_10 (.CI(n35765), .I0(n8339[7]), .I1(GND_net), .CO(n35766));
    SB_LUT4 add_4427_9_lut (.I0(GND_net), .I1(n8339[6]), .I2(GND_net), 
            .I3(n35764), .O(n8310[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4770_17 (.CI(n36199), .I0(n9624[14]), .I1(GND_net), .CO(n36200));
    SB_CARRY add_4427_9 (.CI(n35764), .I0(n8339[6]), .I1(GND_net), .CO(n35765));
    SB_LUT4 add_4427_8_lut (.I0(GND_net), .I1(n8339[5]), .I2(n692), .I3(n35763), 
            .O(n8310[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_3_lut (.I0(GND_net), .I1(n9047[0]), .I2(n234_adj_3556), 
            .I3(n36505), .O(n9027[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_16_lut (.I0(GND_net), .I1(n9624[13]), .I2(GND_net), 
            .I3(n36198), .O(n9591[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_8 (.CI(n35763), .I0(n8339[5]), .I1(n692), .CO(n35764));
    SB_LUT4 add_4427_7_lut (.I0(GND_net), .I1(n8339[4]), .I2(n595), .I3(n35762), 
            .O(n8310[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4770_16 (.CI(n36198), .I0(n9624[13]), .I1(GND_net), .CO(n36199));
    SB_CARRY add_4427_7 (.CI(n35762), .I0(n8339[4]), .I1(n595), .CO(n35763));
    SB_LUT4 add_4427_6_lut (.I0(GND_net), .I1(n8339[3]), .I2(n498), .I3(n35761), 
            .O(n8310[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i410_2_lut (.I0(\Kd[6] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n610_adj_3557));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4783_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9722[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4783_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4460_3 (.CI(n36505), .I0(n9047[0]), .I1(n234_adj_3556), 
            .CO(n36506));
    SB_LUT4 add_4770_15_lut (.I0(GND_net), .I1(n9624[12]), .I2(GND_net), 
            .I3(n36197), .O(n9591[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40037_4_lut (.I0(\PID_CONTROLLER.result [23]), .I1(n50655), 
            .I2(pwm_23__N_3310[23]), .I3(n47953), .O(n47940));
    defparam i40037_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_4427_6 (.CI(n35761), .I0(n8339[3]), .I1(n498), .CO(n35762));
    SB_LUT4 add_4427_5_lut (.I0(GND_net), .I1(n8339[2]), .I2(n401_c), 
            .I3(n35760), .O(n8310[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_23__I_833_i30_3_lut (.I0(n28_adj_3527), .I1(pwm_23__N_3310[16]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(GND_net), .O(n30_adj_3558));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i134_2_lut (.I0(\Kd[2] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4770_15 (.CI(n36197), .I0(n9624[12]), .I1(GND_net), .CO(n36198));
    SB_CARRY add_4427_5 (.CI(n35760), .I0(n8339[2]), .I1(n401_c), .CO(n35761));
    SB_LUT4 add_4427_4_lut (.I0(GND_net), .I1(n8339[1]), .I2(n304), .I3(n35759), 
            .O(n8310[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4460_2_lut (.I0(GND_net), .I1(n44), .I2(n137), .I3(GND_net), 
            .O(n9027[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4460_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_14_lut (.I0(GND_net), .I1(n9624[11]), .I2(GND_net), 
            .I3(n36196), .O(n9591[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4427_4 (.CI(n35759), .I0(n8339[1]), .I1(n304), .CO(n35760));
    SB_LUT4 add_4427_3_lut (.I0(GND_net), .I1(n8339[0]), .I2(n207), .I3(n35758), 
            .O(n8310[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39809_3_lut (.I0(n48422), .I1(pwm_23__N_3310[24]), .I2(n43813), 
            .I3(GND_net), .O(n47712));   // verilog/motorControl.v(44[31:51])
    defparam i39809_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4473_6 (.CI(n36936), .I0(n9555[3]), .I1(n399), .CO(n36937));
    SB_LUT4 i40040_4_lut (.I0(\PID_CONTROLLER.result [23]), .I1(n50655), 
            .I2(pwm_23__N_3310[23]), .I3(n48797), .O(n47943));
    defparam i40040_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_4427_3 (.CI(n35758), .I0(n8339[0]), .I1(n207), .CO(n35759));
    SB_LUT4 add_4427_2_lut (.I0(GND_net), .I1(n17_adj_3559), .I2(n110), 
            .I3(GND_net), .O(n8310[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4427_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4770_14 (.CI(n36196), .I0(n9624[11]), .I1(GND_net), .CO(n36197));
    SB_CARRY add_4427_2 (.CI(GND_net), .I0(n17_adj_3559), .I1(n110), .CO(n35758));
    SB_LUT4 i40398_4_lut (.I0(n47712), .I1(n30_adj_3558), .I2(n43813), 
            .I3(n47940), .O(n48301));   // verilog/motorControl.v(44[31:51])
    defparam i40398_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4426_29_lut (.I0(GND_net), .I1(n8310[26]), .I2(GND_net), 
            .I3(n35757), .O(n8280[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39807_3_lut (.I0(n48711), .I1(pwm_23__N_3310[21]), .I2(\PID_CONTROLLER.result [21]), 
            .I3(GND_net), .O(n47710));   // verilog/motorControl.v(44[31:51])
    defparam i39807_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40566_4_lut (.I0(n47710), .I1(n48301), .I2(n43813), .I3(n47943), 
            .O(n48469));   // verilog/motorControl.v(44[31:51])
    defparam i40566_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4770_13_lut (.I0(GND_net), .I1(n9624[10]), .I2(GND_net), 
            .I3(n36195), .O(n9591[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i4_4_lut  (.I0(deadband[0]), .I1(\PID_CONTROLLER.result [1]), 
            .I2(deadband[1]), .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3560));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i4_4_lut .LUT_INIT = 16'h4d0c;
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n57[1]), 
            .I3(n34649), .O(pwm_23__N_3310[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40534_3_lut (.I0(n4_adj_3560), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(n27_adj_3), .I3(GND_net), .O(n48437));   // verilog/motorControl.v(44[10:27])
    defparam i40534_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_17_add_3_3 (.CI(n34649), .I0(GND_net), .I1(n57[1]), 
            .CO(n34650));
    SB_CARRY add_4460_2 (.CI(GND_net), .I0(n44), .I1(n137), .CO(n36505));
    SB_CARRY add_4770_13 (.CI(n36195), .I0(n9624[10]), .I1(GND_net), .CO(n36196));
    SB_CARRY mult_14_add_1216_5 (.CI(n36844), .I0(n1802[2]), .I1(n308_adj_3555), 
            .CO(n36845));
    SB_CARRY add_4783_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36714));
    SB_LUT4 add_4459_20_lut (.I0(GND_net), .I1(n9027[17]), .I2(GND_net), 
            .I3(n36504), .O(n9006[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_12_lut (.I0(GND_net), .I1(n9624[9]), .I2(GND_net), 
            .I3(n36194), .O(n9591[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40535_3_lut (.I0(n48437), .I1(\PID_CONTROLLER.result [14]), 
            .I2(n29_c), .I3(GND_net), .O(n48438));   // verilog/motorControl.v(44[10:27])
    defparam i40535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4426_28_lut (.I0(GND_net), .I1(n8310[25]), .I2(GND_net), 
            .I3(n35756), .O(n8280[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_28 (.CI(n35756), .I0(n8310[25]), .I1(GND_net), .CO(n35757));
    SB_CARRY add_4770_12 (.CI(n36194), .I0(n9624[9]), .I1(GND_net), .CO(n36195));
    SB_LUT4 add_4426_27_lut (.I0(GND_net), .I1(n8310[24]), .I2(GND_net), 
            .I3(n35755), .O(n8280[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_27 (.CI(n35755), .I0(n8310[24]), .I1(GND_net), .CO(n35756));
    SB_LUT4 add_4459_19_lut (.I0(GND_net), .I1(n9027[16]), .I2(GND_net), 
            .I3(n36503), .O(n9006[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_11_lut (.I0(GND_net), .I1(n9624[8]), .I2(GND_net), 
            .I3(n36193), .O(n9591[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_26_lut (.I0(GND_net), .I1(n8310[23]), .I2(GND_net), 
            .I3(n35754), .O(n8280[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_26 (.CI(n35754), .I0(n8310[23]), .I1(GND_net), .CO(n35755));
    SB_CARRY add_4770_11 (.CI(n36193), .I0(n9624[8]), .I1(GND_net), .CO(n36194));
    SB_LUT4 add_4426_25_lut (.I0(GND_net), .I1(n8310[22]), .I2(GND_net), 
            .I3(n35753), .O(n8280[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_25 (.CI(n35753), .I0(n8310[22]), .I1(GND_net), .CO(n35754));
    SB_LUT4 mult_14_i196_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i196_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_4784_14_lut (.I0(GND_net), .I1(n9753[11]), .I2(GND_net), 
            .I3(n36713), .O(n9738[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_19 (.CI(n36503), .I0(n9027[16]), .I1(GND_net), .CO(n36504));
    SB_LUT4 add_4770_10_lut (.I0(GND_net), .I1(n9624[7]), .I2(GND_net), 
            .I3(n36192), .O(n9591[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_24_lut (.I0(GND_net), .I1(n8310[21]), .I2(GND_net), 
            .I3(n35752), .O(n8280[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_24 (.CI(n35752), .I0(n8310[21]), .I1(GND_net), .CO(n35753));
    SB_CARRY add_4770_10 (.CI(n36192), .I0(n9624[7]), .I1(GND_net), .CO(n36193));
    SB_LUT4 add_4426_23_lut (.I0(GND_net), .I1(n8310[20]), .I2(GND_net), 
            .I3(n35751), .O(n8280[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_23 (.CI(n35751), .I0(n8310[20]), .I1(GND_net), .CO(n35752));
    SB_LUT4 i39359_4_lut (.I0(n33), .I1(n31), .I2(n29_c), .I3(n47266), 
            .O(n47262));
    defparam i39359_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4459_18_lut (.I0(GND_net), .I1(n9027[15]), .I2(GND_net), 
            .I3(n36502), .O(n9006[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_9_lut (.I0(GND_net), .I1(n9624[6]), .I2(GND_net), 
            .I3(n36191), .O(n9591[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_22_lut (.I0(GND_net), .I1(n8310[19]), .I2(GND_net), 
            .I3(n35750), .O(n8280[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_22 (.CI(n35750), .I0(n8310[19]), .I1(GND_net), .CO(n35751));
    SB_LUT4 mult_12_i475_2_lut (.I0(\Kd[7] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n707_adj_3562));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i475_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4770_9 (.CI(n36191), .I0(n9624[6]), .I1(GND_net), .CO(n36192));
    SB_LUT4 add_4426_21_lut (.I0(GND_net), .I1(n8310[18]), .I2(GND_net), 
            .I3(n35749), .O(n8280[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_21 (.CI(n35749), .I0(n8310[18]), .I1(GND_net), .CO(n35750));
    SB_LUT4 i40944_4_lut (.I0(n30_adj_3533), .I1(n10_adj_3563), .I2(n35), 
            .I3(n47260), .O(n48847));   // verilog/motorControl.v(44[10:27])
    defparam i40944_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4473_5_lut (.I0(GND_net), .I1(n9555[2]), .I2(n326), .I3(n36935), 
            .O(n9225[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i199_2_lut (.I0(\Kd[3] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n295));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1216_4_lut (.I0(GND_net), .I1(n1802[1]), .I2(n235_adj_3565), 
            .I3(n36843), .O(n1801[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_13_lut (.I0(GND_net), .I1(n9753[10]), .I2(GND_net), 
            .I3(n36712), .O(n9738[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_18 (.CI(n36502), .I0(n9027[15]), .I1(GND_net), .CO(n36503));
    SB_LUT4 add_4770_8_lut (.I0(GND_net), .I1(n9624[5]), .I2(n545), .I3(n36190), 
            .O(n9591[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_20_lut (.I0(GND_net), .I1(n8310[17]), .I2(GND_net), 
            .I3(n35748), .O(n8280[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_20 (.CI(n35748), .I0(n8310[17]), .I1(GND_net), .CO(n35749));
    SB_CARRY add_4770_8 (.CI(n36190), .I0(n9624[5]), .I1(n545), .CO(n36191));
    SB_LUT4 add_4426_19_lut (.I0(GND_net), .I1(n8310[16]), .I2(GND_net), 
            .I3(n35747), .O(n8280[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_19 (.CI(n35747), .I0(n8310[16]), .I1(GND_net), .CO(n35748));
    SB_LUT4 add_4459_17_lut (.I0(GND_net), .I1(n9027[14]), .I2(GND_net), 
            .I3(n36501), .O(n9006[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_7_lut (.I0(GND_net), .I1(n9624[4]), .I2(n472), .I3(n36189), 
            .O(n9591[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_18_lut (.I0(GND_net), .I1(n8310[15]), .I2(GND_net), 
            .I3(n35746), .O(n8280[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_18 (.CI(n35746), .I0(n8310[15]), .I1(GND_net), .CO(n35747));
    SB_CARRY add_4770_7 (.CI(n36189), .I0(n9624[4]), .I1(n472), .CO(n36190));
    SB_LUT4 add_4426_17_lut (.I0(GND_net), .I1(n8310[14]), .I2(GND_net), 
            .I3(n35745), .O(n8280[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_17 (.CI(n35745), .I0(n8310[14]), .I1(GND_net), .CO(n35746));
    SB_CARRY add_4784_13 (.CI(n36712), .I0(n9753[10]), .I1(GND_net), .CO(n36713));
    SB_CARRY add_4459_17 (.CI(n36501), .I0(n9027[14]), .I1(GND_net), .CO(n36502));
    SB_LUT4 add_4770_6_lut (.I0(GND_net), .I1(n9624[3]), .I2(n399), .I3(n36188), 
            .O(n9591[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_16_lut (.I0(GND_net), .I1(n8310[13]), .I2(GND_net), 
            .I3(n35744), .O(n8280[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_16 (.CI(n35744), .I0(n8310[13]), .I1(GND_net), .CO(n35745));
    SB_CARRY add_4770_6 (.CI(n36188), .I0(n9624[3]), .I1(n399), .CO(n36189));
    SB_LUT4 add_4426_15_lut (.I0(GND_net), .I1(n8310[12]), .I2(GND_net), 
            .I3(n35743), .O(n8280[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_15 (.CI(n35743), .I0(n8310[12]), .I1(GND_net), .CO(n35744));
    SB_LUT4 add_4459_16_lut (.I0(GND_net), .I1(n9027[13]), .I2(GND_net), 
            .I3(n36500), .O(n9006[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[8]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4770_5_lut (.I0(GND_net), .I1(n9624[2]), .I2(n326), .I3(n36187), 
            .O(n9591[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_14_lut (.I0(GND_net), .I1(n8310[11]), .I2(GND_net), 
            .I3(n35742), .O(n8280[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_14 (.CI(n35742), .I0(n8310[11]), .I1(GND_net), .CO(n35743));
    SB_CARRY add_4770_5 (.CI(n36187), .I0(n9624[2]), .I1(n326), .CO(n36188));
    SB_LUT4 add_4426_13_lut (.I0(GND_net), .I1(n8310[10]), .I2(GND_net), 
            .I3(n35741), .O(n8280[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_13 (.CI(n35741), .I0(n8310[10]), .I1(GND_net), .CO(n35742));
    SB_CARRY mult_14_add_1216_4 (.CI(n36843), .I0(n1802[1]), .I1(n235_adj_3565), 
            .CO(n36844));
    SB_LUT4 add_4784_12_lut (.I0(GND_net), .I1(n9753[9]), .I2(GND_net), 
            .I3(n36711), .O(n9738[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_16 (.CI(n36500), .I0(n9027[13]), .I1(GND_net), .CO(n36501));
    SB_LUT4 add_4770_4_lut (.I0(GND_net), .I1(n9624[1]), .I2(n253), .I3(n36186), 
            .O(n9591[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_12_lut (.I0(GND_net), .I1(n8310[9]), .I2(GND_net), 
            .I3(n35740), .O(n8280[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_12 (.CI(n35740), .I0(n8310[9]), .I1(GND_net), .CO(n35741));
    SB_CARRY add_4770_4 (.CI(n36186), .I0(n9624[1]), .I1(n253), .CO(n36187));
    SB_LUT4 add_4426_11_lut (.I0(GND_net), .I1(n8310[8]), .I2(GND_net), 
            .I3(n35739), .O(n8280[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_11 (.CI(n35739), .I0(n8310[8]), .I1(GND_net), .CO(n35740));
    SB_LUT4 add_4459_15_lut (.I0(GND_net), .I1(n9027[12]), .I2(GND_net), 
            .I3(n36499), .O(n9006[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4770_3_lut (.I0(GND_net), .I1(n9624[0]), .I2(n180_adj_3549), 
            .I3(n36185), .O(n9591[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_10_lut (.I0(GND_net), .I1(n8310[7]), .I2(GND_net), 
            .I3(n35738), .O(n8280[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_10 (.CI(n35738), .I0(n8310[7]), .I1(GND_net), .CO(n35739));
    SB_CARRY add_4770_3 (.CI(n36185), .I0(n9624[0]), .I1(n180_adj_3549), 
            .CO(n36186));
    SB_LUT4 add_4426_9_lut (.I0(GND_net), .I1(n8310[6]), .I2(GND_net), 
            .I3(n35737), .O(n8280[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_9 (.CI(n35737), .I0(n8310[6]), .I1(GND_net), .CO(n35738));
    SB_CARRY add_4784_12 (.CI(n36711), .I0(n9753[9]), .I1(GND_net), .CO(n36712));
    SB_CARRY add_4459_15 (.CI(n36499), .I0(n9027[12]), .I1(GND_net), .CO(n36500));
    SB_LUT4 add_4770_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9591[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4770_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_8_lut (.I0(GND_net), .I1(n8310[5]), .I2(n689), .I3(n35736), 
            .O(n8280[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4770_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36185));
    SB_CARRY add_4426_8 (.CI(n35736), .I0(n8310[5]), .I1(n689), .CO(n35737));
    SB_LUT4 add_4426_7_lut (.I0(GND_net), .I1(n8310[4]), .I2(n592), .I3(n35735), 
            .O(n8280[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4459_14_lut (.I0(GND_net), .I1(n9027[11]), .I2(GND_net), 
            .I3(n36498), .O(n9006[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_19_lut (.I0(GND_net), .I1(n9654[16]), .I2(GND_net), 
            .I3(n36184), .O(n9624[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_7 (.CI(n35735), .I0(n8310[4]), .I1(n592), .CO(n35736));
    SB_LUT4 add_4773_18_lut (.I0(GND_net), .I1(n9654[15]), .I2(GND_net), 
            .I3(n36183), .O(n9624[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_6_lut (.I0(GND_net), .I1(n8310[3]), .I2(n495), .I3(n35734), 
            .O(n8280[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_6 (.CI(n35734), .I0(n8310[3]), .I1(n495), .CO(n35735));
    SB_LUT4 i39789_3_lut (.I0(n48438), .I1(\PID_CONTROLLER.result [15]), 
            .I2(n31), .I3(GND_net), .O(n47692));   // verilog/motorControl.v(44[10:27])
    defparam i39789_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4473_5 (.CI(n36935), .I0(n9555[2]), .I1(n326), .CO(n36936));
    SB_LUT4 add_4426_5_lut (.I0(GND_net), .I1(n8310[2]), .I2(n398), .I3(n35733), 
            .O(n8280[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_3_lut (.I0(GND_net), .I1(n1802[0]), .I2(n162), 
            .I3(n36842), .O(n1801[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_11_lut (.I0(GND_net), .I1(n9753[8]), .I2(GND_net), 
            .I3(n36710), .O(n9738[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_14 (.CI(n36498), .I0(n9027[11]), .I1(GND_net), .CO(n36499));
    SB_CARRY add_4773_18 (.CI(n36183), .I0(n9654[15]), .I1(GND_net), .CO(n36184));
    SB_CARRY add_4426_5 (.CI(n35733), .I0(n8310[2]), .I1(n398), .CO(n35734));
    SB_LUT4 add_4426_4_lut (.I0(GND_net), .I1(n8310[1]), .I2(n301), .I3(n35732), 
            .O(n8280[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_4 (.CI(n35732), .I0(n8310[1]), .I1(n301), .CO(n35733));
    SB_LUT4 mult_12_i264_2_lut (.I0(\Kd[4] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n392));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4773_17_lut (.I0(GND_net), .I1(n9654[14]), .I2(GND_net), 
            .I3(n36182), .O(n9624[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_3_lut (.I0(GND_net), .I1(n8310[0]), .I2(n204), .I3(n35731), 
            .O(n8280[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_3 (.CI(n35731), .I0(n8310[0]), .I1(n204), .CO(n35732));
    SB_LUT4 add_4459_13_lut (.I0(GND_net), .I1(n9027[10]), .I2(GND_net), 
            .I3(n36497), .O(n9006[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_17 (.CI(n36182), .I0(n9654[14]), .I1(GND_net), .CO(n36183));
    SB_LUT4 add_4773_16_lut (.I0(GND_net), .I1(n9654[13]), .I2(GND_net), 
            .I3(n36181), .O(n9624[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_2_lut (.I0(GND_net), .I1(n14), .I2(n107_adj_3567), 
            .I3(GND_net), .O(n8280[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_2 (.CI(GND_net), .I0(n14), .I1(n107_adj_3567), .CO(n35731));
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n25957), .I1(GND_net), .I2(n57[0]), 
            .I3(VCC_net), .O(n46520)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n57[0]), 
            .CO(n34649));
    SB_CARRY add_4784_11 (.CI(n36710), .I0(n9753[8]), .I1(GND_net), .CO(n36711));
    SB_CARRY add_4459_13 (.CI(n36497), .I0(n9027[10]), .I1(GND_net), .CO(n36498));
    SB_LUT4 add_4473_4_lut (.I0(GND_net), .I1(n9555[1]), .I2(n253), .I3(n36934), 
            .O(n9225[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_10_lut (.I0(GND_net), .I1(n9753[7]), .I2(GND_net), 
            .I3(n36709), .O(n9738[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4459_12_lut (.I0(GND_net), .I1(n9027[9]), .I2(GND_net), 
            .I3(n36496), .O(n9006[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_10 (.CI(n36709), .I0(n9753[7]), .I1(GND_net), .CO(n36710));
    SB_LUT4 add_4425_30_lut (.I0(GND_net), .I1(n8280[27]), .I2(GND_net), 
            .I3(n35730), .O(n8249[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_16 (.CI(n36181), .I0(n9654[13]), .I1(GND_net), .CO(n36182));
    SB_CARRY add_4459_12 (.CI(n36496), .I0(n9027[9]), .I1(GND_net), .CO(n36497));
    SB_LUT4 add_4773_15_lut (.I0(GND_net), .I1(n9654[12]), .I2(GND_net), 
            .I3(n36180), .O(n9624[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_15 (.CI(n36180), .I0(n9654[12]), .I1(GND_net), .CO(n36181));
    SB_LUT4 unary_minus_70_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(GATES_5__N_3405), 
            .I3(n34765), .O(n853)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_4 (.CI(n36934), .I0(n9555[1]), .I1(n253), .CO(n36935));
    SB_LUT4 add_4425_29_lut (.I0(GND_net), .I1(n8280[26]), .I2(GND_net), 
            .I3(n35729), .O(n8249[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_29 (.CI(n35729), .I0(n8280[26]), .I1(GND_net), .CO(n35730));
    SB_LUT4 add_4773_14_lut (.I0(GND_net), .I1(n9654[11]), .I2(GND_net), 
            .I3(n36179), .O(n9624[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_24_lut (.I0(n852[18]), .I1(GND_net), .I2(n63[22]), 
            .I3(n34764), .O(n44276)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_70_add_3_24 (.CI(n34764), .I0(GND_net), .I1(n63[22]), 
            .CO(n34765));
    SB_CARRY mult_14_add_1216_3 (.CI(n36842), .I0(n1802[0]), .I1(n162), 
            .CO(n36843));
    SB_LUT4 i41105_4_lut (.I0(n47692), .I1(n48847), .I2(n35), .I3(n47262), 
            .O(n49008));   // verilog/motorControl.v(44[10:27])
    defparam i41105_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41106_3_lut (.I0(n49008), .I1(\PID_CONTROLLER.result [18]), 
            .I2(n37), .I3(GND_net), .O(n49009));   // verilog/motorControl.v(44[10:27])
    defparam i41106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i329_2_lut (.I0(\Kd[5] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n489));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i329_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4773_14 (.CI(n36179), .I0(n9654[11]), .I1(GND_net), .CO(n36180));
    SB_LUT4 unary_minus_70_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n63[21]), 
            .I3(n34763), .O(n855)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_28_lut (.I0(GND_net), .I1(n8280[25]), .I2(GND_net), 
            .I3(n35728), .O(n8249[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_28 (.CI(n35728), .I0(n8280[25]), .I1(GND_net), .CO(n35729));
    SB_LUT4 i41069_3_lut (.I0(n49009), .I1(\PID_CONTROLLER.result[19] ), 
            .I2(n39), .I3(GND_net), .O(n48972));   // verilog/motorControl.v(44[10:27])
    defparam i41069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41169_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(n49036), .O(n49072));
    defparam i41169_4_lut.LUT_INIT = 16'hff7e;
    SB_CARRY unary_minus_70_add_3_23 (.CI(n34763), .I0(GND_net), .I1(n63[21]), 
            .CO(n34764));
    SB_LUT4 add_4473_3_lut (.I0(GND_net), .I1(n9555[0]), .I2(n180_adj_3549), 
            .I3(n36933), .O(n9225[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n63[20]), 
            .I3(n34762), .O(n856)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_9_lut (.I0(GND_net), .I1(n9753[6]), .I2(GND_net), 
            .I3(n36708), .O(n9738[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_27_lut (.I0(GND_net), .I1(n8280[24]), .I2(GND_net), 
            .I3(n35727), .O(n8249[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40992_4_lut (.I0(n47702), .I1(n48893), .I2(n50608), .I3(n48592), 
            .O(n48895));   // verilog/motorControl.v(44[10:27])
    defparam i40992_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4459_11_lut (.I0(GND_net), .I1(n9027[8]), .I2(GND_net), 
            .I3(n36495), .O(n9006[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_13_lut (.I0(GND_net), .I1(n9654[10]), .I2(GND_net), 
            .I3(n36178), .O(n9624[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_2_lut (.I0(GND_net), .I1(n20_adj_3571), .I2(n89), 
            .I3(GND_net), .O(n1801[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_22 (.CI(n34762), .I0(GND_net), .I1(n63[20]), 
            .CO(n34763));
    SB_LUT4 i39795_3_lut (.I0(n48972), .I1(\PID_CONTROLLER.result [20]), 
            .I2(n41), .I3(GND_net), .O(n47698));   // verilog/motorControl.v(44[10:27])
    defparam i39795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_833_i64_3_lut (.I0(n48469), .I1(\PID_CONTROLLER.result [31]), 
            .I2(pwm_23__N_3310[24]), .I3(GND_net), .O(pwm_23__N_3309));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i64_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4459_11 (.CI(n36495), .I0(n9027[8]), .I1(GND_net), .CO(n36496));
    SB_CARRY add_4773_13 (.CI(n36178), .I0(n9654[10]), .I1(GND_net), .CO(n36179));
    SB_LUT4 add_4773_12_lut (.I0(GND_net), .I1(n9654[9]), .I2(GND_net), 
            .I3(n36177), .O(n9624[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_27 (.CI(n35727), .I0(n8280[24]), .I1(GND_net), .CO(n35728));
    SB_LUT4 add_4425_26_lut (.I0(GND_net), .I1(n8280[23]), .I2(GND_net), 
            .I3(n35726), .O(n8249[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_9 (.CI(n36708), .I0(n9753[6]), .I1(GND_net), .CO(n36709));
    SB_CARRY mult_14_add_1216_2 (.CI(GND_net), .I0(n20_adj_3571), .I1(n89), 
            .CO(n36842));
    SB_LUT4 i40994_3_lut (.I0(n47698), .I1(n48895), .I2(n49072), .I3(GND_net), 
            .O(n48897));   // verilog/motorControl.v(44[10:27])
    defparam i40994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i245_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n364));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i245_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_4459_10_lut (.I0(GND_net), .I1(n9027[7]), .I2(GND_net), 
            .I3(n36494), .O(n9006[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_8_lut (.I0(GND_net), .I1(n9753[5]), .I2(n545), .I3(n36707), 
            .O(n9738[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_12 (.CI(n36177), .I0(n9654[9]), .I1(GND_net), .CO(n36178));
    SB_CARRY add_4459_10 (.CI(n36494), .I0(n9027[7]), .I1(GND_net), .CO(n36495));
    SB_CARRY add_4425_26 (.CI(n35726), .I0(n8280[23]), .I1(GND_net), .CO(n35727));
    SB_LUT4 add_4459_9_lut (.I0(GND_net), .I1(n9027[6]), .I2(GND_net), 
            .I3(n36493), .O(n9006[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[9]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4425_25_lut (.I0(GND_net), .I1(n8280[22]), .I2(GND_net), 
            .I3(n35725), .O(n8249[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n63[19]), 
            .I3(n34761), .O(n857)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_9 (.CI(n36493), .I0(n9027[6]), .I1(GND_net), .CO(n36494));
    SB_LUT4 add_4459_8_lut (.I0(GND_net), .I1(n9027[5]), .I2(n716), .I3(n36492), 
            .O(n9006[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_25 (.CI(n35725), .I0(n8280[22]), .I1(GND_net), .CO(n35726));
    SB_LUT4 add_4425_24_lut (.I0(GND_net), .I1(n8280[21]), .I2(GND_net), 
            .I3(n35724), .O(n8249[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_11_lut (.I0(GND_net), .I1(n9654[8]), .I2(GND_net), 
            .I3(n36176), .O(n9624[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_24 (.CI(n35724), .I0(n8280[21]), .I1(GND_net), .CO(n35725));
    SB_LUT4 pwm_23__I_832_4_lut (.I0(n48897), .I1(pwm_23__N_3309), .I2(deadband[23]), 
            .I3(\PID_CONTROLLER.result [31]), .O(pwm_23__N_3307));   // verilog/motorControl.v(44[10:51])
    defparam pwm_23__I_832_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 add_4425_23_lut (.I0(GND_net), .I1(n8280[20]), .I2(GND_net), 
            .I3(n35723), .O(n8249[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_8 (.CI(n36707), .I0(n9753[5]), .I1(n545), .CO(n36708));
    SB_CARRY add_4773_11 (.CI(n36176), .I0(n9654[8]), .I1(GND_net), .CO(n36177));
    SB_CARRY add_4425_23 (.CI(n35723), .I0(n8280[20]), .I1(GND_net), .CO(n35724));
    SB_CARRY unary_minus_70_add_3_21 (.CI(n34761), .I0(GND_net), .I1(n63[19]), 
            .CO(n34762));
    SB_LUT4 unary_minus_70_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n63[18]), 
            .I3(n34760), .O(n852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_8 (.CI(n36492), .I0(n9027[5]), .I1(n716), .CO(n36493));
    SB_LUT4 add_4784_7_lut (.I0(GND_net), .I1(n9753[4]), .I2(n472), .I3(n36706), 
            .O(n9738[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4459_7_lut (.I0(GND_net), .I1(n9027[4]), .I2(n619), .I3(n36491), 
            .O(n9006[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_10_lut (.I0(GND_net), .I1(n9654[7]), .I2(GND_net), 
            .I3(n36175), .O(n9624[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_20 (.CI(n34760), .I0(GND_net), .I1(n63[18]), 
            .CO(n34761));
    SB_LUT4 add_4425_22_lut (.I0(GND_net), .I1(n8280[19]), .I2(GND_net), 
            .I3(n35722), .O(n8249[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_22 (.CI(n35722), .I0(n8280[19]), .I1(GND_net), .CO(n35723));
    SB_LUT4 unary_minus_70_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n63[17]), 
            .I3(n34759), .O(n859)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_7 (.CI(n36491), .I0(n9027[4]), .I1(n619), .CO(n36492));
    SB_CARRY unary_minus_70_add_3_19 (.CI(n34759), .I0(GND_net), .I1(n63[17]), 
            .CO(n34760));
    SB_CARRY add_4773_10 (.CI(n36175), .I0(n9654[7]), .I1(GND_net), .CO(n36176));
    SB_LUT4 add_4773_9_lut (.I0(GND_net), .I1(n9654[6]), .I2(GND_net), 
            .I3(n36174), .O(n9624[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_9 (.CI(n36174), .I0(n9654[6]), .I1(GND_net), .CO(n36175));
    SB_CARRY add_4473_3 (.CI(n36933), .I0(n9555[0]), .I1(n180_adj_3549), 
            .CO(n36934));
    SB_LUT4 unary_minus_70_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n63[16]), 
            .I3(n34758), .O(n860)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_8_lut (.I0(GND_net), .I1(n9654[5]), .I2(n545), .I3(n36173), 
            .O(n9624[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_24_lut (.I0(GND_net), .I1(n1801[21]), .I2(GND_net), 
            .I3(n36840), .O(n1800[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_7 (.CI(n36706), .I0(n9753[4]), .I1(n472), .CO(n36707));
    SB_LUT4 add_4459_6_lut (.I0(GND_net), .I1(n9027[3]), .I2(n522), .I3(n36490), 
            .O(n9006[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_21_lut (.I0(GND_net), .I1(n8280[18]), .I2(GND_net), 
            .I3(n35721), .O(n8249[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_21 (.CI(n35721), .I0(n8280[18]), .I1(GND_net), .CO(n35722));
    SB_CARRY add_4773_8 (.CI(n36173), .I0(n9654[5]), .I1(n545), .CO(n36174));
    SB_LUT4 add_4425_20_lut (.I0(GND_net), .I1(n8280[17]), .I2(GND_net), 
            .I3(n35720), .O(n8249[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_20 (.CI(n35720), .I0(n8280[17]), .I1(GND_net), .CO(n35721));
    SB_LUT4 add_4425_19_lut (.I0(GND_net), .I1(n8280[16]), .I2(GND_net), 
            .I3(n35719), .O(n8249[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_19 (.CI(n35719), .I0(n8280[16]), .I1(GND_net), .CO(n35720));
    SB_LUT4 add_4773_7_lut (.I0(GND_net), .I1(n9654[4]), .I2(n472), .I3(n36172), 
            .O(n9624[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_18_lut (.I0(GND_net), .I1(n8280[15]), .I2(GND_net), 
            .I3(n35718), .O(n8249[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_18 (.CI(n35718), .I0(n8280[15]), .I1(GND_net), .CO(n35719));
    SB_CARRY unary_minus_70_add_3_18 (.CI(n34758), .I0(GND_net), .I1(n63[16]), 
            .CO(n34759));
    SB_LUT4 unary_minus_70_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n63[15]), 
            .I3(n34757), .O(n861)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_7 (.CI(n36172), .I0(n9654[4]), .I1(n472), .CO(n36173));
    SB_CARRY unary_minus_70_add_3_17 (.CI(n34757), .I0(GND_net), .I1(n63[15]), 
            .CO(n34758));
    SB_CARRY mult_14_add_1215_24 (.CI(n36840), .I0(n1801[21]), .I1(GND_net), 
            .CO(n1699));
    SB_LUT4 unary_minus_70_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n63[14]), 
            .I3(n34756), .O(n862)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_6 (.CI(n36490), .I0(n9027[3]), .I1(n522), .CO(n36491));
    SB_LUT4 add_4773_6_lut (.I0(GND_net), .I1(n9654[3]), .I2(n399), .I3(n36171), 
            .O(n9624[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4459_5_lut (.I0(GND_net), .I1(n9027[2]), .I2(n425), .I3(n36489), 
            .O(n9006[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_17_lut (.I0(GND_net), .I1(n8280[14]), .I2(GND_net), 
            .I3(n35717), .O(n8249[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_17 (.CI(n35717), .I0(n8280[14]), .I1(GND_net), .CO(n35718));
    SB_CARRY add_4773_6 (.CI(n36171), .I0(n9654[3]), .I1(n399), .CO(n36172));
    SB_LUT4 add_4425_16_lut (.I0(GND_net), .I1(n8280[13]), .I2(GND_net), 
            .I3(n35716), .O(n8249[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_16 (.CI(n35716), .I0(n8280[13]), .I1(GND_net), .CO(n35717));
    SB_CARRY unary_minus_70_add_3_16 (.CI(n34756), .I0(GND_net), .I1(n63[14]), 
            .CO(n34757));
    SB_LUT4 unary_minus_70_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n63[13]), 
            .I3(n34755), .O(n863)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_6_lut (.I0(GND_net), .I1(n9753[3]), .I2(n399), .I3(n36705), 
            .O(n9738[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_5 (.CI(n36489), .I0(n9027[2]), .I1(n425), .CO(n36490));
    SB_LUT4 add_4773_5_lut (.I0(GND_net), .I1(n9654[2]), .I2(n326), .I3(n36170), 
            .O(n9624[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_15_lut (.I0(GND_net), .I1(n8280[12]), .I2(GND_net), 
            .I3(n35715), .O(n8249[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_6 (.CI(n36705), .I0(n9753[3]), .I1(n399), .CO(n36706));
    SB_CARRY add_4425_15 (.CI(n35715), .I0(n8280[12]), .I1(GND_net), .CO(n35716));
    SB_LUT4 add_4459_4_lut (.I0(GND_net), .I1(n9027[1]), .I2(n328), .I3(n36488), 
            .O(n9006[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_15 (.CI(n34755), .I0(GND_net), .I1(n63[13]), 
            .CO(n34756));
    SB_CARRY add_4773_5 (.CI(n36170), .I0(n9654[2]), .I1(n326), .CO(n36171));
    SB_LUT4 add_4425_14_lut (.I0(GND_net), .I1(n8280[11]), .I2(GND_net), 
            .I3(n35714), .O(n8249[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n63[12]), 
            .I3(n34754), .O(n864)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_5_lut (.I0(GND_net), .I1(n9753[2]), .I2(n326), .I3(n36704), 
            .O(n9738[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_4 (.CI(n36488), .I0(n9027[1]), .I1(n328), .CO(n36489));
    SB_LUT4 add_4773_4_lut (.I0(GND_net), .I1(n9654[1]), .I2(n253), .I3(n36169), 
            .O(n9624[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_14 (.CI(n35714), .I0(n8280[11]), .I1(GND_net), .CO(n35715));
    SB_CARRY add_4773_4 (.CI(n36169), .I0(n9654[1]), .I1(n253), .CO(n36170));
    SB_LUT4 add_4773_3_lut (.I0(GND_net), .I1(n9654[0]), .I2(n180_adj_3549), 
            .I3(n36168), .O(n9624[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_5 (.CI(n36704), .I0(n9753[2]), .I1(n326), .CO(n36705));
    SB_LUT4 add_4459_3_lut (.I0(GND_net), .I1(n9027[0]), .I2(n231_adj_3581), 
            .I3(n36487), .O(n9006[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_13_lut (.I0(GND_net), .I1(n8280[10]), .I2(GND_net), 
            .I3(n35713), .O(n8249[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_13 (.CI(n35713), .I0(n8280[10]), .I1(GND_net), .CO(n35714));
    SB_CARRY add_4773_3 (.CI(n36168), .I0(n9654[0]), .I1(n180_adj_3549), 
            .CO(n36169));
    SB_LUT4 add_4773_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9624[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_12_lut (.I0(GND_net), .I1(n8280[9]), .I2(GND_net), 
            .I3(n35712), .O(n8249[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_12 (.CI(n35712), .I0(n8280[9]), .I1(GND_net), .CO(n35713));
    SB_CARRY add_4773_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36168));
    SB_CARRY add_4459_3 (.CI(n36487), .I0(n9027[0]), .I1(n231_adj_3581), 
            .CO(n36488));
    SB_LUT4 add_4784_4_lut (.I0(GND_net), .I1(n9753[1]), .I2(n253), .I3(n36703), 
            .O(n9738[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_11_lut (.I0(GND_net), .I1(n8280[8]), .I2(GND_net), 
            .I3(n35711), .O(n8249[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_11 (.CI(n35711), .I0(n8280[8]), .I1(GND_net), .CO(n35712));
    SB_LUT4 add_4776_18_lut (.I0(GND_net), .I1(n9681[15]), .I2(GND_net), 
            .I3(n36167), .O(n9654[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_10_lut (.I0(GND_net), .I1(n8280[7]), .I2(GND_net), 
            .I3(n35710), .O(n8249[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_10 (.CI(n35710), .I0(n8280[7]), .I1(GND_net), .CO(n35711));
    SB_CARRY unary_minus_70_add_3_14 (.CI(n34754), .I0(GND_net), .I1(n63[12]), 
            .CO(n34755));
    SB_LUT4 unary_minus_70_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n63[11]), 
            .I3(n34753), .O(n865)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_13 (.CI(n34753), .I0(GND_net), .I1(n63[11]), 
            .CO(n34754));
    SB_LUT4 add_4425_9_lut (.I0(GND_net), .I1(n8280[6]), .I2(GND_net), 
            .I3(n35709), .O(n8249[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4459_2_lut (.I0(GND_net), .I1(n41_adj_3583), .I2(n134), 
            .I3(GND_net), .O(n9006[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4459_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_9 (.CI(n35709), .I0(n8280[6]), .I1(GND_net), .CO(n35710));
    SB_CARRY add_4784_4 (.CI(n36703), .I0(n9753[1]), .I1(n253), .CO(n36704));
    SB_LUT4 add_4425_8_lut (.I0(GND_net), .I1(n8280[5]), .I2(n686_adj_3584), 
            .I3(n35708), .O(n8249[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4459_2 (.CI(GND_net), .I0(n41_adj_3583), .I1(n134), .CO(n36487));
    SB_LUT4 add_4458_21_lut (.I0(GND_net), .I1(n9006[18]), .I2(GND_net), 
            .I3(n36486), .O(n8984[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_17_lut (.I0(GND_net), .I1(n9681[14]), .I2(GND_net), 
            .I3(n36166), .O(n9654[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_17 (.CI(n36166), .I0(n9681[14]), .I1(GND_net), .CO(n36167));
    SB_CARRY add_4425_8 (.CI(n35708), .I0(n8280[5]), .I1(n686_adj_3584), 
            .CO(n35709));
    SB_LUT4 add_4425_7_lut (.I0(GND_net), .I1(n8280[4]), .I2(n589_adj_3585), 
            .I3(n35707), .O(n8249[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_20_lut (.I0(GND_net), .I1(n9006[17]), .I2(GND_net), 
            .I3(n36485), .O(n8984[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n63[10]), 
            .I3(n34752), .O(n866)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_16_lut (.I0(GND_net), .I1(n9681[13]), .I2(GND_net), 
            .I3(n36165), .O(n9654[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_16 (.CI(n36165), .I0(n9681[13]), .I1(GND_net), .CO(n36166));
    SB_CARRY unary_minus_70_add_3_12 (.CI(n34752), .I0(GND_net), .I1(n63[10]), 
            .CO(n34753));
    SB_CARRY add_4425_7 (.CI(n35707), .I0(n8280[4]), .I1(n589_adj_3585), 
            .CO(n35708));
    SB_LUT4 add_4473_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9225[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_6_lut (.I0(GND_net), .I1(n8280[3]), .I2(n492_adj_3587), 
            .I3(n35706), .O(n8249[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_6 (.CI(n35706), .I0(n8280[3]), .I1(n492_adj_3587), 
            .CO(n35707));
    SB_LUT4 mult_14_add_1215_23_lut (.I0(GND_net), .I1(n1801[20]), .I2(GND_net), 
            .I3(n36839), .O(n1800[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_5_lut (.I0(GND_net), .I1(n8280[2]), .I2(n395_adj_3588), 
            .I3(n35705), .O(n8249[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_15_lut (.I0(GND_net), .I1(n9681[12]), .I2(GND_net), 
            .I3(n36164), .O(n9654[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_5 (.CI(n35705), .I0(n8280[2]), .I1(n395_adj_3588), 
            .CO(n35706));
    SB_CARRY add_4473_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36933));
    SB_LUT4 add_4784_3_lut (.I0(GND_net), .I1(n9753[0]), .I2(n180_adj_3549), 
            .I3(n36702), .O(n9738[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_20 (.CI(n36485), .I0(n9006[17]), .I1(GND_net), .CO(n36486));
    SB_LUT4 add_4425_4_lut (.I0(GND_net), .I1(n8280[1]), .I2(n298_adj_3589), 
            .I3(n35704), .O(n8249[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_4 (.CI(n35704), .I0(n8280[1]), .I1(n298_adj_3589), 
            .CO(n35705));
    SB_CARRY mult_14_add_1215_23 (.CI(n36839), .I0(n1801[20]), .I1(GND_net), 
            .CO(n36840));
    SB_CARRY add_4784_3 (.CI(n36702), .I0(n9753[0]), .I1(n180_adj_3549), 
            .CO(n36703));
    SB_CARRY add_4776_15 (.CI(n36164), .I0(n9681[12]), .I1(GND_net), .CO(n36165));
    SB_LUT4 add_4776_14_lut (.I0(GND_net), .I1(n9681[11]), .I2(GND_net), 
            .I3(n36163), .O(n9654[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_22_lut (.I0(GND_net), .I1(n1801[19]), .I2(GND_net), 
            .I3(n36838), .O(n1800[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n63[9]), 
            .I3(n34751), .O(n867)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_11 (.CI(n34751), .I0(GND_net), .I1(n63[9]), 
            .CO(n34752));
    SB_CARRY mult_14_add_1215_22 (.CI(n36838), .I0(n1801[19]), .I1(GND_net), 
            .CO(n36839));
    SB_LUT4 mult_14_add_1215_21_lut (.I0(GND_net), .I1(n1801[18]), .I2(GND_net), 
            .I3(n36837), .O(n1800[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4425_3_lut (.I0(GND_net), .I1(n8280[0]), .I2(n201_adj_3591), 
            .I3(n35703), .O(n8249[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_21 (.CI(n36837), .I0(n1801[18]), .I1(GND_net), 
            .CO(n36838));
    SB_LUT4 add_4458_19_lut (.I0(GND_net), .I1(n9006[16]), .I2(GND_net), 
            .I3(n36484), .O(n8984[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_14 (.CI(n36163), .I0(n9681[11]), .I1(GND_net), .CO(n36164));
    SB_CARRY add_4425_3 (.CI(n35703), .I0(n8280[0]), .I1(n201_adj_3591), 
            .CO(n35704));
    SB_LUT4 add_4425_2_lut (.I0(GND_net), .I1(n11_adj_3592), .I2(n104_adj_3593), 
            .I3(GND_net), .O(n8249[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4425_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_13_lut (.I0(GND_net), .I1(n9681[10]), .I2(GND_net), 
            .I3(n36162), .O(n9654[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4784_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9738[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4784_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4425_2 (.CI(GND_net), .I0(n11_adj_3592), .I1(n104_adj_3593), 
            .CO(n35703));
    SB_LUT4 mult_14_add_1219_24_lut (.I0(GND_net), .I1(n9201[21]), .I2(GND_net), 
            .I3(n36932), .O(n1804[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_13 (.CI(n36162), .I0(n9681[10]), .I1(GND_net), .CO(n36163));
    SB_LUT4 mult_14_add_1219_23_lut (.I0(GND_net), .I1(n9201[20]), .I2(GND_net), 
            .I3(n36931), .O(n1804[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_32_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n8217[29]), 
            .I2(GND_net), .I3(n35702), .O(n6807[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_70_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n63[8]), 
            .I3(n34750), .O(n868)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4784_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36702));
    SB_LUT4 mult_14_add_1215_20_lut (.I0(GND_net), .I1(n1801[17]), .I2(GND_net), 
            .I3(n36836), .O(n1800[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_31_lut (.I0(GND_net), .I1(n8217[28]), .I2(GND_net), 
            .I3(n35701), .O(n64[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_10 (.CI(n34750), .I0(GND_net), .I1(n63[8]), 
            .CO(n34751));
    SB_CARRY mult_14_add_1215_20 (.CI(n36836), .I0(n1801[17]), .I1(GND_net), 
            .CO(n36837));
    SB_LUT4 unary_minus_70_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n63[7]), 
            .I3(n34749), .O(n869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_13_lut (.I0(GND_net), .I1(n9767[10]), .I2(GND_net), 
            .I3(n36701), .O(n9753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_19 (.CI(n36484), .I0(n9006[16]), .I1(GND_net), .CO(n36485));
    SB_LUT4 add_4458_18_lut (.I0(GND_net), .I1(n9006[15]), .I2(GND_net), 
            .I3(n36483), .O(n8984[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_12_lut (.I0(GND_net), .I1(n9681[9]), .I2(GND_net), 
            .I3(n36161), .O(n9654[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_31 (.CI(n35701), .I0(n8217[28]), .I1(GND_net), 
            .CO(n35702));
    SB_CARRY unary_minus_70_add_3_9 (.CI(n34749), .I0(GND_net), .I1(n63[7]), 
            .CO(n34750));
    SB_LUT4 add_4785_12_lut (.I0(GND_net), .I1(n9767[9]), .I2(GND_net), 
            .I3(n36700), .O(n9753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_23 (.CI(n36931), .I0(n9201[20]), .I1(GND_net), 
            .CO(n36932));
    SB_LUT4 mult_14_add_1215_19_lut (.I0(GND_net), .I1(n1801[16]), .I2(GND_net), 
            .I3(n36835), .O(n1800[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_19 (.CI(n36835), .I0(n1801[16]), .I1(GND_net), 
            .CO(n36836));
    SB_CARRY add_4785_12 (.CI(n36700), .I0(n9767[9]), .I1(GND_net), .CO(n36701));
    SB_CARRY add_4458_18 (.CI(n36483), .I0(n9006[15]), .I1(GND_net), .CO(n36484));
    SB_LUT4 mult_10_add_2137_30_lut (.I0(GND_net), .I1(n8217[27]), .I2(GND_net), 
            .I3(n35700), .O(n64[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n63[6]), 
            .I3(n34748), .O(n870)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_30 (.CI(n35700), .I0(n8217[27]), .I1(GND_net), 
            .CO(n35701));
    SB_LUT4 mult_14_add_1215_18_lut (.I0(GND_net), .I1(n1801[15]), .I2(GND_net), 
            .I3(n36834), .O(n1800[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_8 (.CI(n34748), .I0(GND_net), .I1(n63[6]), 
            .CO(n34749));
    SB_LUT4 add_4785_11_lut (.I0(GND_net), .I1(n9767[8]), .I2(GND_net), 
            .I3(n36699), .O(n9753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_17_lut (.I0(GND_net), .I1(n9006[14]), .I2(GND_net), 
            .I3(n36482), .O(n8984[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_11 (.CI(n36699), .I0(n9767[8]), .I1(GND_net), .CO(n36700));
    SB_CARRY add_4776_12 (.CI(n36161), .I0(n9681[9]), .I1(GND_net), .CO(n36162));
    SB_LUT4 mult_14_add_1219_22_lut (.I0(GND_net), .I1(n9201[19]), .I2(GND_net), 
            .I3(n36930), .O(n1804[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_18 (.CI(n36834), .I0(n1801[15]), .I1(GND_net), 
            .CO(n36835));
    SB_LUT4 add_4776_11_lut (.I0(GND_net), .I1(n9681[8]), .I2(GND_net), 
            .I3(n36160), .O(n9654[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_22 (.CI(n36930), .I0(n9201[19]), .I1(GND_net), 
            .CO(n36931));
    SB_LUT4 mult_14_add_1215_17_lut (.I0(GND_net), .I1(n1801[14]), .I2(GND_net), 
            .I3(n36833), .O(n1800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_10_lut (.I0(GND_net), .I1(n9767[7]), .I2(GND_net), 
            .I3(n36698), .O(n9753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_10 (.CI(n36698), .I0(n9767[7]), .I1(GND_net), .CO(n36699));
    SB_CARRY add_4458_17 (.CI(n36482), .I0(n9006[14]), .I1(GND_net), .CO(n36483));
    SB_LUT4 mult_10_add_2137_29_lut (.I0(GND_net), .I1(n8217[26]), .I2(GND_net), 
            .I3(n35699), .O(n64[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_21_lut (.I0(GND_net), .I1(n9201[18]), .I2(GND_net), 
            .I3(n36929), .O(n1804[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_9_lut (.I0(GND_net), .I1(n9767[6]), .I2(GND_net), 
            .I3(n36697), .O(n9753[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_21 (.CI(n36929), .I0(n9201[18]), .I1(GND_net), 
            .CO(n36930));
    SB_CARRY mult_14_add_1215_17 (.CI(n36833), .I0(n1801[14]), .I1(GND_net), 
            .CO(n36834));
    SB_CARRY add_4776_11 (.CI(n36160), .I0(n9681[8]), .I1(GND_net), .CO(n36161));
    SB_CARRY mult_10_add_2137_29 (.CI(n35699), .I0(n8217[26]), .I1(GND_net), 
            .CO(n35700));
    SB_CARRY add_4785_9 (.CI(n36697), .I0(n9767[6]), .I1(GND_net), .CO(n36698));
    SB_LUT4 mult_10_add_2137_28_lut (.I0(GND_net), .I1(n8217[25]), .I2(GND_net), 
            .I3(n35698), .O(n64[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_10_lut (.I0(GND_net), .I1(n9681[7]), .I2(GND_net), 
            .I3(n36159), .O(n9654[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_10 (.CI(n36159), .I0(n9681[7]), .I1(GND_net), .CO(n36160));
    SB_LUT4 unary_minus_70_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n63[5]), 
            .I3(n34747), .O(n871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_20_lut (.I0(GND_net), .I1(n9201[17]), .I2(GND_net), 
            .I3(n36928), .O(n1804[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_7 (.CI(n34747), .I0(GND_net), .I1(n63[5]), 
            .CO(n34748));
    SB_LUT4 add_4458_16_lut (.I0(GND_net), .I1(n9006[13]), .I2(GND_net), 
            .I3(n36481), .O(n8984[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_16_lut (.I0(GND_net), .I1(n1801[13]), .I2(GND_net), 
            .I3(n36832), .O(n1800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_16 (.CI(n36832), .I0(n1801[13]), .I1(GND_net), 
            .CO(n36833));
    SB_LUT4 add_4776_9_lut (.I0(GND_net), .I1(n9681[6]), .I2(GND_net), 
            .I3(n36158), .O(n9654[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_28 (.CI(n35698), .I0(n8217[25]), .I1(GND_net), 
            .CO(n35699));
    SB_LUT4 add_4785_8_lut (.I0(GND_net), .I1(n9767[5]), .I2(n545), .I3(n36696), 
            .O(n9753[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_8 (.CI(n36696), .I0(n9767[5]), .I1(n545), .CO(n36697));
    SB_LUT4 unary_minus_70_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n63[4]), 
            .I3(n34746), .O(n872)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_27_lut (.I0(GND_net), .I1(n8217[24]), .I2(GND_net), 
            .I3(n35697), .O(n64[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_15_lut (.I0(GND_net), .I1(n1801[12]), .I2(GND_net), 
            .I3(n36831), .O(n1800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_27 (.CI(n35697), .I0(n8217[24]), .I1(GND_net), 
            .CO(n35698));
    SB_CARRY add_4776_9 (.CI(n36158), .I0(n9681[6]), .I1(GND_net), .CO(n36159));
    SB_LUT4 add_4785_7_lut (.I0(GND_net), .I1(n9767[4]), .I2(n472), .I3(n36695), 
            .O(n9753[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_8_lut (.I0(GND_net), .I1(n9681[5]), .I2(n545), .I3(n36157), 
            .O(n9654[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_26_lut (.I0(GND_net), .I1(n8217[23]), .I2(GND_net), 
            .I3(n35696), .O(n64[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_7 (.CI(n36695), .I0(n9767[4]), .I1(n472), .CO(n36696));
    SB_CARRY mult_10_add_2137_26 (.CI(n35696), .I0(n8217[23]), .I1(GND_net), 
            .CO(n35697));
    SB_LUT4 mult_10_add_2137_25_lut (.I0(GND_net), .I1(n8217[22]), .I2(GND_net), 
            .I3(n35695), .O(n64[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_20 (.CI(n36928), .I0(n9201[17]), .I1(GND_net), 
            .CO(n36929));
    SB_LUT4 mult_14_add_1219_19_lut (.I0(GND_net), .I1(n9201[16]), .I2(GND_net), 
            .I3(n36927), .O(n1804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_25 (.CI(n35695), .I0(n8217[22]), .I1(GND_net), 
            .CO(n35696));
    SB_CARRY add_4776_8 (.CI(n36157), .I0(n9681[5]), .I1(n545), .CO(n36158));
    SB_CARRY add_4458_16 (.CI(n36481), .I0(n9006[13]), .I1(GND_net), .CO(n36482));
    SB_CARRY mult_14_add_1219_19 (.CI(n36927), .I0(n9201[16]), .I1(GND_net), 
            .CO(n36928));
    SB_CARRY mult_14_add_1215_15 (.CI(n36831), .I0(n1801[12]), .I1(GND_net), 
            .CO(n36832));
    SB_LUT4 mult_14_add_1215_14_lut (.I0(GND_net), .I1(n1801[11]), .I2(GND_net), 
            .I3(n36830), .O(n1800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_24_lut (.I0(GND_net), .I1(n8217[21]), .I2(GND_net), 
            .I3(n35694), .O(n64[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_6_lut (.I0(GND_net), .I1(n9767[3]), .I2(n399), .I3(n36694), 
            .O(n9753[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_14 (.CI(n36830), .I0(n1801[11]), .I1(GND_net), 
            .CO(n36831));
    SB_LUT4 mult_14_add_1219_18_lut (.I0(GND_net), .I1(n9201[15]), .I2(GND_net), 
            .I3(n36926), .O(n1804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_13_lut (.I0(GND_net), .I1(n1801[10]), .I2(GND_net), 
            .I3(n36829), .O(n1800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_18 (.CI(n36926), .I0(n9201[15]), .I1(GND_net), 
            .CO(n36927));
    SB_CARRY mult_14_add_1215_13 (.CI(n36829), .I0(n1801[10]), .I1(GND_net), 
            .CO(n36830));
    SB_CARRY add_4785_6 (.CI(n36694), .I0(n9767[3]), .I1(n399), .CO(n36695));
    SB_LUT4 add_4458_15_lut (.I0(GND_net), .I1(n9006[12]), .I2(GND_net), 
            .I3(n36480), .O(n8984[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_17_lut (.I0(GND_net), .I1(n9201[14]), .I2(GND_net), 
            .I3(n36925), .O(n1804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_5_lut (.I0(GND_net), .I1(n9767[2]), .I2(n326), .I3(n36693), 
            .O(n9753[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_7_lut (.I0(GND_net), .I1(n9681[4]), .I2(n472), .I3(n36156), 
            .O(n9654[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_12_lut (.I0(GND_net), .I1(n1801[9]), .I2(GND_net), 
            .I3(n36828), .O(n1800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_5 (.CI(n36693), .I0(n9767[2]), .I1(n326), .CO(n36694));
    SB_LUT4 add_4785_4_lut (.I0(GND_net), .I1(n9767[1]), .I2(n253), .I3(n36692), 
            .O(n9753[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_15 (.CI(n36480), .I0(n9006[12]), .I1(GND_net), .CO(n36481));
    SB_CARRY add_4785_4 (.CI(n36692), .I0(n9767[1]), .I1(n253), .CO(n36693));
    SB_LUT4 add_4458_14_lut (.I0(GND_net), .I1(n9006[11]), .I2(GND_net), 
            .I3(n36479), .O(n8984[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_14 (.CI(n36479), .I0(n9006[11]), .I1(GND_net), .CO(n36480));
    SB_CARRY mult_10_add_2137_24 (.CI(n35694), .I0(n8217[21]), .I1(GND_net), 
            .CO(n35695));
    SB_CARRY add_4776_7 (.CI(n36156), .I0(n9681[4]), .I1(n472), .CO(n36157));
    SB_LUT4 mult_10_add_2137_23_lut (.I0(GND_net), .I1(n8217[20]), .I2(GND_net), 
            .I3(n35693), .O(n64[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_6 (.CI(n34746), .I0(GND_net), .I1(n63[4]), 
            .CO(n34747));
    SB_LUT4 unary_minus_70_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n63[3]), 
            .I3(n34745), .O(n873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_6_lut (.I0(GND_net), .I1(n9681[3]), .I2(n399), .I3(n36155), 
            .O(n9654[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_13_lut (.I0(GND_net), .I1(n9006[10]), .I2(GND_net), 
            .I3(n36478), .O(n8984[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4785_3_lut (.I0(GND_net), .I1(n9767[0]), .I2(n180_adj_3549), 
            .I3(n36691), .O(n9753[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_23 (.CI(n35693), .I0(n8217[20]), .I1(GND_net), 
            .CO(n35694));
    SB_CARRY add_4776_6 (.CI(n36155), .I0(n9681[3]), .I1(n399), .CO(n36156));
    SB_LUT4 add_4776_5_lut (.I0(GND_net), .I1(n9681[2]), .I2(n326), .I3(n36154), 
            .O(n9654[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_22_lut (.I0(GND_net), .I1(n8217[19]), .I2(GND_net), 
            .I3(n35692), .O(n64[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_22 (.CI(n35692), .I0(n8217[19]), .I1(GND_net), 
            .CO(n35693));
    SB_LUT4 mult_10_add_2137_21_lut (.I0(GND_net), .I1(n8217[18]), .I2(GND_net), 
            .I3(n35691), .O(n64[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_13 (.CI(n36478), .I0(n9006[10]), .I1(GND_net), .CO(n36479));
    SB_CARRY mult_10_add_2137_21 (.CI(n35691), .I0(n8217[18]), .I1(GND_net), 
            .CO(n35692));
    SB_CARRY add_4776_5 (.CI(n36154), .I0(n9681[2]), .I1(n326), .CO(n36155));
    SB_LUT4 add_4458_12_lut (.I0(GND_net), .I1(n9006[9]), .I2(GND_net), 
            .I3(n36477), .O(n8984[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_4_lut (.I0(GND_net), .I1(n9681[1]), .I2(n253), .I3(n36153), 
            .O(n9654[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_20_lut (.I0(GND_net), .I1(n8217[17]), .I2(GND_net), 
            .I3(n35690), .O(n64[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_12 (.CI(n36828), .I0(n1801[9]), .I1(GND_net), 
            .CO(n36829));
    SB_CARRY mult_14_add_1219_17 (.CI(n36925), .I0(n9201[14]), .I1(GND_net), 
            .CO(n36926));
    SB_CARRY add_4776_4 (.CI(n36153), .I0(n9681[1]), .I1(n253), .CO(n36154));
    SB_LUT4 add_4776_3_lut (.I0(GND_net), .I1(n9681[0]), .I2(n180_adj_3549), 
            .I3(n36152), .O(n9654[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_11_lut (.I0(GND_net), .I1(n1801[8]), .I2(GND_net), 
            .I3(n36827), .O(n1800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4785_3 (.CI(n36691), .I0(n9767[0]), .I1(n180_adj_3549), 
            .CO(n36692));
    SB_CARRY add_4458_12 (.CI(n36477), .I0(n9006[9]), .I1(GND_net), .CO(n36478));
    SB_LUT4 add_4458_11_lut (.I0(GND_net), .I1(n9006[8]), .I2(GND_net), 
            .I3(n36476), .O(n8984[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_5 (.CI(n34745), .I0(GND_net), .I1(n63[3]), 
            .CO(n34746));
    SB_LUT4 unary_minus_70_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n63[2]), 
            .I3(n34744), .O(n874)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4776_3 (.CI(n36152), .I0(n9681[0]), .I1(n180_adj_3549), 
            .CO(n36153));
    SB_CARRY mult_10_add_2137_20 (.CI(n35690), .I0(n8217[17]), .I1(GND_net), 
            .CO(n35691));
    SB_LUT4 mult_10_add_2137_19_lut (.I0(GND_net), .I1(n8217[16]), .I2(GND_net), 
            .I3(n35689), .O(n64[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4776_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9654[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4776_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_19 (.CI(n35689), .I0(n8217[16]), .I1(GND_net), 
            .CO(n35690));
    SB_CARRY unary_minus_70_add_3_4 (.CI(n34744), .I0(GND_net), .I1(n63[2]), 
            .CO(n34745));
    SB_CARRY mult_14_add_1215_11 (.CI(n36827), .I0(n1801[8]), .I1(GND_net), 
            .CO(n36828));
    SB_LUT4 add_4785_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9753[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4785_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n63[1]), 
            .I3(n34743), .O(n875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_11 (.CI(n36476), .I0(n9006[8]), .I1(GND_net), .CO(n36477));
    SB_CARRY add_4785_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36691));
    SB_CARRY add_4776_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36152));
    SB_LUT4 mult_10_add_2137_18_lut (.I0(GND_net), .I1(n8217[15]), .I2(GND_net), 
            .I3(n35688), .O(n64[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_3 (.CI(n34743), .I0(GND_net), .I1(n63[1]), 
            .CO(n34744));
    SB_CARRY mult_10_add_2137_18 (.CI(n35688), .I0(n8217[15]), .I1(GND_net), 
            .CO(n35689));
    SB_LUT4 add_4458_10_lut (.I0(GND_net), .I1(n9006[7]), .I2(GND_net), 
            .I3(n36475), .O(n8984[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_17_lut (.I0(GND_net), .I1(n8217[14]), .I2(GND_net), 
            .I3(n35687), .O(n64[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_16_lut (.I0(GND_net), .I1(n9201[13]), .I2(GND_net), 
            .I3(n36924), .O(n1804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_17 (.CI(n35687), .I0(n8217[14]), .I1(GND_net), 
            .CO(n35688));
    SB_CARRY add_4458_10 (.CI(n36475), .I0(n9006[7]), .I1(GND_net), .CO(n36476));
    SB_LUT4 add_4458_9_lut (.I0(GND_net), .I1(n9006[6]), .I2(GND_net), 
            .I3(n36474), .O(n8984[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_17_lut (.I0(GND_net), .I1(n9705[14]), .I2(GND_net), 
            .I3(n36151), .O(n9681[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_12_lut (.I0(GND_net), .I1(n9780[9]), .I2(GND_net), 
            .I3(n36690), .O(n9767[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_9 (.CI(n36474), .I0(n9006[6]), .I1(GND_net), .CO(n36475));
    SB_LUT4 mult_10_add_2137_16_lut (.I0(GND_net), .I1(n8217[13]), .I2(GND_net), 
            .I3(n35686), .O(n64[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_16 (.CI(n36924), .I0(n9201[13]), .I1(GND_net), 
            .CO(n36925));
    SB_LUT4 add_4779_16_lut (.I0(GND_net), .I1(n9705[13]), .I2(GND_net), 
            .I3(n36150), .O(n9681[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_10_lut (.I0(GND_net), .I1(n1801[7]), .I2(GND_net), 
            .I3(n36826), .O(n1800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_8_lut (.I0(GND_net), .I1(n9006[5]), .I2(n713), .I3(n36473), 
            .O(n8984[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_2_lut (.I0(n25958), .I1(GND_net), .I2(n63[0]), 
            .I3(VCC_net), .O(n46548)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4779_16 (.CI(n36150), .I0(n9705[13]), .I1(GND_net), .CO(n36151));
    SB_LUT4 mult_14_add_1219_15_lut (.I0(GND_net), .I1(n9201[12]), .I2(GND_net), 
            .I3(n36923), .O(n1804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_15_lut (.I0(GND_net), .I1(n9705[12]), .I2(GND_net), 
            .I3(n36149), .O(n9681[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_10 (.CI(n36826), .I0(n1801[7]), .I1(GND_net), 
            .CO(n36827));
    SB_LUT4 add_4786_11_lut (.I0(GND_net), .I1(n9780[8]), .I2(GND_net), 
            .I3(n36689), .O(n9767[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_8 (.CI(n36473), .I0(n9006[5]), .I1(n713), .CO(n36474));
    SB_CARRY add_4779_15 (.CI(n36149), .I0(n9705[12]), .I1(GND_net), .CO(n36150));
    SB_LUT4 add_4458_7_lut (.I0(GND_net), .I1(n9006[4]), .I2(n616), .I3(n36472), 
            .O(n8984[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_15 (.CI(n36923), .I0(n9201[12]), .I1(GND_net), 
            .CO(n36924));
    SB_LUT4 mult_12_i394_2_lut (.I0(\Kd[6] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n586));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_2137_16 (.CI(n35686), .I0(n8217[13]), .I1(GND_net), 
            .CO(n35687));
    SB_LUT4 mult_10_i127_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n176));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i127_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4786_11 (.CI(n36689), .I0(n9780[8]), .I1(GND_net), .CO(n36690));
    SB_LUT4 add_4786_10_lut (.I0(GND_net), .I1(n9780[7]), .I2(GND_net), 
            .I3(n36688), .O(n9767[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_7 (.CI(n36472), .I0(n9006[4]), .I1(n616), .CO(n36473));
    SB_LUT4 mult_14_add_1215_9_lut (.I0(GND_net), .I1(n1801[6]), .I2(GND_net), 
            .I3(n36825), .O(n1800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i459_2_lut (.I0(\Kd[7] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n683));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_14_lut (.I0(GND_net), .I1(n9201[11]), .I2(GND_net), 
            .I3(n36922), .O(n1804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3607));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[10]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4779_14_lut (.I0(GND_net), .I1(n9705[11]), .I2(GND_net), 
            .I3(n36148), .O(n9681[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_15_lut (.I0(GND_net), .I1(n8217[12]), .I2(GND_net), 
            .I3(n35685), .O(n64[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_6_lut (.I0(GND_net), .I1(n9006[3]), .I2(n519), .I3(n36471), 
            .O(n8984[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_14 (.CI(n36922), .I0(n9201[11]), .I1(GND_net), 
            .CO(n36923));
    SB_CARRY mult_14_add_1215_9 (.CI(n36825), .I0(n1801[6]), .I1(GND_net), 
            .CO(n36826));
    SB_CARRY add_4786_10 (.CI(n36688), .I0(n9780[7]), .I1(GND_net), .CO(n36689));
    SB_CARRY add_4458_6 (.CI(n36471), .I0(n9006[3]), .I1(n519), .CO(n36472));
    SB_LUT4 mult_14_add_1215_8_lut (.I0(GND_net), .I1(n1801[5]), .I2(n524), 
            .I3(n36824), .O(n1800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_9_lut (.I0(GND_net), .I1(n9780[6]), .I2(GND_net), 
            .I3(n36687), .O(n9767[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_5_lut (.I0(GND_net), .I1(n9006[2]), .I2(n422), .I3(n36470), 
            .O(n8984[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_14 (.CI(n36148), .I0(n9705[11]), .I1(GND_net), .CO(n36149));
    SB_CARRY mult_10_add_2137_15 (.CI(n35685), .I0(n8217[12]), .I1(GND_net), 
            .CO(n35686));
    SB_LUT4 mult_10_add_2137_14_lut (.I0(GND_net), .I1(n8217[11]), .I2(GND_net), 
            .I3(n35684), .O(n64[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_13_lut (.I0(GND_net), .I1(n9705[10]), .I2(GND_net), 
            .I3(n36147), .O(n9681[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_14 (.CI(n35684), .I0(n8217[11]), .I1(GND_net), 
            .CO(n35685));
    SB_CARRY unary_minus_70_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n63[0]), 
            .CO(n34743));
    SB_CARRY add_4786_9 (.CI(n36687), .I0(n9780[6]), .I1(GND_net), .CO(n36688));
    SB_LUT4 mult_14_i294_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n437));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i294_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_10_add_2137_13_lut (.I0(GND_net), .I1(n8217[10]), .I2(GND_net), 
            .I3(n35683), .O(n64[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4458_5 (.CI(n36470), .I0(n9006[2]), .I1(n422), .CO(n36471));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n467));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_8_lut (.I0(GND_net), .I1(n9780[5]), .I2(n545), .I3(n36686), 
            .O(n9767[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i379_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n564));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(n6_adj_3612), .I1(n467), .I2(n9612[2]), .I3(GND_net), 
            .O(n9577[3]));   // verilog/motorControl.v(43[17:23])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_4458_4_lut (.I0(GND_net), .I1(n9006[1]), .I2(n325), .I3(n36469), 
            .O(n8984[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_13 (.CI(n35683), .I0(n8217[10]), .I1(GND_net), 
            .CO(n35684));
    SB_CARRY add_4779_13 (.CI(n36147), .I0(n9705[10]), .I1(GND_net), .CO(n36148));
    SB_CARRY add_4458_4 (.CI(n36469), .I0(n9006[1]), .I1(n325), .CO(n36470));
    SB_LUT4 mult_10_add_2137_12_lut (.I0(GND_net), .I1(n8217[9]), .I2(GND_net), 
            .I3(n35682), .O(n64[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_13_lut (.I0(GND_net), .I1(n9201[10]), .I2(GND_net), 
            .I3(n36921), .O(n1804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_13 (.CI(n36921), .I0(n9201[10]), .I1(GND_net), 
            .CO(n36922));
    SB_LUT4 mult_14_add_1219_12_lut (.I0(GND_net), .I1(n9201[9]), .I2(GND_net), 
            .I3(n36920), .O(n1804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4458_3_lut (.I0(GND_net), .I1(n9006[0]), .I2(n228_adj_3613), 
            .I3(n36468), .O(n8984[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_12 (.CI(n36920), .I0(n9201[9]), .I1(GND_net), 
            .CO(n36921));
    SB_CARRY mult_14_add_1215_8 (.CI(n36824), .I0(n1801[5]), .I1(n524), 
            .CO(n36825));
    SB_CARRY add_4786_8 (.CI(n36686), .I0(n9780[5]), .I1(n545), .CO(n36687));
    SB_LUT4 add_4779_12_lut (.I0(GND_net), .I1(n9705[9]), .I2(GND_net), 
            .I3(n36146), .O(n9681[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_7_lut (.I0(GND_net), .I1(n1801[4]), .I2(n451_c), 
            .I3(n36823), .O(n1800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_12 (.CI(n35682), .I0(n8217[9]), .I1(GND_net), 
            .CO(n35683));
    SB_LUT4 unary_minus_23_add_3_25_lut (.I0(\PID_CONTROLLER.result [23]), 
            .I1(n49785), .I2(n61[31]), .I3(n34742), .O(n448)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_23_add_3_24_lut (.I0(\PID_CONTROLLER.result [22]), 
            .I1(n49785), .I2(n61[22]), .I3(n34741), .O(n449)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_24 (.CI(n34741), .I0(n49785), .I1(n61[22]), 
            .CO(n34742));
    SB_CARRY add_4458_3 (.CI(n36468), .I0(n9006[0]), .I1(n228_adj_3613), 
            .CO(n36469));
    SB_LUT4 mult_10_add_2137_11_lut (.I0(GND_net), .I1(n8217[8]), .I2(GND_net), 
            .I3(n35681), .O(n64[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_11 (.CI(n35681), .I0(n8217[8]), .I1(GND_net), 
            .CO(n35682));
    SB_CARRY add_4779_12 (.CI(n36146), .I0(n9705[9]), .I1(GND_net), .CO(n36147));
    SB_CARRY mult_14_add_1215_7 (.CI(n36823), .I0(n1801[4]), .I1(n451_c), 
            .CO(n36824));
    SB_LUT4 add_4779_11_lut (.I0(GND_net), .I1(n9705[8]), .I2(GND_net), 
            .I3(n36145), .O(n9681[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_11 (.CI(n36145), .I0(n9705[8]), .I1(GND_net), .CO(n36146));
    SB_LUT4 add_4458_2_lut (.I0(GND_net), .I1(n38), .I2(n131_adj_3617), 
            .I3(GND_net), .O(n8984[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4458_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_10_lut (.I0(GND_net), .I1(n8217[7]), .I2(GND_net), 
            .I3(n35680), .O(n64[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_7_lut (.I0(GND_net), .I1(n9780[4]), .I2(n472), .I3(n36685), 
            .O(n9767[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_7 (.CI(n36685), .I0(n9780[4]), .I1(n472), .CO(n36686));
    SB_CARRY add_4458_2 (.CI(GND_net), .I0(n38), .I1(n131_adj_3617), .CO(n36468));
    SB_LUT4 add_4779_10_lut (.I0(GND_net), .I1(n9705[7]), .I2(GND_net), 
            .I3(n36144), .O(n9681[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4457_22_lut (.I0(GND_net), .I1(n8984[19]), .I2(GND_net), 
            .I3(n36467), .O(n8961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_10 (.CI(n36144), .I0(n9705[7]), .I1(GND_net), .CO(n36145));
    SB_LUT4 add_4779_9_lut (.I0(GND_net), .I1(n9705[6]), .I2(GND_net), 
            .I3(n36143), .O(n9681[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_9 (.CI(n36143), .I0(n9705[6]), .I1(GND_net), .CO(n36144));
    SB_CARRY mult_10_add_2137_10 (.CI(n35680), .I0(n8217[7]), .I1(GND_net), 
            .CO(n35681));
    SB_LUT4 add_4779_8_lut (.I0(GND_net), .I1(n9705[5]), .I2(n545), .I3(n36142), 
            .O(n9681[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_6_lut (.I0(GND_net), .I1(n1801[3]), .I2(n378), 
            .I3(n36822), .O(n1800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_8 (.CI(n36142), .I0(n9705[5]), .I1(n545), .CO(n36143));
    SB_LUT4 add_4457_21_lut (.I0(GND_net), .I1(n8984[18]), .I2(GND_net), 
            .I3(n36466), .O(n8961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_21 (.CI(n36466), .I0(n8984[18]), .I1(GND_net), .CO(n36467));
    SB_LUT4 mult_10_add_2137_9_lut (.I0(GND_net), .I1(n8217[6]), .I2(GND_net), 
            .I3(n35679), .O(n64[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_7_lut (.I0(GND_net), .I1(n9705[4]), .I2(n472), .I3(n36141), 
            .O(n9681[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_9 (.CI(n35679), .I0(n8217[6]), .I1(GND_net), 
            .CO(n35680));
    SB_LUT4 add_4457_20_lut (.I0(GND_net), .I1(n8984[17]), .I2(GND_net), 
            .I3(n36465), .O(n8961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_8_lut (.I0(GND_net), .I1(n8217[5]), .I2(n680_adj_3618), 
            .I3(n35678), .O(n64[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_6_lut (.I0(GND_net), .I1(n9780[3]), .I2(n399), .I3(n36684), 
            .O(n9767[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_20 (.CI(n36465), .I0(n8984[17]), .I1(GND_net), .CO(n36466));
    SB_CARRY mult_10_add_2137_8 (.CI(n35678), .I0(n8217[5]), .I1(n680_adj_3618), 
            .CO(n35679));
    SB_CARRY add_4779_7 (.CI(n36141), .I0(n9705[4]), .I1(n472), .CO(n36142));
    SB_LUT4 add_4457_19_lut (.I0(GND_net), .I1(n8984[16]), .I2(GND_net), 
            .I3(n36464), .O(n8961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_6 (.CI(n36822), .I0(n1801[3]), .I1(n378), 
            .CO(n36823));
    SB_CARRY add_4786_6 (.CI(n36684), .I0(n9780[3]), .I1(n399), .CO(n36685));
    SB_CARRY add_4457_19 (.CI(n36464), .I0(n8984[16]), .I1(GND_net), .CO(n36465));
    SB_LUT4 add_4779_6_lut (.I0(GND_net), .I1(n9705[3]), .I2(n399), .I3(n36140), 
            .O(n9681[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_7_lut (.I0(GND_net), .I1(n8217[4]), .I2(n583_adj_3620), 
            .I3(n35677), .O(n64[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_6 (.CI(n36140), .I0(n9705[3]), .I1(n399), .CO(n36141));
    SB_CARRY mult_10_add_2137_7 (.CI(n35677), .I0(n8217[4]), .I1(n583_adj_3620), 
            .CO(n35678));
    SB_LUT4 add_4779_5_lut (.I0(GND_net), .I1(n9705[2]), .I2(n326), .I3(n36139), 
            .O(n9681[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_6_lut (.I0(GND_net), .I1(n8217[3]), .I2(n486_adj_3621), 
            .I3(n35676), .O(n64[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_6 (.CI(n35676), .I0(n8217[3]), .I1(n486_adj_3621), 
            .CO(n35677));
    SB_LUT4 mult_10_i190_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n273));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i190_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4779_5 (.CI(n36139), .I0(n9705[2]), .I1(n326), .CO(n36140));
    SB_LUT4 add_4786_5_lut (.I0(GND_net), .I1(n9780[2]), .I2(n326), .I3(n36683), 
            .O(n9767[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4457_18_lut (.I0(GND_net), .I1(n8984[15]), .I2(GND_net), 
            .I3(n36463), .O(n8961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_5_lut (.I0(GND_net), .I1(n8217[2]), .I2(n389_adj_3622), 
            .I3(n35675), .O(n64[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_4_lut (.I0(GND_net), .I1(n9705[1]), .I2(n253), .I3(n36138), 
            .O(n9681[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_18 (.CI(n36463), .I0(n8984[15]), .I1(GND_net), .CO(n36464));
    SB_LUT4 mult_10_i62_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i62_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_2137_5 (.CI(n35675), .I0(n8217[2]), .I1(n389_adj_3622), 
            .CO(n35676));
    SB_LUT4 unary_minus_23_add_3_23_lut (.I0(\PID_CONTROLLER.result [21]), 
            .I1(n49785), .I2(n61[21]), .I3(n34740), .O(n450)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4779_4 (.CI(n36138), .I0(n9705[1]), .I1(n253), .CO(n36139));
    SB_LUT4 mult_10_add_2137_4_lut (.I0(GND_net), .I1(n8217[1]), .I2(n292_adj_3624), 
            .I3(n35674), .O(n64[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_3_lut (.I0(GND_net), .I1(n9705[0]), .I2(n180_adj_3549), 
            .I3(n36137), .O(n9681[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_4 (.CI(n35674), .I0(n8217[1]), .I1(n292_adj_3624), 
            .CO(n35675));
    SB_CARRY add_4779_3 (.CI(n36137), .I0(n9705[0]), .I1(n180_adj_3549), 
            .CO(n36138));
    SB_LUT4 add_4779_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9681[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_23 (.CI(n34740), .I0(n49785), .I1(n61[21]), 
            .CO(n34741));
    SB_CARRY add_4786_5 (.CI(n36683), .I0(n9780[2]), .I1(n326), .CO(n36684));
    SB_LUT4 add_4457_17_lut (.I0(GND_net), .I1(n8984[14]), .I2(GND_net), 
            .I3(n36462), .O(n8961[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_17 (.CI(n36462), .I0(n8984[14]), .I1(GND_net), .CO(n36463));
    SB_CARRY add_4779_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36137));
    SB_LUT4 add_4782_16_lut (.I0(GND_net), .I1(n9722[13]), .I2(GND_net), 
            .I3(n36136), .O(n9705[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_3_lut (.I0(GND_net), .I1(n8217[0]), .I2(n195_adj_3625), 
            .I3(n35673), .O(n64[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_15_lut (.I0(GND_net), .I1(n9722[12]), .I2(GND_net), 
            .I3(n36135), .O(n9705[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_11_lut (.I0(GND_net), .I1(n9201[8]), .I2(GND_net), 
            .I3(n36919), .O(n1804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_3 (.CI(n35673), .I0(n8217[0]), .I1(n195_adj_3625), 
            .CO(n35674));
    SB_LUT4 mult_14_add_1215_5_lut (.I0(GND_net), .I1(n1801[2]), .I2(n305), 
            .I3(n36821), .O(n1800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_4_lut (.I0(GND_net), .I1(n9780[1]), .I2(n253), .I3(n36682), 
            .O(n9767[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_22_lut (.I0(\PID_CONTROLLER.result [20]), 
            .I1(n49785), .I2(n61[20]), .I3(n34739), .O(n451)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4457_16_lut (.I0(GND_net), .I1(n8984[13]), .I2(GND_net), 
            .I3(n36461), .O(n8961[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_22 (.CI(n34739), .I0(n49785), .I1(n61[20]), 
            .CO(n34740));
    SB_CARRY add_4786_4 (.CI(n36682), .I0(n9780[1]), .I1(n253), .CO(n36683));
    SB_CARRY add_4457_16 (.CI(n36461), .I0(n8984[13]), .I1(GND_net), .CO(n36462));
    SB_LUT4 unary_minus_23_add_3_21_lut (.I0(\PID_CONTROLLER.result[19] ), 
            .I1(n49785), .I2(n61[19]), .I3(n34738), .O(n23926)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4457_15_lut (.I0(GND_net), .I1(n8984[12]), .I2(GND_net), 
            .I3(n36460), .O(n8961[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_3_lut (.I0(GND_net), .I1(n9780[0]), .I2(n180_adj_3549), 
            .I3(n36681), .O(n9767[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_11 (.CI(n36919), .I0(n9201[8]), .I1(GND_net), 
            .CO(n36920));
    SB_CARRY add_4782_15 (.CI(n36135), .I0(n9722[12]), .I1(GND_net), .CO(n36136));
    SB_CARRY add_4457_15 (.CI(n36460), .I0(n8984[12]), .I1(GND_net), .CO(n36461));
    SB_LUT4 add_4782_14_lut (.I0(GND_net), .I1(n9722[11]), .I2(GND_net), 
            .I3(n36134), .O(n9705[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3630), .I2(n98_adj_3631), 
            .I3(GND_net), .O(n64[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_10_lut (.I0(GND_net), .I1(n9201[7]), .I2(GND_net), 
            .I3(n36918), .O(n1804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_5 (.CI(n36821), .I0(n1801[2]), .I1(n305), 
            .CO(n36822));
    SB_CARRY add_4786_3 (.CI(n36681), .I0(n9780[0]), .I1(n180_adj_3549), 
            .CO(n36682));
    SB_LUT4 add_4457_14_lut (.I0(GND_net), .I1(n8984[11]), .I2(GND_net), 
            .I3(n36459), .O(n8961[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_14 (.CI(n36134), .I0(n9722[11]), .I1(GND_net), .CO(n36135));
    SB_CARRY mult_10_add_2137_2 (.CI(GND_net), .I0(n5_adj_3630), .I1(n98_adj_3631), 
            .CO(n35673));
    SB_LUT4 add_4766_7_lut (.I0(GND_net), .I1(n44039), .I2(n658), .I3(n35672), 
            .O(n9547[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9767[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4766_6_lut (.I0(GND_net), .I1(n9584[3]), .I2(n561), .I3(n35671), 
            .O(n9547[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n370_adj_3633));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_23_add_3_21 (.CI(n34738), .I0(n49785), .I1(n61[19]), 
            .CO(n34739));
    SB_CARRY add_4766_6 (.CI(n35671), .I0(n9584[3]), .I1(n561), .CO(n35672));
    SB_LUT4 mult_14_add_1215_4_lut (.I0(GND_net), .I1(n1801[1]), .I2(n232_adj_3635), 
            .I3(n36820), .O(n1800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_14 (.CI(n36459), .I0(n8984[11]), .I1(GND_net), .CO(n36460));
    SB_CARRY mult_14_add_1215_4 (.CI(n36820), .I0(n1801[1]), .I1(n232_adj_3635), 
            .CO(n36821));
    SB_LUT4 add_4457_13_lut (.I0(GND_net), .I1(n8984[10]), .I2(GND_net), 
            .I3(n36458), .O(n8961[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29089_3_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n34094), .I2(n34487), 
            .I3(GND_net), .O(n9577[1]));   // verilog/motorControl.v(43[17:23])
    defparam i29089_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 unary_minus_23_add_3_20_lut (.I0(\PID_CONTROLLER.result [18]), 
            .I1(n49785), .I2(n61[18]), .I3(n34737), .O(n453)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4782_13_lut (.I0(GND_net), .I1(n9722[10]), .I2(GND_net), 
            .I3(n36133), .O(n9705[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_13 (.CI(n36133), .I0(n9722[10]), .I1(GND_net), .CO(n36134));
    SB_CARRY add_4786_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36681));
    SB_LUT4 mult_14_add_1215_3_lut (.I0(GND_net), .I1(n1801[0]), .I2(n159), 
            .I3(n36819), .O(n1800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4787_11_lut (.I0(GND_net), .I1(n9792[8]), .I2(GND_net), 
            .I3(n36680), .O(n9780[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_20 (.CI(n34737), .I0(n49785), .I1(n61[18]), 
            .CO(n34738));
    SB_CARRY add_4457_13 (.CI(n36458), .I0(n8984[10]), .I1(GND_net), .CO(n36459));
    SB_LUT4 add_4787_10_lut (.I0(GND_net), .I1(n9792[7]), .I2(GND_net), 
            .I3(n36679), .O(n9780[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4457_12_lut (.I0(GND_net), .I1(n8984[9]), .I2(GND_net), 
            .I3(n36457), .O(n8961[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_12 (.CI(n36457), .I0(n8984[9]), .I1(GND_net), .CO(n36458));
    SB_LUT4 add_4782_12_lut (.I0(GND_net), .I1(n9722[9]), .I2(GND_net), 
            .I3(n36132), .O(n9705[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_12 (.CI(n36132), .I0(n9722[9]), .I1(GND_net), .CO(n36133));
    SB_LUT4 unary_minus_23_add_3_19_lut (.I0(\PID_CONTROLLER.result[17] ), 
            .I1(n49785), .I2(n61[17]), .I3(n34736), .O(n23686)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4457_11_lut (.I0(GND_net), .I1(n8984[8]), .I2(GND_net), 
            .I3(n36456), .O(n8961[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_11_lut (.I0(GND_net), .I1(n9722[8]), .I2(GND_net), 
            .I3(n36131), .O(n9705[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_11 (.CI(n36456), .I0(n8984[8]), .I1(GND_net), .CO(n36457));
    SB_CARRY add_4782_11 (.CI(n36131), .I0(n9722[8]), .I1(GND_net), .CO(n36132));
    SB_LUT4 add_4782_10_lut (.I0(GND_net), .I1(n9722[7]), .I2(GND_net), 
            .I3(n36130), .O(n9705[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_10 (.CI(n36130), .I0(n9722[7]), .I1(GND_net), .CO(n36131));
    SB_CARRY add_4787_10 (.CI(n36679), .I0(n9792[7]), .I1(GND_net), .CO(n36680));
    SB_LUT4 add_4766_5_lut (.I0(GND_net), .I1(n9618[2]), .I2(n470_c), 
            .I3(n35670), .O(n9547[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4766_5 (.CI(n35670), .I0(n9618[2]), .I1(n470_c), .CO(n35671));
    SB_LUT4 add_4766_4_lut (.I0(GND_net), .I1(n9584[1]), .I2(n373), .I3(n35669), 
            .O(n9547[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4766_4 (.CI(n35669), .I0(n9584[1]), .I1(n373), .CO(n35670));
    SB_CARRY mult_14_add_1215_3 (.CI(n36819), .I0(n1801[0]), .I1(n159), 
            .CO(n36820));
    SB_CARRY unary_minus_23_add_3_19 (.CI(n34736), .I0(n49785), .I1(n61[17]), 
            .CO(n34737));
    SB_LUT4 add_4457_10_lut (.I0(GND_net), .I1(n8984[7]), .I2(GND_net), 
            .I3(n36455), .O(n8961[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_9_lut (.I0(GND_net), .I1(n9722[6]), .I2(GND_net), 
            .I3(n36129), .O(n9705[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4787_9_lut (.I0(GND_net), .I1(n9792[6]), .I2(GND_net), 
            .I3(n36678), .O(n9780[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_9 (.CI(n36129), .I0(n9722[6]), .I1(GND_net), .CO(n36130));
    SB_CARRY add_4787_9 (.CI(n36678), .I0(n9792[6]), .I1(GND_net), .CO(n36679));
    SB_LUT4 add_4766_3_lut (.I0(GND_net), .I1(n9584[0]), .I2(n276), .I3(n35668), 
            .O(n9547[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_18_lut (.I0(\PID_CONTROLLER.result [16]), 
            .I1(n49785), .I2(n61[16]), .I3(n34735), .O(n455)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4782_8_lut (.I0(GND_net), .I1(n9722[5]), .I2(n545), .I3(n36128), 
            .O(n9705[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4766_3 (.CI(n35668), .I0(n9584[0]), .I1(n276), .CO(n35669));
    SB_CARRY add_4782_8 (.CI(n36128), .I0(n9722[5]), .I1(n545), .CO(n36129));
    SB_CARRY add_4457_10 (.CI(n36455), .I0(n8984[7]), .I1(GND_net), .CO(n36456));
    SB_LUT4 add_4457_9_lut (.I0(GND_net), .I1(n8984[6]), .I2(GND_net), 
            .I3(n36454), .O(n8961[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4787_8_lut (.I0(GND_net), .I1(n9792[5]), .I2(n545), .I3(n36677), 
            .O(n9780[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4766_2_lut (.I0(GND_net), .I1(n83), .I2(n179), .I3(GND_net), 
            .O(n9547[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_7_lut (.I0(GND_net), .I1(n9722[4]), .I2(n472), .I3(n36127), 
            .O(n9705[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4766_2 (.CI(GND_net), .I0(n83), .I1(n179), .CO(n35668));
    SB_LUT4 add_4424_31_lut (.I0(GND_net), .I1(n8249[28]), .I2(GND_net), 
            .I3(n35667), .O(n8217[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i440_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n655));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4424_30_lut (.I0(GND_net), .I1(n8249[27]), .I2(GND_net), 
            .I3(n35666), .O(n8217[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4787_8 (.CI(n36677), .I0(n9792[5]), .I1(n545), .CO(n36678));
    SB_CARRY add_4457_9 (.CI(n36454), .I0(n8984[6]), .I1(GND_net), .CO(n36455));
    SB_CARRY mult_14_add_1219_10 (.CI(n36918), .I0(n9201[7]), .I1(GND_net), 
            .CO(n36919));
    SB_CARRY add_4782_7 (.CI(n36127), .I0(n9722[4]), .I1(n472), .CO(n36128));
    SB_CARRY add_4424_30 (.CI(n35666), .I0(n8249[27]), .I1(GND_net), .CO(n35667));
    SB_LUT4 add_4457_8_lut (.I0(GND_net), .I1(n8984[5]), .I2(n710), .I3(n36453), 
            .O(n8961[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_29_lut (.I0(GND_net), .I1(n8249[26]), .I2(GND_net), 
            .I3(n35665), .O(n8217[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_18 (.CI(n34735), .I0(n49785), .I1(n61[16]), 
            .CO(n34736));
    SB_LUT4 i28783_4_lut (.I0(n9612[2]), .I1(\Kp[4] ), .I2(n6_adj_3612), 
            .I3(\PID_CONTROLLER.err[31] ), .O(n8_adj_3640));   // verilog/motorControl.v(43[17:23])
    defparam i28783_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_14_add_1219_9_lut (.I0(GND_net), .I1(n9201[6]), .I2(GND_net), 
            .I3(n36917), .O(n1804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_2_lut (.I0(GND_net), .I1(n17_adj_3642), .I2(n86), 
            .I3(GND_net), .O(n1800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4787_7_lut (.I0(GND_net), .I1(n9792[4]), .I2(n472), .I3(n36676), 
            .O(n9780[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_8 (.CI(n36453), .I0(n8984[5]), .I1(n710), .CO(n36454));
    SB_LUT4 add_4782_6_lut (.I0(GND_net), .I1(n9722[3]), .I2(n399), .I3(n36126), 
            .O(n9705[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_17_lut (.I0(\PID_CONTROLLER.result [15]), 
            .I1(n49785), .I2(n61[15]), .I3(n34734), .O(n456)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mult_14_add_1215_2 (.CI(GND_net), .I0(n17_adj_3642), .I1(n86), 
            .CO(n36819));
    SB_CARRY add_4787_7 (.CI(n36676), .I0(n9792[4]), .I1(n472), .CO(n36677));
    SB_CARRY add_4424_29 (.CI(n35665), .I0(n8249[26]), .I1(GND_net), .CO(n35666));
    SB_LUT4 add_4457_7_lut (.I0(GND_net), .I1(n8984[4]), .I2(n613), .I3(n36452), 
            .O(n8961[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_6 (.CI(n36126), .I0(n9722[3]), .I1(n399), .CO(n36127));
    SB_LUT4 add_4424_28_lut (.I0(GND_net), .I1(n8249[25]), .I2(GND_net), 
            .I3(n35664), .O(n8217[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_5_lut (.I0(GND_net), .I1(n9722[2]), .I2(n326), .I3(n36125), 
            .O(n9705[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_5 (.CI(n36125), .I0(n9722[2]), .I1(n326), .CO(n36126));
    SB_CARRY add_4424_28 (.CI(n35664), .I0(n8249[25]), .I1(GND_net), .CO(n35665));
    SB_LUT4 add_4782_4_lut (.I0(GND_net), .I1(n9722[1]), .I2(n253), .I3(n36124), 
            .O(n9705[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_24_lut (.I0(GND_net), .I1(n1800[21]), .I2(GND_net), 
            .I3(n36817), .O(n1799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_27_lut (.I0(GND_net), .I1(n8249[24]), .I2(GND_net), 
            .I3(n35663), .O(n8217[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_4 (.CI(n36124), .I0(n9722[1]), .I1(n253), .CO(n36125));
    SB_CARRY add_4424_27 (.CI(n35663), .I0(n8249[24]), .I1(GND_net), .CO(n35664));
    SB_LUT4 i28718_4_lut (.I0(n9577[1]), .I1(\Kp[3] ), .I2(n4_adj_3644), 
            .I3(\PID_CONTROLLER.err[31] ), .O(n6_adj_3645));   // verilog/motorControl.v(43[17:23])
    defparam i28718_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4424_26_lut (.I0(GND_net), .I1(n8249[23]), .I2(GND_net), 
            .I3(n35662), .O(n8217[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_9 (.CI(n36917), .I0(n9201[6]), .I1(GND_net), 
            .CO(n36918));
    SB_CARRY mult_14_add_1214_24 (.CI(n36817), .I0(n1800[21]), .I1(GND_net), 
            .CO(n1695));
    SB_LUT4 add_4787_6_lut (.I0(GND_net), .I1(n9792[3]), .I2(n399), .I3(n36675), 
            .O(n9780[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_7 (.CI(n36452), .I0(n8984[4]), .I1(n613), .CO(n36453));
    SB_LUT4 i5_4_lut (.I0(n34487), .I1(\Kp[3] ), .I2(\Kp[4] ), .I3(\Kp[5] ), 
            .O(n44310));   // verilog/motorControl.v(43[17:23])
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 add_4782_3_lut (.I0(GND_net), .I1(n9722[0]), .I2(n180_adj_3549), 
            .I3(n36123), .O(n9705[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_3 (.CI(n36123), .I0(n9722[0]), .I1(n180_adj_3549), 
            .CO(n36124));
    SB_LUT4 i6_4_lut (.I0(n34094), .I1(n6_adj_3645), .I2(n4_adj_3646), 
            .I3(n8_adj_3640), .O(n14_adj_3647));   // verilog/motorControl.v(43[17:23])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4457_6_lut (.I0(GND_net), .I1(n8984[3]), .I2(n516_adj_3648), 
            .I3(n36451), .O(n8961[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9705[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36123));
    SB_CARRY add_4457_6 (.CI(n36451), .I0(n8984[3]), .I1(n516_adj_3648), 
            .CO(n36452));
    SB_LUT4 i7_3_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n14_adj_3647), 
            .I2(n44310), .I3(GND_net), .O(n43598));   // verilog/motorControl.v(43[17:23])
    defparam i7_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 add_4457_5_lut (.I0(GND_net), .I1(n8984[2]), .I2(n419), .I3(n36450), 
            .O(n8961[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_26 (.CI(n35662), .I0(n8249[23]), .I1(GND_net), .CO(n35663));
    SB_LUT4 add_4448_31_lut (.I0(GND_net), .I1(n8741[28]), .I2(GND_net), 
            .I3(n36122), .O(n8709[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_30_lut (.I0(GND_net), .I1(n8741[27]), .I2(GND_net), 
            .I3(n36121), .O(n8709[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_30 (.CI(n36121), .I0(n8741[27]), .I1(GND_net), .CO(n36122));
    SB_LUT4 add_4424_25_lut (.I0(GND_net), .I1(n8249[22]), .I2(GND_net), 
            .I3(n35661), .O(n8217[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_25 (.CI(n35661), .I0(n8249[22]), .I1(GND_net), .CO(n35662));
    SB_CARRY add_4457_5 (.CI(n36450), .I0(n8984[2]), .I1(n419), .CO(n36451));
    SB_LUT4 add_4448_29_lut (.I0(GND_net), .I1(n8741[26]), .I2(GND_net), 
            .I3(n36120), .O(n8709[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_24_lut (.I0(GND_net), .I1(n8249[21]), .I2(GND_net), 
            .I3(n35660), .O(n8217[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_24 (.CI(n35660), .I0(n8249[21]), .I1(GND_net), .CO(n35661));
    SB_LUT4 add_4424_23_lut (.I0(GND_net), .I1(n8249[20]), .I2(GND_net), 
            .I3(n35659), .O(n8217[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_29 (.CI(n36120), .I0(n8741[26]), .I1(GND_net), .CO(n36121));
    SB_CARRY add_4424_23 (.CI(n35659), .I0(n8249[20]), .I1(GND_net), .CO(n35660));
    SB_LUT4 add_4424_22_lut (.I0(GND_net), .I1(n8249[19]), .I2(GND_net), 
            .I3(n35658), .O(n8217[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_22 (.CI(n35658), .I0(n8249[19]), .I1(GND_net), .CO(n35659));
    SB_LUT4 unary_minus_21_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[11]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4787_6 (.CI(n36675), .I0(n9792[3]), .I1(n399), .CO(n36676));
    SB_LUT4 add_4457_4_lut (.I0(GND_net), .I1(n8984[1]), .I2(n322), .I3(n36449), 
            .O(n8961[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_4 (.CI(n36449), .I0(n8984[1]), .I1(n322), .CO(n36450));
    SB_LUT4 add_4448_28_lut (.I0(GND_net), .I1(n8741[25]), .I2(GND_net), 
            .I3(n36119), .O(n8709[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_17 (.CI(n34734), .I0(n49785), .I1(n61[15]), 
            .CO(n34735));
    SB_LUT4 add_4424_21_lut (.I0(GND_net), .I1(n8249[18]), .I2(GND_net), 
            .I3(n35657), .O(n8217[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_8_lut (.I0(GND_net), .I1(n9201[5]), .I2(n536), 
            .I3(n36916), .O(n1804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_23_lut (.I0(GND_net), .I1(n1800[20]), .I2(GND_net), 
            .I3(n36816), .O(n1799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3650));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_28678_33_lut (.I0(GND_net), .I1(n66[31]), .I2(n6817[0]), 
            .I3(n34898), .O(\PID_CONTROLLER.result_31__N_3353 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_8 (.CI(n36916), .I0(n9201[5]), .I1(n536), 
            .CO(n36917));
    SB_CARRY add_4424_21 (.CI(n35657), .I0(n8249[18]), .I1(GND_net), .CO(n35658));
    SB_LUT4 add_4424_20_lut (.I0(GND_net), .I1(n8249[17]), .I2(GND_net), 
            .I3(n35656), .O(n8217[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3651));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3652));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_7_lut (.I0(GND_net), .I1(n9201[4]), .I2(n463_c), 
            .I3(n36915), .O(n1804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_23 (.CI(n36816), .I0(n1800[20]), .I1(GND_net), 
            .CO(n36817));
    SB_CARRY add_4448_28 (.CI(n36119), .I0(n8741[25]), .I1(GND_net), .CO(n36120));
    SB_LUT4 add_4787_5_lut (.I0(GND_net), .I1(n9792[2]), .I2(n326), .I3(n36674), 
            .O(n9780[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i199_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n295_adj_3653));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i199_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4424_20 (.CI(n35656), .I0(n8249[17]), .I1(GND_net), .CO(n35657));
    SB_LUT4 add_4457_3_lut (.I0(GND_net), .I1(n8984[0]), .I2(n225_adj_3654), 
            .I3(n36448), .O(n8961[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_27_lut (.I0(GND_net), .I1(n8741[24]), .I2(GND_net), 
            .I3(n36118), .O(n8709[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_27 (.CI(n36118), .I0(n8741[24]), .I1(GND_net), .CO(n36119));
    SB_CARRY add_4787_5 (.CI(n36674), .I0(n9792[2]), .I1(n326), .CO(n36675));
    SB_CARRY add_4457_3 (.CI(n36448), .I0(n8984[0]), .I1(n225_adj_3654), 
            .CO(n36449));
    SB_LUT4 add_4457_2_lut (.I0(GND_net), .I1(n35_adj_3655), .I2(n128_adj_3656), 
            .I3(GND_net), .O(n8961[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4457_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_19_lut (.I0(GND_net), .I1(n8249[16]), .I2(GND_net), 
            .I3(n35655), .O(n8217[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_19 (.CI(n35655), .I0(n8249[16]), .I1(GND_net), .CO(n35656));
    SB_LUT4 add_4448_26_lut (.I0(GND_net), .I1(n8741[23]), .I2(GND_net), 
            .I3(n36117), .O(n8709[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i264_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n392_adj_3657));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i343_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n510_adj_3658));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i343_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_add_1214_22_lut (.I0(GND_net), .I1(n1800[19]), .I2(GND_net), 
            .I3(n36815), .O(n1799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_16_lut (.I0(\PID_CONTROLLER.result [14]), 
            .I1(n49785), .I2(n61[14]), .I3(n34733), .O(n457)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4424_18_lut (.I0(GND_net), .I1(n8249[15]), .I2(GND_net), 
            .I3(n35654), .O(n8217[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4457_2 (.CI(GND_net), .I0(n35_adj_3655), .I1(n128_adj_3656), 
            .CO(n36448));
    SB_LUT4 add_4456_23_lut (.I0(GND_net), .I1(n8961[20]), .I2(GND_net), 
            .I3(n36447), .O(n8937[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4787_4_lut (.I0(GND_net), .I1(n9792[1]), .I2(n253), .I3(n36673), 
            .O(n9780[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_18 (.CI(n35654), .I0(n8249[15]), .I1(GND_net), .CO(n35655));
    SB_LUT4 add_4424_17_lut (.I0(GND_net), .I1(n8249[14]), .I2(GND_net), 
            .I3(n35653), .O(n8217[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i280_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n416_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[16]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n513));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n610));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i422_2_lut (.I0(\Kd[6] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n628));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4448_26 (.CI(n36117), .I0(n8741[23]), .I1(GND_net), .CO(n36118));
    SB_LUT4 add_4456_22_lut (.I0(GND_net), .I1(n8961[19]), .I2(GND_net), 
            .I3(n36446), .O(n8937[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_17 (.CI(n35653), .I0(n8249[14]), .I1(GND_net), .CO(n35654));
    SB_LUT4 mult_10_i329_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n489_adj_3660));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i329_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_7 (.CI(n36915), .I0(n9201[4]), .I1(n463_c), 
            .CO(n36916));
    SB_CARRY mult_14_add_1214_22 (.CI(n36815), .I0(n1800[19]), .I1(GND_net), 
            .CO(n36816));
    SB_LUT4 add_4424_16_lut (.I0(GND_net), .I1(n8249[13]), .I2(GND_net), 
            .I3(n35652), .O(n8217[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n586_adj_3661));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_28678_32_lut (.I0(GND_net), .I1(n66[30]), .I2(n191[30]), 
            .I3(n34897), .O(\PID_CONTROLLER.result_31__N_3353 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i392_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3662));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i392_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_4456_22 (.CI(n36446), .I0(n8961[19]), .I1(GND_net), .CO(n36447));
    SB_CARRY add_4787_4 (.CI(n36673), .I0(n9792[1]), .I1(n253), .CO(n36674));
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n683_adj_3663));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4456_21_lut (.I0(GND_net), .I1(n8961[18]), .I2(GND_net), 
            .I3(n36445), .O(n8937[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_16 (.CI(n34733), .I0(n49785), .I1(n61[14]), 
            .CO(n34734));
    SB_LUT4 mult_14_add_1219_6_lut (.I0(GND_net), .I1(n9201[3]), .I2(n390), 
            .I3(n36914), .O(n1804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_25_lut (.I0(GND_net), .I1(n8741[22]), .I2(GND_net), 
            .I3(n36116), .O(n8709[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[12]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[13]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1214_21_lut (.I0(GND_net), .I1(n1800[18]), .I2(GND_net), 
            .I3(n36814), .O(n1799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_15_lut (.I0(\PID_CONTROLLER.result[13] ), 
            .I1(n49785), .I2(n61[13]), .I3(n34732), .O(n23155)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4424_16 (.CI(n35652), .I0(n8249[13]), .I1(GND_net), .CO(n35653));
    SB_CARRY add_4456_21 (.CI(n36445), .I0(n8961[18]), .I1(GND_net), .CO(n36446));
    SB_CARRY add_4448_25 (.CI(n36116), .I0(n8741[22]), .I1(GND_net), .CO(n36117));
    SB_LUT4 add_4424_15_lut (.I0(GND_net), .I1(n8249[12]), .I2(GND_net), 
            .I3(n35651), .O(n8217[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_15 (.CI(n35651), .I0(n8249[12]), .I1(GND_net), .CO(n35652));
    SB_LUT4 add_4456_20_lut (.I0(GND_net), .I1(n8961[17]), .I2(GND_net), 
            .I3(n36444), .O(n8937[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_14_lut (.I0(GND_net), .I1(n8249[11]), .I2(GND_net), 
            .I3(n35650), .O(n8217[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_24_lut (.I0(GND_net), .I1(n8741[21]), .I2(GND_net), 
            .I3(n36115), .O(n8709[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_24 (.CI(n36115), .I0(n8741[21]), .I1(GND_net), .CO(n36116));
    SB_LUT4 mult_14_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4448_23_lut (.I0(GND_net), .I1(n8741[20]), .I2(GND_net), 
            .I3(n36114), .O(n8709[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_6 (.CI(n36914), .I0(n9201[3]), .I1(n390), 
            .CO(n36915));
    SB_LUT4 add_4787_3_lut (.I0(GND_net), .I1(n9792[0]), .I2(n180_adj_3549), 
            .I3(n36672), .O(n9780[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_20 (.CI(n36444), .I0(n8961[17]), .I1(GND_net), .CO(n36445));
    SB_CARRY add_4424_14 (.CI(n35650), .I0(n8249[11]), .I1(GND_net), .CO(n35651));
    SB_CARRY add_4787_3 (.CI(n36672), .I0(n9792[0]), .I1(n180_adj_3549), 
            .CO(n36673));
    SB_CARRY add_4448_23 (.CI(n36114), .I0(n8741[20]), .I1(GND_net), .CO(n36115));
    SB_LUT4 add_4448_22_lut (.I0(GND_net), .I1(n8741[19]), .I2(GND_net), 
            .I3(n36113), .O(n8709[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_13_lut (.I0(GND_net), .I1(n8249[10]), .I2(GND_net), 
            .I3(n35649), .O(n8217[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_13 (.CI(n35649), .I0(n8249[10]), .I1(GND_net), .CO(n35650));
    SB_CARRY add_4448_22 (.CI(n36113), .I0(n8741[19]), .I1(GND_net), .CO(n36114));
    SB_LUT4 add_4424_12_lut (.I0(GND_net), .I1(n8249[9]), .I2(GND_net), 
            .I3(n35648), .O(n8217[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i475_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n707));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4456_19_lut (.I0(GND_net), .I1(n8961[16]), .I2(GND_net), 
            .I3(n36443), .O(n8937[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_21_lut (.I0(GND_net), .I1(n8741[18]), .I2(GND_net), 
            .I3(n36112), .O(n8709[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_32 (.CI(n34897), .I0(n66[30]), .I1(n191[30]), .CO(n34898));
    SB_LUT4 add_4787_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9780[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4787_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_12 (.CI(n35648), .I0(n8249[9]), .I1(GND_net), .CO(n35649));
    SB_CARRY add_4448_21 (.CI(n36112), .I0(n8741[18]), .I1(GND_net), .CO(n36113));
    SB_LUT4 add_4424_11_lut (.I0(GND_net), .I1(n8249[8]), .I2(GND_net), 
            .I3(n35647), .O(n8217[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_11 (.CI(n35647), .I0(n8249[8]), .I1(GND_net), .CO(n35648));
    SB_LUT4 unary_minus_21_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[14]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i87_2_lut (.I0(\Kd[1] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n128_adj_3656));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4448_20_lut (.I0(GND_net), .I1(n8741[17]), .I2(GND_net), 
            .I3(n36111), .O(n8709[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_19 (.CI(n36443), .I0(n8961[16]), .I1(GND_net), .CO(n36444));
    SB_CARRY add_4448_20 (.CI(n36111), .I0(n8741[17]), .I1(GND_net), .CO(n36112));
    SB_LUT4 add_4424_10_lut (.I0(GND_net), .I1(n8249[7]), .I2(GND_net), 
            .I3(n35646), .O(n8217[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_10 (.CI(n35646), .I0(n8249[7]), .I1(GND_net), .CO(n35647));
    SB_LUT4 mult_12_i24_2_lut (.I0(\Kd[0] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3655));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4424_9_lut (.I0(GND_net), .I1(n8249[6]), .I2(GND_net), 
            .I3(n35645), .O(n8217[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_19_lut (.I0(GND_net), .I1(n8741[16]), .I2(GND_net), 
            .I3(n36110), .O(n8709[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_15 (.CI(n34732), .I0(n49785), .I1(n61[13]), 
            .CO(n34733));
    SB_LUT4 unary_minus_23_add_3_14_lut (.I0(\PID_CONTROLLER.result [12]), 
            .I1(n49785), .I2(n61[12]), .I3(n34731), .O(n459)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mult_12_i152_2_lut (.I0(\Kd[2] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n225_adj_3654));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4424_9 (.CI(n35645), .I0(n8249[6]), .I1(GND_net), .CO(n35646));
    SB_LUT4 add_4424_8_lut (.I0(GND_net), .I1(n8249[5]), .I2(n683_adj_3663), 
            .I3(n35644), .O(n8217[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4787_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36672));
    SB_LUT4 mult_12_i217_2_lut (.I0(\Kd[3] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4788_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(n36671), .O(n9792[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_18_lut (.I0(GND_net), .I1(n8961[15]), .I2(GND_net), 
            .I3(n36442), .O(n8937[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_18 (.CI(n36442), .I0(n8961[15]), .I1(GND_net), .CO(n36443));
    SB_CARRY add_4448_19 (.CI(n36110), .I0(n8741[16]), .I1(GND_net), .CO(n36111));
    SB_CARRY add_4424_8 (.CI(n35644), .I0(n8249[5]), .I1(n683_adj_3663), 
            .CO(n35645));
    SB_LUT4 mult_12_i282_2_lut (.I0(\Kd[4] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n419));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4448_18_lut (.I0(GND_net), .I1(n8741[15]), .I2(GND_net), 
            .I3(n36109), .O(n8709[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_18 (.CI(n36109), .I0(n8741[15]), .I1(GND_net), .CO(n36110));
    SB_LUT4 add_4456_17_lut (.I0(GND_net), .I1(n8961[14]), .I2(GND_net), 
            .I3(n36441), .O(n8937[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4788_9_lut (.I0(GND_net), .I1(n583_adj_3662), .I2(GND_net), 
            .I3(n36670), .O(n9792[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_7_lut (.I0(GND_net), .I1(n8249[4]), .I2(n586_adj_3661), 
            .I3(n35643), .O(n8217[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_17_lut (.I0(GND_net), .I1(n8741[14]), .I2(GND_net), 
            .I3(n36108), .O(n8709[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_17 (.CI(n36108), .I0(n8741[14]), .I1(GND_net), .CO(n36109));
    SB_LUT4 mult_14_add_1219_5_lut (.I0(GND_net), .I1(n9201[2]), .I2(n317), 
            .I3(n36913), .O(n1804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_21 (.CI(n36814), .I0(n1800[18]), .I1(GND_net), 
            .CO(n36815));
    SB_CARRY add_4456_17 (.CI(n36441), .I0(n8961[14]), .I1(GND_net), .CO(n36442));
    SB_CARRY add_4424_7 (.CI(n35643), .I0(n8249[4]), .I1(n586_adj_3661), 
            .CO(n35644));
    SB_CARRY add_4788_9 (.CI(n36670), .I0(n583_adj_3662), .I1(GND_net), 
            .CO(n36671));
    SB_LUT4 add_4456_16_lut (.I0(GND_net), .I1(n8961[13]), .I2(GND_net), 
            .I3(n36440), .O(n8937[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_16_lut (.I0(GND_net), .I1(n8741[13]), .I2(GND_net), 
            .I3(n36107), .O(n8709[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4424_6_lut (.I0(GND_net), .I1(n8249[3]), .I2(n489_adj_3660), 
            .I3(n35642), .O(n8217[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_16 (.CI(n36107), .I0(n8741[13]), .I1(GND_net), .CO(n36108));
    SB_LUT4 mult_12_i347_2_lut (.I0(\Kd[5] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n516_adj_3648));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4788_8_lut (.I0(GND_net), .I1(n510_adj_3658), .I2(n545), 
            .I3(n36669), .O(n9792[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_16 (.CI(n36440), .I0(n8961[13]), .I1(GND_net), .CO(n36441));
    SB_LUT4 mult_12_i412_2_lut (.I0(\Kd[6] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[15]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4448_15_lut (.I0(GND_net), .I1(n8741[12]), .I2(GND_net), 
            .I3(n36106), .O(n8709[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_15 (.CI(n36106), .I0(n8741[12]), .I1(GND_net), .CO(n36107));
    SB_LUT4 add_4448_14_lut (.I0(GND_net), .I1(n8741[11]), .I2(GND_net), 
            .I3(n36105), .O(n8709[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_15_lut (.I0(GND_net), .I1(n8961[12]), .I2(GND_net), 
            .I3(n36439), .O(n8937[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_6 (.CI(n35642), .I0(n8249[3]), .I1(n489_adj_3660), 
            .CO(n35643));
    SB_LUT4 add_4424_5_lut (.I0(GND_net), .I1(n8249[2]), .I2(n392_adj_3657), 
            .I3(n35641), .O(n8217[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_14 (.CI(n36105), .I0(n8741[11]), .I1(GND_net), .CO(n36106));
    SB_CARRY add_4456_15 (.CI(n36439), .I0(n8961[12]), .I1(GND_net), .CO(n36440));
    SB_LUT4 add_4448_13_lut (.I0(GND_net), .I1(n8741[10]), .I2(GND_net), 
            .I3(n36104), .O(n8709[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4424_5 (.CI(n35641), .I0(n8249[2]), .I1(n392_adj_3657), 
            .CO(n35642));
    SB_LUT4 add_4424_4_lut (.I0(GND_net), .I1(n8249[1]), .I2(n295_adj_3653), 
            .I3(n35640), .O(n8217[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_4 (.CI(n35640), .I0(n8249[1]), .I1(n295_adj_3653), 
            .CO(n35641));
    SB_CARRY add_4788_8 (.CI(n36669), .I0(n510_adj_3658), .I1(n545), .CO(n36670));
    SB_LUT4 mult_14_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3642));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i477_2_lut (.I0(\Kd[7] ), .I1(n58[10]), .I2(GND_net), 
            .I3(GND_net), .O(n710));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4424_3_lut (.I0(GND_net), .I1(n8249[0]), .I2(n198_adj_3652), 
            .I3(n35639), .O(n8217[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_14_lut (.I0(GND_net), .I1(n8961[11]), .I2(GND_net), 
            .I3(n36438), .O(n8937[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_13 (.CI(n36104), .I0(n8741[10]), .I1(GND_net), .CO(n36105));
    SB_LUT4 add_28678_31_lut (.I0(GND_net), .I1(n66[29]), .I2(n191[29]), 
            .I3(n34896), .O(\PID_CONTROLLER.result_31__N_3353 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4424_3 (.CI(n35639), .I0(n8249[0]), .I1(n198_adj_3652), 
            .CO(n35640));
    SB_LUT4 add_4424_2_lut (.I0(GND_net), .I1(n8_adj_3651), .I2(n101_adj_3650), 
            .I3(GND_net), .O(n8217[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4424_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_14 (.CI(n34731), .I0(n49785), .I1(n61[12]), 
            .CO(n34732));
    SB_LUT4 unary_minus_23_add_3_13_lut (.I0(\PID_CONTROLLER.result [11]), 
            .I1(n49785), .I2(n61[11]), .I3(n34730), .O(n460)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4424_2 (.CI(GND_net), .I0(n8_adj_3651), .I1(n101_adj_3650), 
            .CO(n35639));
    SB_LUT4 mult_12_i127_2_lut (.I0(\Kd[1] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n179));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i127_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4765_7_lut (.I0(GND_net), .I1(n43598), .I2(n655), .I3(n35638), 
            .O(n9539[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_5 (.CI(n36913), .I0(n9201[2]), .I1(n317), 
            .CO(n36914));
    SB_CARRY add_4456_14 (.CI(n36438), .I0(n8961[11]), .I1(GND_net), .CO(n36439));
    SB_LUT4 add_4456_13_lut (.I0(GND_net), .I1(n8961[10]), .I2(GND_net), 
            .I3(n36437), .O(n8937[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_13 (.CI(n36437), .I0(n8961[10]), .I1(GND_net), .CO(n36438));
    SB_LUT4 add_4448_12_lut (.I0(GND_net), .I1(n8741[9]), .I2(GND_net), 
            .I3(n36103), .O(n8709[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_12_lut (.I0(GND_net), .I1(n8961[9]), .I2(GND_net), 
            .I3(n36436), .O(n8937[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_12 (.CI(n36103), .I0(n8741[9]), .I1(GND_net), .CO(n36104));
    SB_LUT4 add_4765_6_lut (.I0(GND_net), .I1(n9577[3]), .I2(n564), .I3(n35637), 
            .O(n9539[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_20_lut (.I0(GND_net), .I1(n1800[17]), .I2(GND_net), 
            .I3(n36813), .O(n1799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[16]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4765_6 (.CI(n35637), .I0(n9577[3]), .I1(n564), .CO(n35638));
    SB_LUT4 mult_12_i190_2_lut (.I0(\Kd[2] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n276));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i190_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4448_11_lut (.I0(GND_net), .I1(n8741[8]), .I2(GND_net), 
            .I3(n36102), .O(n8709[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_11 (.CI(n36102), .I0(n8741[8]), .I1(GND_net), .CO(n36103));
    SB_CARRY add_28678_31 (.CI(n34896), .I0(n66[29]), .I1(n191[29]), .CO(n34897));
    SB_LUT4 add_4448_10_lut (.I0(GND_net), .I1(n8741[7]), .I2(GND_net), 
            .I3(n36101), .O(n8709[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4788_7_lut (.I0(GND_net), .I1(n437), .I2(n472), .I3(n36668), 
            .O(n9792[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4765_5_lut (.I0(GND_net), .I1(n9577[2]), .I2(n467), .I3(n35636), 
            .O(n9539[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4765_5 (.CI(n35636), .I0(n9577[2]), .I1(n467), .CO(n35637));
    SB_CARRY unary_minus_23_add_3_13 (.CI(n34730), .I0(n49785), .I1(n61[11]), 
            .CO(n34731));
    SB_LUT4 unary_minus_21_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[17]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[18]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3635));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_23_add_3_12_lut (.I0(\PID_CONTROLLER.result[10] ), 
            .I1(n49785), .I2(n61[10]), .I3(n34729), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4765_4_lut (.I0(GND_net), .I1(n9577[1]), .I2(n370_adj_3633), 
            .I3(n35635), .O(n9539[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4765_4 (.CI(n35635), .I0(n9577[1]), .I1(n370_adj_3633), 
            .CO(n35636));
    SB_CARRY add_4456_12 (.CI(n36436), .I0(n8961[9]), .I1(GND_net), .CO(n36437));
    SB_LUT4 add_28678_30_lut (.I0(GND_net), .I1(n66[28]), .I2(n191[28]), 
            .I3(n34895), .O(\PID_CONTROLLER.result_31__N_3353 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_11_lut (.I0(GND_net), .I1(n8961[8]), .I2(GND_net), 
            .I3(n36435), .O(n8937[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4765_3_lut (.I0(GND_net), .I1(n9577[0]), .I2(n273), .I3(n35634), 
            .O(n9539[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_10 (.CI(n36101), .I0(n8741[7]), .I1(GND_net), .CO(n36102));
    SB_CARRY unary_minus_23_add_3_12 (.CI(n34729), .I0(n49785), .I1(n61[10]), 
            .CO(n34730));
    SB_LUT4 add_4448_9_lut (.I0(GND_net), .I1(n8741[6]), .I2(GND_net), 
            .I3(n36100), .O(n8709[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4765_3 (.CI(n35634), .I0(n9577[0]), .I1(n273), .CO(n35635));
    SB_LUT4 mult_14_add_1219_4_lut (.I0(GND_net), .I1(n9201[1]), .I2(n244_adj_3607), 
            .I3(n36912), .O(n1804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_20 (.CI(n36813), .I0(n1800[17]), .I1(GND_net), 
            .CO(n36814));
    SB_CARRY add_4448_9 (.CI(n36100), .I0(n8741[6]), .I1(GND_net), .CO(n36101));
    SB_LUT4 mult_14_add_1214_19_lut (.I0(GND_net), .I1(n1800[16]), .I2(GND_net), 
            .I3(n36812), .O(n1799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4448_8_lut (.I0(GND_net), .I1(n8741[5]), .I2(n683), .I3(n36099), 
            .O(n8709[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4765_2_lut (.I0(GND_net), .I1(n80), .I2(n176), .I3(GND_net), 
            .O(n9539[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4765_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4765_2 (.CI(GND_net), .I0(n80), .I1(n176), .CO(n35634));
    SB_CARRY add_28678_30 (.CI(n34895), .I0(n66[28]), .I1(n191[28]), .CO(n34896));
    SB_CARRY add_4448_8 (.CI(n36099), .I0(n8741[5]), .I1(n683), .CO(n36100));
    SB_CARRY mult_14_add_1214_19 (.CI(n36812), .I0(n1800[16]), .I1(GND_net), 
            .CO(n36813));
    SB_CARRY add_4788_7 (.CI(n36668), .I0(n437), .I1(n472), .CO(n36669));
    SB_LUT4 mult_12_i62_2_lut (.I0(\Kd[0] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i62_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4456_11 (.CI(n36435), .I0(n8961[8]), .I1(GND_net), .CO(n36436));
    SB_LUT4 add_4448_7_lut (.I0(GND_net), .I1(n8741[4]), .I2(n586), .I3(n36098), 
            .O(n8709[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_7 (.CI(n36098), .I0(n8741[4]), .I1(n586), .CO(n36099));
    SB_LUT4 unary_minus_23_add_3_11_lut (.I0(\PID_CONTROLLER.result [9]), 
            .I1(n49785), .I2(n61[9]), .I3(n34728), .O(n462)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_11 (.CI(n34728), .I0(n49785), .I1(n61[9]), 
            .CO(n34729));
    SB_LUT4 add_4788_6_lut (.I0(GND_net), .I1(n364), .I2(n399), .I3(n36667), 
            .O(n9792[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(\Kd[2] ), .I1(\Kd[0] ), .I2(n58[25]), .I3(\Kd[1] ), 
            .O(n4_adj_3668));   // verilog/motorControl.v(43[26:45])
    defparam i2_4_lut.LUT_INIT = 16'ha080;
    SB_LUT4 add_4448_6_lut (.I0(GND_net), .I1(n8741[3]), .I2(n489), .I3(n36097), 
            .O(n8709[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_6 (.CI(n36097), .I0(n8741[3]), .I1(n489), .CO(n36098));
    SB_LUT4 mult_12_i253_2_lut (.I0(\Kd[3] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n373));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28976_3_lut (.I0(n58[25]), .I1(n34377), .I2(n34352), .I3(GND_net), 
            .O(n9584[1]));   // verilog/motorControl.v(43[26:45])
    defparam i28976_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_12_i316_2_lut (.I0(\Kd[4] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n470_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4456_10_lut (.I0(GND_net), .I1(n8961[7]), .I2(GND_net), 
            .I3(n36434), .O(n8937[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i377_2_lut (.I0(\Kd[5] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n561));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4456_10 (.CI(n36434), .I0(n8961[7]), .I1(GND_net), .CO(n36435));
    SB_LUT4 add_4456_9_lut (.I0(GND_net), .I1(n8961[6]), .I2(GND_net), 
            .I3(n36433), .O(n8937[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_4 (.CI(n36912), .I0(n9201[1]), .I1(n244_adj_3607), 
            .CO(n36913));
    SB_LUT4 add_4448_5_lut (.I0(GND_net), .I1(n8741[2]), .I2(n392), .I3(n36096), 
            .O(n8709[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4788_6 (.CI(n36667), .I0(n364), .I1(n399), .CO(n36668));
    SB_LUT4 mult_14_add_1214_18_lut (.I0(GND_net), .I1(n1800[15]), .I2(GND_net), 
            .I3(n36811), .O(n1799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_29_lut (.I0(GND_net), .I1(n66[27]), .I2(n191[27]), 
            .I3(n34894), .O(\PID_CONTROLLER.result_31__N_3353 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i487_2_lut (.I0(\Kd[7] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n725));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_23_add_3_10_lut (.I0(\PID_CONTROLLER.result [8]), 
            .I1(n49785), .I2(n61[8]), .I3(n34727), .O(n463)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mult_12_i442_2_lut (.I0(\Kd[6] ), .I1(n58[25]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i442_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4448_5 (.CI(n36096), .I0(n8741[2]), .I1(n392), .CO(n36097));
    SB_LUT4 unary_minus_17_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[17]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4448_4_lut (.I0(GND_net), .I1(n8741[1]), .I2(n295), .I3(n36095), 
            .O(n8709[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut_adj_842 (.I0(n34377), .I1(n7_adj_3670), .I2(n8_adj_3671), 
            .I3(n8_adj_3672), .O(n44039));   // verilog/motorControl.v(43[26:45])
    defparam i5_4_lut_adj_842.LUT_INIT = 16'h6996;
    SB_CARRY add_4456_9 (.CI(n36433), .I0(n8961[6]), .I1(GND_net), .CO(n36434));
    SB_LUT4 add_4456_8_lut (.I0(GND_net), .I1(n8961[5]), .I2(n707_adj_3562), 
            .I3(n36432), .O(n8937[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_18 (.CI(n36811), .I0(n1800[15]), .I1(GND_net), 
            .CO(n36812));
    SB_LUT4 add_4788_5_lut (.I0(GND_net), .I1(n291), .I2(n326), .I3(n36666), 
            .O(n9792[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_29 (.CI(n34894), .I0(n66[27]), .I1(n191[27]), .CO(n34895));
    SB_CARRY unary_minus_23_add_3_10 (.CI(n34727), .I0(n49785), .I1(n61[8]), 
            .CO(n34728));
    SB_CARRY add_4448_4 (.CI(n36095), .I0(n8741[1]), .I1(n295), .CO(n36096));
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3631));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3630));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[19]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4788_5 (.CI(n36666), .I0(n291), .I1(n326), .CO(n36667));
    SB_LUT4 add_4448_3_lut (.I0(GND_net), .I1(n8741[0]), .I2(n198), .I3(n36094), 
            .O(n8709[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_8 (.CI(n36432), .I0(n8961[5]), .I1(n707_adj_3562), 
            .CO(n36433));
    SB_LUT4 add_4456_7_lut (.I0(GND_net), .I1(n8961[4]), .I2(n610_adj_3557), 
            .I3(n36431), .O(n8937[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[20]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4448_3 (.CI(n36094), .I0(n8741[0]), .I1(n198), .CO(n36095));
    SB_LUT4 add_4448_2_lut (.I0(GND_net), .I1(n8_adj_3551), .I2(n101), 
            .I3(GND_net), .O(n8709[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4448_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4448_2 (.CI(GND_net), .I0(n8_adj_3551), .I1(n101), .CO(n36094));
    SB_LUT4 mult_14_add_1219_3_lut (.I0(GND_net), .I1(n9201[0]), .I2(n171), 
            .I3(n36911), .O(n1804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4447_8_lut (.I0(GND_net), .I1(n9539[5]), .I2(n752), .I3(n36093), 
            .O(n8700[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4447_7_lut (.I0(GND_net), .I1(n9539[4]), .I2(n655), .I3(n36092), 
            .O(n8700[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4788_4_lut (.I0(GND_net), .I1(n218_adj_3548), .I2(n253), 
            .I3(n36665), .O(n9792[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_7 (.CI(n36431), .I0(n8961[4]), .I1(n610_adj_3557), 
            .CO(n36432));
    SB_CARRY add_4447_7 (.CI(n36092), .I0(n9539[4]), .I1(n655), .CO(n36093));
    SB_LUT4 add_4447_6_lut (.I0(GND_net), .I1(n9539[3]), .I2(n564), .I3(n36091), 
            .O(n8700[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_6_lut (.I0(GND_net), .I1(n8961[3]), .I2(n513_adj_3544), 
            .I3(n36430), .O(n8937[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_17_lut (.I0(GND_net), .I1(n1800[14]), .I2(GND_net), 
            .I3(n36810), .O(n1799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4447_6 (.CI(n36091), .I0(n9539[3]), .I1(n564), .CO(n36092));
    SB_CARRY add_4788_4 (.CI(n36665), .I0(n218_adj_3548), .I1(n253), .CO(n36666));
    SB_LUT4 add_4447_5_lut (.I0(GND_net), .I1(n9539[2]), .I2(n467), .I3(n36090), 
            .O(n8700[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4456_6 (.CI(n36430), .I0(n8961[3]), .I1(n513_adj_3544), 
            .CO(n36431));
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3625));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4447_5 (.CI(n36090), .I0(n9539[2]), .I1(n467), .CO(n36091));
    SB_LUT4 add_4447_4_lut (.I0(GND_net), .I1(n9539[1]), .I2(n370_adj_3633), 
            .I3(n36089), .O(n8700[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4456_5_lut (.I0(GND_net), .I1(n8961[2]), .I2(n416_adj_3536), 
            .I3(n36429), .O(n8937[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_3 (.CI(n36911), .I0(n9201[0]), .I1(n171), 
            .CO(n36912));
    SB_CARRY add_4447_4 (.CI(n36089), .I0(n9539[1]), .I1(n370_adj_3633), 
            .CO(n36090));
    SB_LUT4 add_28678_28_lut (.I0(GND_net), .I1(n66[26]), .I2(n191[26]), 
            .I3(n34893), .O(\PID_CONTROLLER.result_31__N_3353 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_17 (.CI(n36810), .I0(n1800[14]), .I1(GND_net), 
            .CO(n36811));
    SB_LUT4 unary_minus_23_add_3_9_lut (.I0(\PID_CONTROLLER.result [7]), .I1(n49785), 
            .I2(n61[7]), .I3(n34726), .O(n464)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4447_3_lut (.I0(GND_net), .I1(n9539[0]), .I2(n273), .I3(n36088), 
            .O(n8700[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4447_3 (.CI(n36088), .I0(n9539[0]), .I1(n273), .CO(n36089));
    SB_LUT4 add_4447_2_lut (.I0(GND_net), .I1(n80), .I2(n176), .I3(GND_net), 
            .O(n8700[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4447_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n98_adj_3534), 
            .I3(GND_net), .O(n1804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_16_lut (.I0(GND_net), .I1(n1800[13]), .I2(GND_net), 
            .I3(n36809), .O(n1799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n695));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i197_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n292_adj_3624));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[21]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4788_3_lut (.I0(GND_net), .I1(n145), .I2(n180_adj_3549), 
            .I3(n36664), .O(n9792[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_9 (.CI(n34726), .I0(n49785), .I1(n61[7]), 
            .CO(n34727));
    SB_CARRY add_4456_5 (.CI(n36429), .I0(n8961[2]), .I1(n416_adj_3536), 
            .CO(n36430));
    SB_LUT4 add_4456_4_lut (.I0(GND_net), .I1(n8961[1]), .I2(n319_adj_3530), 
            .I3(n36428), .O(n8937[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4447_2 (.CI(GND_net), .I0(n80), .I1(n176), .CO(n36088));
    SB_CARRY add_4456_4 (.CI(n36428), .I0(n8961[1]), .I1(n319_adj_3530), 
            .CO(n36429));
    SB_LUT4 add_4446_9_lut (.I0(GND_net), .I1(n8700[6]), .I2(GND_net), 
            .I3(n36087), .O(n8690[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_8_lut (.I0(GND_net), .I1(n8700[5]), .I2(n749), .I3(n36086), 
            .O(n8690[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4788_3 (.CI(n36664), .I0(n145), .I1(n180_adj_3549), .CO(n36665));
    SB_CARRY mult_14_add_1219_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n98_adj_3534), 
            .CO(n36911));
    SB_LUT4 mult_10_i262_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n389_adj_3622));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4788_2_lut (.I0(GND_net), .I1(n72), .I2(n107), .I3(GND_net), 
            .O(n9792[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4788_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_8 (.CI(n36086), .I0(n8700[5]), .I1(n749), .CO(n36087));
    SB_CARRY add_28678_28 (.CI(n34893), .I0(n66[26]), .I1(n191[26]), .CO(n34894));
    SB_CARRY mult_14_add_1214_16 (.CI(n36809), .I0(n1800[13]), .I1(GND_net), 
            .CO(n36810));
    SB_LUT4 mult_10_i327_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n486_adj_3621));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4456_3_lut (.I0(GND_net), .I1(n8961[0]), .I2(n222_adj_3526), 
            .I3(n36427), .O(n8937[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_8_lut (.I0(\PID_CONTROLLER.result[6] ), .I1(n49785), 
            .I2(n61[6]), .I3(n34725), .O(n1_adj_3674)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_8 (.CI(n34725), .I0(n49785), .I1(n61[6]), 
            .CO(n34726));
    SB_CARRY add_4788_2 (.CI(GND_net), .I0(n72), .I1(n107), .CO(n36664));
    SB_CARRY add_4456_3 (.CI(n36427), .I0(n8961[0]), .I1(n222_adj_3526), 
            .CO(n36428));
    SB_LUT4 add_28678_27_lut (.I0(GND_net), .I1(n66[25]), .I2(n191[25]), 
            .I3(n34892), .O(\PID_CONTROLLER.result_31__N_3353 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_7_lut (.I0(\PID_CONTROLLER.result [5]), .I1(n49785), 
            .I2(n61[5]), .I3(n34724), .O(n466)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_4446_7_lut (.I0(GND_net), .I1(n8700[4]), .I2(n652), .I3(n36085), 
            .O(n8690[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_7 (.CI(n36085), .I0(n8700[4]), .I1(n652), .CO(n36086));
    SB_LUT4 add_4472_23_lut (.I0(GND_net), .I1(n9225[20]), .I2(GND_net), 
            .I3(n36663), .O(n9201[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i392_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3620));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4446_6_lut (.I0(GND_net), .I1(n8700[3]), .I2(n555), .I3(n36084), 
            .O(n8690[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_24_lut (.I0(GND_net), .I1(n1804[21]), .I2(GND_net), 
            .I3(n36909), .O(n1803[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n680_adj_3618));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_28678_27 (.CI(n34892), .I0(n66[25]), .I1(n191[25]), .CO(n34893));
    SB_LUT4 mult_14_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4456_2_lut (.I0(GND_net), .I1(n32_adj_3523), .I2(n125_adj_3521), 
            .I3(GND_net), .O(n8937[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4456_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_15_lut (.I0(GND_net), .I1(n1800[12]), .I2(GND_net), 
            .I3(n36808), .O(n1799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_6 (.CI(n36084), .I0(n8700[3]), .I1(n555), .CO(n36085));
    SB_CARRY unary_minus_23_add_3_7 (.CI(n34724), .I0(n49785), .I1(n61[5]), 
            .CO(n34725));
    SB_LUT4 add_4446_5_lut (.I0(GND_net), .I1(n8700[2]), .I2(n458_adj_3519), 
            .I3(n36083), .O(n8690[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_22_lut (.I0(GND_net), .I1(n9225[19]), .I2(GND_net), 
            .I3(n36662), .O(n9201[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_6_lut (.I0(\PID_CONTROLLER.result[4] ), .I1(n49785), 
            .I2(n61[4]), .I3(n34723), .O(n1_adj_3675)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4456_2 (.CI(GND_net), .I0(n32_adj_3523), .I1(n125_adj_3521), 
            .CO(n36427));
    SB_CARRY mult_14_add_1214_15 (.CI(n36808), .I0(n1800[12]), .I1(GND_net), 
            .CO(n36809));
    SB_LUT4 mult_12_i89_2_lut (.I0(\Kd[1] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_3617));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i89_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4446_5 (.CI(n36083), .I0(n8700[2]), .I1(n458_adj_3519), 
            .CO(n36084));
    SB_LUT4 add_4455_24_lut (.I0(GND_net), .I1(n8937[21]), .I2(GND_net), 
            .I3(n36426), .O(n8912[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_4_lut (.I0(GND_net), .I1(n8700[1]), .I2(n361), .I3(n36082), 
            .O(n8690[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_4 (.CI(n36082), .I0(n8700[1]), .I1(n361), .CO(n36083));
    SB_CARRY add_4472_22 (.CI(n36662), .I0(n9225[19]), .I1(GND_net), .CO(n36663));
    SB_LUT4 add_4455_23_lut (.I0(GND_net), .I1(n8937[20]), .I2(GND_net), 
            .I3(n36425), .O(n8912[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_23 (.CI(n36425), .I0(n8937[20]), .I1(GND_net), .CO(n36426));
    SB_LUT4 add_4446_3_lut (.I0(GND_net), .I1(n8700[0]), .I2(n264), .I3(n36081), 
            .O(n8690[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i26_2_lut (.I0(\Kd[0] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4455_22_lut (.I0(GND_net), .I1(n8937[19]), .I2(GND_net), 
            .I3(n36424), .O(n8912[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_3 (.CI(n36081), .I0(n8700[0]), .I1(n264), .CO(n36082));
    SB_LUT4 add_4446_2_lut (.I0(GND_net), .I1(n80), .I2(n167), .I3(GND_net), 
            .O(n8690[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[22]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4446_2 (.CI(GND_net), .I0(n80), .I1(n167), .CO(n36081));
    SB_CARRY add_4455_22 (.CI(n36424), .I0(n8937[19]), .I1(GND_net), .CO(n36425));
    SB_LUT4 LessThan_22_i41_2_lut (.I0(\PID_CONTROLLER.result [20]), .I1(n67[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3676));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4445_10_lut (.I0(GND_net), .I1(n8690[7]), .I2(GND_net), 
            .I3(n36080), .O(n8679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_26_lut (.I0(GND_net), .I1(n66[24]), .I2(n191[24]), 
            .I3(n34891), .O(\PID_CONTROLLER.result_31__N_3353 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_6 (.CI(n34723), .I0(n49785), .I1(n61[4]), 
            .CO(n34724));
    SB_LUT4 LessThan_22_i45_2_lut (.I0(\PID_CONTROLLER.result [22]), .I1(n67[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_3678));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i43_2_lut (.I0(\PID_CONTROLLER.result [21]), .I1(n67[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_3680));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4445_9_lut (.I0(GND_net), .I1(n8690[6]), .I2(GND_net), 
            .I3(n36079), .O(n8679[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4445_9 (.CI(n36079), .I0(n8690[6]), .I1(GND_net), .CO(n36080));
    SB_LUT4 add_4472_21_lut (.I0(GND_net), .I1(n9225[18]), .I2(GND_net), 
            .I3(n36661), .O(n9201[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_21_lut (.I0(GND_net), .I1(n8937[18]), .I2(GND_net), 
            .I3(n36423), .O(n8912[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4445_8_lut (.I0(GND_net), .I1(n8690[5]), .I2(n746), .I3(n36078), 
            .O(n8679[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4445_8 (.CI(n36078), .I0(n8690[5]), .I1(n746), .CO(n36079));
    SB_LUT4 add_4445_7_lut (.I0(GND_net), .I1(n8690[4]), .I2(n649), .I3(n36077), 
            .O(n8679[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_5_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n49785), 
            .I2(n61[3]), .I3(n34722), .O(n468)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4445_7 (.CI(n36077), .I0(n8690[4]), .I1(n649), .CO(n36078));
    SB_CARRY add_4455_21 (.CI(n36423), .I0(n8937[18]), .I1(GND_net), .CO(n36424));
    SB_CARRY unary_minus_23_add_3_5 (.CI(n34722), .I0(n49785), .I1(n61[3]), 
            .CO(n34723));
    SB_LUT4 add_13_add_1_28678_add_1_33_lut (.I0(GND_net), .I1(n6821[8]), 
            .I2(n6807[0]), .I3(n36991), .O(n66[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_21 (.CI(n36661), .I0(n9225[18]), .I1(GND_net), .CO(n36662));
    SB_LUT4 mult_14_add_1214_14_lut (.I0(GND_net), .I1(n1800[11]), .I2(GND_net), 
            .I3(n36807), .O(n1799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i37_2_lut (.I0(\PID_CONTROLLER.result [18]), .I1(n67[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3681));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_14_add_1218_24 (.CI(n36909), .I0(n1804[21]), .I1(GND_net), 
            .CO(n1711));
    SB_CARRY mult_14_add_1214_14 (.CI(n36807), .I0(n1800[11]), .I1(GND_net), 
            .CO(n36808));
    SB_LUT4 add_4472_20_lut (.I0(GND_net), .I1(n9225[17]), .I2(GND_net), 
            .I3(n36660), .O(n9201[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_20 (.CI(n36660), .I0(n9225[17]), .I1(GND_net), .CO(n36661));
    SB_LUT4 add_4472_19_lut (.I0(GND_net), .I1(n9225[16]), .I2(GND_net), 
            .I3(n36659), .O(n9201[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_20_lut (.I0(GND_net), .I1(n8937[17]), .I2(GND_net), 
            .I3(n36422), .O(n8912[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_20 (.CI(n36422), .I0(n8937[17]), .I1(GND_net), .CO(n36423));
    SB_LUT4 add_4455_19_lut (.I0(GND_net), .I1(n8937[16]), .I2(GND_net), 
            .I3(n36421), .O(n8912[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4445_6_lut (.I0(GND_net), .I1(n8690[3]), .I2(n552), .I3(n36076), 
            .O(n8679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4445_6 (.CI(n36076), .I0(n8690[3]), .I1(n552), .CO(n36077));
    SB_LUT4 add_4445_5_lut (.I0(GND_net), .I1(n8690[2]), .I2(n455_adj_3509), 
            .I3(n36075), .O(n8679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_19 (.CI(n36421), .I0(n8937[16]), .I1(GND_net), .CO(n36422));
    SB_CARRY add_28678_26 (.CI(n34891), .I0(n66[24]), .I1(n191[24]), .CO(n34892));
    SB_LUT4 LessThan_22_i29_2_lut (.I0(\PID_CONTROLLER.result [14]), .I1(n67[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3682));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i31_2_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n67[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_3683));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4445_5 (.CI(n36075), .I0(n8690[2]), .I1(n455_adj_3509), 
            .CO(n36076));
    SB_LUT4 add_13_add_1_28678_add_1_32_lut (.I0(GND_net), .I1(n6821[7]), 
            .I2(n64[30]), .I3(n36990), .O(n66[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4445_4_lut (.I0(GND_net), .I1(n8690[1]), .I2(n358), .I3(n36074), 
            .O(n8679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4445_4 (.CI(n36074), .I0(n8690[1]), .I1(n358), .CO(n36075));
    SB_LUT4 add_4445_3_lut (.I0(GND_net), .I1(n8690[0]), .I2(n261), .I3(n36073), 
            .O(n8679[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_19 (.CI(n36659), .I0(n9225[16]), .I1(GND_net), .CO(n36660));
    SB_LUT4 LessThan_22_i23_2_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n67[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3684));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_28678_25_lut (.I0(GND_net), .I1(n66[23]), .I2(n191[23]), 
            .I3(n34890), .O(\PID_CONTROLLER.result_31__N_3353 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_18_lut (.I0(GND_net), .I1(n9225[15]), .I2(GND_net), 
            .I3(n36658), .O(n9201[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_18_lut (.I0(GND_net), .I1(n8937[15]), .I2(GND_net), 
            .I3(n36420), .O(n8912[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_4_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n49785), 
            .I2(n61[2]), .I3(n34721), .O(n469)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_28678_25 (.CI(n34890), .I0(n66[23]), .I1(n191[23]), .CO(n34891));
    SB_CARRY add_4445_3 (.CI(n36073), .I0(n8690[0]), .I1(n261), .CO(n36074));
    SB_CARRY add_4472_18 (.CI(n36658), .I0(n9225[15]), .I1(GND_net), .CO(n36659));
    SB_LUT4 add_28678_24_lut (.I0(GND_net), .I1(n66[22]), .I2(n191[22]), 
            .I3(n34889), .O(\PID_CONTROLLER.result_31__N_3353 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_4 (.CI(n34721), .I0(n49785), .I1(n61[2]), 
            .CO(n34722));
    SB_LUT4 add_4445_2_lut (.I0(GND_net), .I1(n71), .I2(n164), .I3(GND_net), 
            .O(n8679[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4445_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4445_2 (.CI(GND_net), .I0(n71), .I1(n164), .CO(n36073));
    SB_LUT4 sub_11_add_2_27_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n60[26]), .I3(n34624), .O(n58[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_18 (.CI(n36420), .I0(n8937[15]), .I1(GND_net), .CO(n36421));
    SB_LUT4 sub_11_add_2_26_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n60[26]), .I3(n34623), .O(n58[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_13_lut (.I0(GND_net), .I1(n1800[10]), .I2(GND_net), 
            .I3(n36806), .O(n1799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_17_lut (.I0(GND_net), .I1(n9225[14]), .I2(GND_net), 
            .I3(n36657), .O(n9201[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_17_lut (.I0(GND_net), .I1(n8937[14]), .I2(GND_net), 
            .I3(n36419), .O(n8912[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_11_lut (.I0(GND_net), .I1(n8679[8]), .I2(GND_net), 
            .I3(n36072), .O(n8667[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_10_lut (.I0(GND_net), .I1(n8679[7]), .I2(GND_net), 
            .I3(n36071), .O(n8667[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_17 (.CI(n36419), .I0(n8937[14]), .I1(GND_net), .CO(n36420));
    SB_CARRY add_4444_10 (.CI(n36071), .I0(n8679[7]), .I1(GND_net), .CO(n36072));
    SB_LUT4 add_4444_9_lut (.I0(GND_net), .I1(n8679[6]), .I2(GND_net), 
            .I3(n36070), .O(n8667[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_17 (.CI(n36657), .I0(n9225[14]), .I1(GND_net), .CO(n36658));
    SB_LUT4 add_4455_16_lut (.I0(GND_net), .I1(n8937[13]), .I2(GND_net), 
            .I3(n36418), .O(n8912[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_9 (.CI(n36070), .I0(n8679[6]), .I1(GND_net), .CO(n36071));
    SB_LUT4 add_4444_8_lut (.I0(GND_net), .I1(n8679[5]), .I2(n743), .I3(n36069), 
            .O(n8667[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i25_2_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n67[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3686));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_23_add_3_3_lut (.I0(\PID_CONTROLLER.result [1]), .I1(n49785), 
            .I2(n61[1]), .I3(n34720), .O(n470)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_4455_16 (.CI(n36418), .I0(n8937[13]), .I1(GND_net), .CO(n36419));
    SB_LUT4 add_4455_15_lut (.I0(GND_net), .I1(n8937[12]), .I2(GND_net), 
            .I3(n36417), .O(n8912[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_8 (.CI(n36069), .I0(n8679[5]), .I1(n743), .CO(n36070));
    SB_LUT4 mult_14_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_28678_add_1_32 (.CI(n36990), .I0(n6821[7]), .I1(n64[30]), 
            .CO(n36991));
    SB_LUT4 add_13_add_1_28678_add_1_31_lut (.I0(GND_net), .I1(n6821[6]), 
            .I2(n64[29]), .I3(n36989), .O(n66[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_31 (.CI(n36989), .I0(n6821[6]), .I1(n64[29]), 
            .CO(n36990));
    SB_LUT4 mult_14_add_1218_23_lut (.I0(GND_net), .I1(n1804[20]), .I2(GND_net), 
            .I3(n36908), .O(n1803[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_13 (.CI(n36806), .I0(n1800[10]), .I1(GND_net), 
            .CO(n36807));
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[4]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4444_7_lut (.I0(GND_net), .I1(n8679[4]), .I2(n646), .I3(n36068), 
            .O(n8667[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_24 (.CI(n34889), .I0(n66[22]), .I1(n191[22]), .CO(n34890));
    SB_CARRY add_4444_7 (.CI(n36068), .I0(n8679[4]), .I1(n646), .CO(n36069));
    SB_LUT4 add_28678_23_lut (.I0(GND_net), .I1(n66[21]), .I2(n191[21]), 
            .I3(n34888), .O(\PID_CONTROLLER.result_31__N_3353 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_3 (.CI(n34720), .I0(n49785), .I1(n61[1]), 
            .CO(n34721));
    SB_CARRY add_4455_15 (.CI(n36417), .I0(n8937[12]), .I1(GND_net), .CO(n36418));
    SB_LUT4 add_4472_16_lut (.I0(GND_net), .I1(n9225[13]), .I2(GND_net), 
            .I3(n36656), .O(n9201[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_26 (.CI(n34623), .I0(\PID_CONTROLLER.err_prev[31] ), 
            .I1(n60[26]), .CO(n34624));
    SB_LUT4 add_4444_6_lut (.I0(GND_net), .I1(n8679[3]), .I2(n549), .I3(n36067), 
            .O(n8667[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_2_lut (.I0(\PID_CONTROLLER.result [0]), .I1(n49785), 
            .I2(n61[0]), .I3(VCC_net), .O(n471)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_22_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n67[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3688));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_11_add_2_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[23] ), 
            .I2(n60[23]), .I3(n34622), .O(n58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_23 (.CI(n34888), .I0(n66[21]), .I1(n191[21]), .CO(n34889));
    SB_LUT4 add_4455_14_lut (.I0(GND_net), .I1(n8937[11]), .I2(GND_net), 
            .I3(n36416), .O(n8912[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_6 (.CI(n36067), .I0(n8679[3]), .I1(n549), .CO(n36068));
    SB_LUT4 mult_14_add_1214_12_lut (.I0(GND_net), .I1(n1800[9]), .I2(GND_net), 
            .I3(n36805), .O(n1799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_14 (.CI(n36416), .I0(n8937[11]), .I1(GND_net), .CO(n36417));
    SB_LUT4 LessThan_22_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n67[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3690));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_28678_22_lut (.I0(GND_net), .I1(n66[20]), .I2(n191[20]), 
            .I3(n34887), .O(\PID_CONTROLLER.result_31__N_3353 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_5_lut (.I0(GND_net), .I1(n8679[2]), .I2(n452), .I3(n36066), 
            .O(n8667[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_13_lut (.I0(GND_net), .I1(n8937[10]), .I2(GND_net), 
            .I3(n36415), .O(n8912[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_25 (.CI(n34622), .I0(\PID_CONTROLLER.err_prev[23] ), 
            .I1(n60[23]), .CO(n34623));
    SB_CARRY mult_14_add_1214_12 (.CI(n36805), .I0(n1800[9]), .I1(GND_net), 
            .CO(n36806));
    SB_CARRY add_4444_5 (.CI(n36066), .I0(n8679[2]), .I1(n452), .CO(n36067));
    SB_LUT4 add_13_add_1_28678_add_1_30_lut (.I0(GND_net), .I1(n6821[5]), 
            .I2(n64[28]), .I3(n36988), .O(n66[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_30 (.CI(n36988), .I0(n6821[5]), .I1(n64[28]), 
            .CO(n36989));
    SB_LUT4 add_4444_4_lut (.I0(GND_net), .I1(n8679[1]), .I2(n355), .I3(n36065), 
            .O(n8667[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_23 (.CI(n36908), .I0(n1804[20]), .I1(GND_net), 
            .CO(n36909));
    SB_CARRY add_4444_4 (.CI(n36065), .I0(n8679[1]), .I1(n355), .CO(n36066));
    SB_CARRY add_4455_13 (.CI(n36415), .I0(n8937[10]), .I1(GND_net), .CO(n36416));
    SB_CARRY add_28678_22 (.CI(n34887), .I0(n66[20]), .I1(n191[20]), .CO(n34888));
    SB_CARRY add_4472_16 (.CI(n36656), .I0(n9225[13]), .I1(GND_net), .CO(n36657));
    SB_LUT4 add_4455_12_lut (.I0(GND_net), .I1(n8937[9]), .I2(GND_net), 
            .I3(n36414), .O(n8912[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4444_3_lut (.I0(GND_net), .I1(n8679[0]), .I2(n258), .I3(n36064), 
            .O(n8667[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_12 (.CI(n36414), .I0(n8937[9]), .I1(GND_net), .CO(n36415));
    SB_LUT4 add_4472_15_lut (.I0(GND_net), .I1(n9225[12]), .I2(GND_net), 
            .I3(n36655), .O(n9201[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_11_lut (.I0(GND_net), .I1(n8937[8]), .I2(GND_net), 
            .I3(n36413), .O(n8912[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i33_2_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n67[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_3692));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i11_2_lut (.I0(\PID_CONTROLLER.result [5]), .I1(n67[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3693));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4455_11 (.CI(n36413), .I0(n8937[8]), .I1(GND_net), .CO(n36414));
    SB_LUT4 add_28678_21_lut (.I0(GND_net), .I1(n66[19]), .I2(n191[19]), 
            .I3(n34886), .O(\PID_CONTROLLER.result_31__N_3353 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_29_lut (.I0(GND_net), .I1(n6821[4]), 
            .I2(n64[27]), .I3(n36987), .O(n66[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_2 (.CI(VCC_net), .I0(n49785), .I1(n61[0]), 
            .CO(n34720));
    SB_LUT4 mult_14_add_1218_22_lut (.I0(GND_net), .I1(n1804[19]), .I2(GND_net), 
            .I3(n36907), .O(n1803[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_15 (.CI(n36655), .I0(n9225[12]), .I1(GND_net), .CO(n36656));
    SB_LUT4 add_4472_14_lut (.I0(GND_net), .I1(n9225[11]), .I2(GND_net), 
            .I3(n36654), .O(n9201[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_29 (.CI(n36987), .I0(n6821[4]), .I1(n64[27]), 
            .CO(n36988));
    SB_LUT4 LessThan_22_i15_2_lut (.I0(\PID_CONTROLLER.result [7]), .I1(n67[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3695));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_add_1214_11_lut (.I0(GND_net), .I1(n1800[8]), .I2(GND_net), 
            .I3(n36804), .O(n1799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_22 (.CI(n36907), .I0(n1804[19]), .I1(GND_net), 
            .CO(n36908));
    SB_LUT4 add_4455_10_lut (.I0(GND_net), .I1(n8937[7]), .I2(GND_net), 
            .I3(n36412), .O(n8912[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_21 (.CI(n34886), .I0(n66[19]), .I1(n191[19]), .CO(n34887));
    SB_CARRY add_4472_14 (.CI(n36654), .I0(n9225[11]), .I1(GND_net), .CO(n36655));
    SB_CARRY add_4444_3 (.CI(n36064), .I0(n8679[0]), .I1(n258), .CO(n36065));
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(n61[31]), 
            .I3(n34719), .O(n67[24])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_10 (.CI(n36412), .I0(n8937[7]), .I1(GND_net), .CO(n36413));
    SB_LUT4 add_4444_2_lut (.I0(GND_net), .I1(n68), .I2(n161), .I3(GND_net), 
            .O(n8667[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4444_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4444_2 (.CI(GND_net), .I0(n68), .I1(n161), .CO(n36064));
    SB_LUT4 add_28678_20_lut (.I0(GND_net), .I1(n66[18]), .I2(n191[18]), 
            .I3(n34885), .O(\PID_CONTROLLER.result_31__N_3353 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_28_lut (.I0(GND_net), .I1(n6821[3]), 
            .I2(n64[26]), .I3(n36986), .O(n66[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i32_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[31]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39199_4_lut (.I0(n27_adj_5), .I1(n15_adj_3695), .I2(n13_adj_6), 
            .I3(n11_adj_3693), .O(n47101));
    defparam i39199_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_14_add_1214_11 (.CI(n36804), .I0(n1800[8]), .I1(GND_net), 
            .CO(n36805));
    SB_CARRY add_13_add_1_28678_add_1_28 (.CI(n36986), .I0(n6821[3]), .I1(n64[26]), 
            .CO(n36987));
    SB_LUT4 add_4455_9_lut (.I0(GND_net), .I1(n8937[6]), .I2(GND_net), 
            .I3(n36411), .O(n8912[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4443_12_lut (.I0(GND_net), .I1(n8667[9]), .I2(GND_net), 
            .I3(n36063), .O(n8654[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_21_lut (.I0(GND_net), .I1(n1804[18]), .I2(GND_net), 
            .I3(n36906), .O(n1803[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4443_11_lut (.I0(GND_net), .I1(n8667[8]), .I2(GND_net), 
            .I3(n36062), .O(n8654[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i12_3_lut (.I0(n67[7]), .I1(n67[16]), .I2(n33_adj_3692), 
            .I3(GND_net), .O(n12_adj_3698));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_11_add_2_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[22] ), 
            .I2(n60[22]), .I3(n34621), .O(n58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_20 (.CI(n34885), .I0(n66[18]), .I1(n191[18]), .CO(n34886));
    SB_CARRY sub_11_add_2_24 (.CI(n34621), .I0(\PID_CONTROLLER.err_prev[22] ), 
            .I1(n60[22]), .CO(n34622));
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n61[31]), 
            .I3(n34718), .O(n67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_9 (.CI(n36411), .I0(n8937[6]), .I1(GND_net), .CO(n36412));
    SB_LUT4 add_28678_19_lut (.I0(GND_net), .I1(n66[17]), .I2(n191[17]), 
            .I3(n34884), .O(\PID_CONTROLLER.result_31__N_3353 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[21] ), 
            .I2(n60[21]), .I3(n34620), .O(n58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n34718), .I0(GND_net), .I1(n61[31]), 
            .CO(n34719));
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n61[22]), 
            .I3(n34717), .O(n67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_11 (.CI(n36062), .I0(n8667[8]), .I1(GND_net), .CO(n36063));
    SB_CARRY mult_14_add_1218_21 (.CI(n36906), .I0(n1804[18]), .I1(GND_net), 
            .CO(n36907));
    SB_CARRY add_28678_19 (.CI(n34884), .I0(n66[17]), .I1(n191[17]), .CO(n34885));
    SB_LUT4 LessThan_22_i10_3_lut (.I0(n67[5]), .I1(n414), .I2(n13_adj_6), 
            .I3(GND_net), .O(n10_adj_3701));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i30_3_lut (.I0(n12_adj_3698), .I1(n403), .I2(n35_adj_7), 
            .I3(GND_net), .O(n30_adj_3703));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_add_1218_20_lut (.I0(GND_net), .I1(n1804[17]), .I2(GND_net), 
            .I3(n36905), .O(n1803[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_8_lut (.I0(GND_net), .I1(n8937[5]), .I2(n704_adj_3704), 
            .I3(n36410), .O(n8912[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1190__i0 (.Q(Kd_delay_counter[0]), .C(clk32MHz), 
           .D(n69[0]));   // verilog/motorControl.v(55[27:47])
    SB_LUT4 mult_14_add_1214_10_lut (.I0(GND_net), .I1(n1800[7]), .I2(GND_net), 
            .I3(n36803), .O(n1799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_20 (.CI(n36905), .I0(n1804[17]), .I1(GND_net), 
            .CO(n36906));
    SB_LUT4 add_4443_10_lut (.I0(GND_net), .I1(n8667[7]), .I2(GND_net), 
            .I3(n36061), .O(n8654[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_24 (.CI(n34717), .I0(GND_net), .I1(n61[22]), 
            .CO(n34718));
    SB_LUT4 add_13_add_1_28678_add_1_27_lut (.I0(GND_net), .I1(n6821[2]), 
            .I2(n64[25]), .I3(n36985), .O(n66[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_10 (.CI(n36061), .I0(n8667[7]), .I1(GND_net), .CO(n36062));
    SB_CARRY mult_14_add_1214_10 (.CI(n36803), .I0(n1800[7]), .I1(GND_net), 
            .CO(n36804));
    SB_LUT4 add_4443_9_lut (.I0(GND_net), .I1(n8667[6]), .I2(GND_net), 
            .I3(n36060), .O(n8654[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_9 (.CI(n36060), .I0(n8667[6]), .I1(GND_net), .CO(n36061));
    SB_LUT4 add_4472_13_lut (.I0(GND_net), .I1(n9225[10]), .I2(GND_net), 
            .I3(n36653), .O(n9201[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_19_lut (.I0(GND_net), .I1(n1804[16]), .I2(GND_net), 
            .I3(n36904), .O(n1803[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_18_lut (.I0(GND_net), .I1(n66[16]), .I2(n191[16]), 
            .I3(n34883), .O(\PID_CONTROLLER.result_31__N_3353 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_9_lut (.I0(GND_net), .I1(n1800[6]), .I2(GND_net), 
            .I3(n36802), .O(n1799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_13 (.CI(n36653), .I0(n9225[10]), .I1(GND_net), .CO(n36654));
    SB_CARRY add_4455_8 (.CI(n36410), .I0(n8937[5]), .I1(n704_adj_3704), 
            .CO(n36411));
    SB_LUT4 add_4443_8_lut (.I0(GND_net), .I1(n8667[5]), .I2(n740), .I3(n36059), 
            .O(n8654[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_12_lut (.I0(GND_net), .I1(n9225[9]), .I2(GND_net), 
            .I3(n36652), .O(n9201[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39999_4_lut (.I0(n13_adj_6), .I1(n11_adj_3693), .I2(n9_adj_8), 
            .I3(n47118), .O(n47902));
    defparam i39999_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_4443_8 (.CI(n36059), .I0(n8667[5]), .I1(n740), .CO(n36060));
    SB_LUT4 i39995_4_lut (.I0(n19_adj_3690), .I1(n17_adj_3688), .I2(n15_adj_3695), 
            .I3(n47902), .O(n47898));
    defparam i39995_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_4443_7_lut (.I0(GND_net), .I1(n8667[4]), .I2(n643), .I3(n36058), 
            .O(n8654[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n61[21]), 
            .I3(n34716), .O(n67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_18 (.CI(n34883), .I0(n66[16]), .I1(n191[16]), .CO(n34884));
    SB_LUT4 i40886_4_lut (.I0(n25_adj_3686), .I1(n23_adj_3684), .I2(n21_adj_9), 
            .I3(n47898), .O(n48789));
    defparam i40886_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4455_7_lut (.I0(GND_net), .I1(n8937[4]), .I2(n607_adj_3708), 
            .I3(n36409), .O(n8912[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_23 (.CI(n34620), .I0(\PID_CONTROLLER.err_prev[21] ), 
            .I1(n60[21]), .CO(n34621));
    SB_CARRY add_4443_7 (.CI(n36058), .I0(n8667[4]), .I1(n643), .CO(n36059));
    SB_LUT4 sub_11_add_2_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[20] ), 
            .I2(n60[20]), .I3(n34619), .O(n58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_27 (.CI(n36985), .I0(n6821[2]), .I1(n64[25]), 
            .CO(n36986));
    SB_CARRY add_4455_7 (.CI(n36409), .I0(n8937[4]), .I1(n607_adj_3708), 
            .CO(n36410));
    SB_LUT4 add_4443_6_lut (.I0(GND_net), .I1(n8667[3]), .I2(n546), .I3(n36057), 
            .O(n8654[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_9 (.CI(n36802), .I0(n1800[6]), .I1(GND_net), 
            .CO(n36803));
    SB_CARRY add_4472_12 (.CI(n36652), .I0(n9225[9]), .I1(GND_net), .CO(n36653));
    SB_LUT4 i40364_4_lut (.I0(n31_adj_3683), .I1(n29_adj_3682), .I2(n27_adj_5), 
            .I3(n48789), .O(n48267));
    defparam i40364_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_4472_11_lut (.I0(GND_net), .I1(n9225[8]), .I2(GND_net), 
            .I3(n36651), .O(n9201[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_17_lut (.I0(GND_net), .I1(n66[15]), .I2(n191[15]), 
            .I3(n34882), .O(\PID_CONTROLLER.result_31__N_3353 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_11 (.CI(n36651), .I0(n9225[8]), .I1(GND_net), .CO(n36652));
    SB_LUT4 add_4472_10_lut (.I0(GND_net), .I1(n9225[7]), .I2(GND_net), 
            .I3(n36650), .O(n9201[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_6_lut (.I0(GND_net), .I1(n8937[3]), .I2(n510_adj_3710), 
            .I3(n36408), .O(n8912[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_17 (.CI(n34882), .I0(n66[15]), .I1(n191[15]), .CO(n34883));
    SB_LUT4 add_13_add_1_28678_add_1_26_lut (.I0(GND_net), .I1(n6821[1]), 
            .I2(n64[24]), .I3(n36984), .O(n66[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_19 (.CI(n36904), .I0(n1804[16]), .I1(GND_net), 
            .CO(n36905));
    SB_LUT4 mult_14_add_1214_8_lut (.I0(GND_net), .I1(n1800[5]), .I2(n521), 
            .I3(n36801), .O(n1799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41009_4_lut (.I0(n37_adj_3681), .I1(n35_adj_7), .I2(n33_adj_3692), 
            .I3(n48267), .O(n48912));
    defparam i41009_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_4472_10 (.CI(n36650), .I0(n9225[7]), .I1(GND_net), .CO(n36651));
    SB_CARRY unary_minus_21_add_3_23 (.CI(n34716), .I0(GND_net), .I1(n61[21]), 
            .CO(n34717));
    SB_CARRY add_4455_6 (.CI(n36408), .I0(n8937[3]), .I1(n510_adj_3710), 
            .CO(n36409));
    SB_LUT4 add_4455_5_lut (.I0(GND_net), .I1(n8937[2]), .I2(n413_adj_3712), 
            .I3(n36407), .O(n8912[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n61[20]), 
            .I3(n34715), .O(n67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_26 (.CI(n36984), .I0(n6821[1]), .I1(n64[24]), 
            .CO(n36985));
    SB_CARRY add_4443_6 (.CI(n36057), .I0(n8667[3]), .I1(n546), .CO(n36058));
    SB_CARRY mult_14_add_1214_8 (.CI(n36801), .I0(n1800[5]), .I1(n521), 
            .CO(n36802));
    SB_LUT4 add_4443_5_lut (.I0(GND_net), .I1(n8667[2]), .I2(n449_adj_3713), 
            .I3(n36056), .O(n8654[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_9_lut (.I0(GND_net), .I1(n9225[6]), .I2(GND_net), 
            .I3(n36649), .O(n9201[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4455_5 (.CI(n36407), .I0(n8937[2]), .I1(n413_adj_3712), 
            .CO(n36408));
    SB_CARRY add_4443_5 (.CI(n36056), .I0(n8667[2]), .I1(n449_adj_3713), 
            .CO(n36057));
    SB_LUT4 add_4443_4_lut (.I0(GND_net), .I1(n8667[1]), .I2(n352), .I3(n36055), 
            .O(n8654[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_4_lut (.I0(GND_net), .I1(n8937[1]), .I2(n316_adj_3714), 
            .I3(n36406), .O(n8912[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_4 (.CI(n36055), .I0(n8667[1]), .I1(n352), .CO(n36056));
    SB_LUT4 i40508_3_lut (.I0(n6_adj_3715), .I1(n410), .I2(n21_adj_9), 
            .I3(GND_net), .O(n48411));   // verilog/motorControl.v(47[21:37])
    defparam i40508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40509_3_lut (.I0(n48411), .I1(n67[11]), .I2(n23_adj_3684), 
            .I3(GND_net), .O(n48412));   // verilog/motorControl.v(47[21:37])
    defparam i40509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4443_3_lut (.I0(GND_net), .I1(n8667[0]), .I2(n255), .I3(n36054), 
            .O(n8654[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_9 (.CI(n36649), .I0(n9225[6]), .I1(GND_net), .CO(n36650));
    SB_LUT4 LessThan_22_i16_3_lut (.I0(n67[9]), .I1(n67[21]), .I2(n43_adj_3680), 
            .I3(GND_net), .O(n16_adj_3717));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4455_4 (.CI(n36406), .I0(n8937[1]), .I1(n316_adj_3714), 
            .CO(n36407));
    SB_CARRY add_4443_3 (.CI(n36054), .I0(n8667[0]), .I1(n255), .CO(n36055));
    SB_LUT4 add_4443_2_lut (.I0(GND_net), .I1(n65), .I2(n158), .I3(GND_net), 
            .O(n8654[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4443_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4443_2 (.CI(GND_net), .I0(n65), .I1(n158), .CO(n36054));
    SB_LUT4 add_4455_3_lut (.I0(GND_net), .I1(n8937[0]), .I2(n219_adj_3718), 
            .I3(n36405), .O(n8912[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_13_lut (.I0(GND_net), .I1(n8654[10]), .I2(GND_net), 
            .I3(n36053), .O(n8640[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_12_lut (.I0(GND_net), .I1(n8654[9]), .I2(GND_net), 
            .I3(n36052), .O(n8640[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i8_3_lut (.I0(n416), .I1(n67[8]), .I2(n17_adj_3688), 
            .I3(GND_net), .O(n8_adj_3720));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4455_3 (.CI(n36405), .I0(n8937[0]), .I1(n219_adj_3718), 
            .CO(n36406));
    SB_CARRY add_4442_12 (.CI(n36052), .I0(n8654[9]), .I1(GND_net), .CO(n36053));
    SB_LUT4 add_4442_11_lut (.I0(GND_net), .I1(n8654[8]), .I2(GND_net), 
            .I3(n36051), .O(n8640[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_16_lut (.I0(GND_net), .I1(n66[14]), .I2(n191[14]), 
            .I3(n34881), .O(\PID_CONTROLLER.result_31__N_3353 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i24_3_lut (.I0(n16_adj_3717), .I1(n67[22]), .I2(n45_adj_3678), 
            .I3(GND_net), .O(n24_adj_3721));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39205_4_lut (.I0(n21_adj_9), .I1(n19_adj_3690), .I2(n17_adj_3688), 
            .I3(n9_adj_8), .O(n47107));
    defparam i39205_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4442_11 (.CI(n36051), .I0(n8654[8]), .I1(GND_net), .CO(n36052));
    SB_LUT4 i39185_4_lut (.I0(n43_adj_3680), .I1(n25_adj_3686), .I2(n23_adj_3684), 
            .I3(n47107), .O(n47087));
    defparam i39185_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n34715), .I0(GND_net), .I1(n61[20]), 
            .CO(n34716));
    SB_LUT4 i41025_4_lut (.I0(n24_adj_3721), .I1(n8_adj_3720), .I2(n45_adj_3678), 
            .I3(n47085), .O(n48928));   // verilog/motorControl.v(47[21:37])
    defparam i41025_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_13_add_1_28678_add_1_25_lut (.I0(GND_net), .I1(n6821[0]), 
            .I2(n64[23]), .I3(n36983), .O(n66[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n61[19]), 
            .I3(n34714), .O(n401)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_16 (.CI(n34881), .I0(n66[14]), .I1(n191[14]), .CO(n34882));
    SB_LUT4 i39825_3_lut (.I0(n48412), .I1(n67[12]), .I2(n25_adj_3686), 
            .I3(GND_net), .O(n47728));   // verilog/motorControl.v(47[21:37])
    defparam i39825_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_11_add_2_22 (.CI(n34619), .I0(\PID_CONTROLLER.err_prev[20] ), 
            .I1(n60[20]), .CO(n34620));
    SB_LUT4 i3_3_lut (.I0(\PID_CONTROLLER.result [30]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(n67[24]), .I3(GND_net), .O(n10_adj_3723));   // verilog/motorControl.v(47[21:37])
    defparam i3_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 add_4442_10_lut (.I0(GND_net), .I1(n8654[7]), .I2(GND_net), 
            .I3(n36050), .O(n8640[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4455_2_lut (.I0(GND_net), .I1(n29_adj_3724), .I2(n122_adj_3725), 
            .I3(GND_net), .O(n8912[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4455_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_8_lut (.I0(GND_net), .I1(n9225[5]), .I2(n545), .I3(n36648), 
            .O(n9201[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_8 (.CI(n36648), .I0(n9225[5]), .I1(n545), .CO(n36649));
    SB_LUT4 sub_11_add_2_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[19] ), 
            .I2(n60[19]), .I3(n34618), .O(n58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_10 (.CI(n36050), .I0(n8654[7]), .I1(GND_net), .CO(n36051));
    SB_CARRY unary_minus_21_add_3_21 (.CI(n34714), .I0(GND_net), .I1(n61[19]), 
            .CO(n34715));
    SB_LUT4 i1_3_lut (.I0(\PID_CONTROLLER.result [26]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(n67[24]), .I3(GND_net), .O(n8_adj_3728));   // verilog/motorControl.v(47[21:37])
    defparam i1_3_lut.LUT_INIT = 16'h7e7e;
    SB_CARRY add_4455_2 (.CI(GND_net), .I0(n29_adj_3724), .I1(n122_adj_3725), 
            .CO(n36405));
    SB_LUT4 add_4454_25_lut (.I0(GND_net), .I1(n8912[22]), .I2(GND_net), 
            .I3(n36404), .O(n8886[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_9_lut (.I0(GND_net), .I1(n8654[6]), .I2(GND_net), 
            .I3(n36049), .O(n8640[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_9 (.CI(n36049), .I0(n8654[6]), .I1(GND_net), .CO(n36050));
    SB_LUT4 mult_14_i340_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i340_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4442_8_lut (.I0(GND_net), .I1(n8654[5]), .I2(n737), .I3(n36048), 
            .O(n8640[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_15_lut (.I0(GND_net), .I1(n66[13]), .I2(n191[13]), 
            .I3(n34880), .O(\PID_CONTROLLER.result_31__N_3353 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_15 (.CI(n34880), .I0(n66[13]), .I1(n191[13]), .CO(n34881));
    SB_LUT4 add_4454_24_lut (.I0(GND_net), .I1(n8912[21]), .I2(GND_net), 
            .I3(n36403), .O(n8886[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1191__i0 (.Q(pwm_count[0]), .C(clk32MHz), .D(n70[0]));   // verilog/motorControl.v(110[18:29])
    SB_LUT4 i5_4_lut_adj_843 (.I0(\PID_CONTROLLER.result [28]), .I1(n10_adj_3723), 
            .I2(\PID_CONTROLLER.result [25]), .I3(n67[24]), .O(n12_adj_3730));   // verilog/motorControl.v(47[21:37])
    defparam i5_4_lut_adj_843.LUT_INIT = 16'hdffe;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[5]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_22_i4_3_lut (.I0(n46522), .I1(n67[1]), .I2(\PID_CONTROLLER.result [1]), 
            .I3(GND_net), .O(n4_adj_3732));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40506_3_lut (.I0(n4_adj_3732), .I1(n407), .I2(n27_adj_5), 
            .I3(GND_net), .O(n48409));   // verilog/motorControl.v(47[21:37])
    defparam i40506_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4442_8 (.CI(n36048), .I0(n8654[5]), .I1(n737), .CO(n36049));
    SB_LUT4 add_4442_7_lut (.I0(GND_net), .I1(n8654[4]), .I2(n640), .I3(n36047), 
            .O(n8640[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_25 (.CI(n36983), .I0(n6821[0]), .I1(n64[23]), 
            .CO(n36984));
    SB_CARRY add_4454_24 (.CI(n36403), .I0(n8912[21]), .I1(GND_net), .CO(n36404));
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n61[18]), 
            .I3(n34713), .O(n67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_23_lut (.I0(GND_net), .I1(n8912[20]), .I2(GND_net), 
            .I3(n36402), .O(n8886[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_20 (.CI(n34713), .I0(GND_net), .I1(n61[18]), 
            .CO(n34714));
    SB_LUT4 mult_14_add_1214_7_lut (.I0(GND_net), .I1(n1800[4]), .I2(n448_adj_3735), 
            .I3(n36800), .O(n1799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_7 (.CI(n36047), .I0(n8654[4]), .I1(n640), .CO(n36048));
    SB_CARRY sub_11_add_2_21 (.CI(n34618), .I0(\PID_CONTROLLER.err_prev[19] ), 
            .I1(n60[19]), .CO(n34619));
    SB_LUT4 i40507_3_lut (.I0(n48409), .I1(n67[14]), .I2(n29_adj_3682), 
            .I3(GND_net), .O(n48410));   // verilog/motorControl.v(47[21:37])
    defparam i40507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4472_7_lut (.I0(GND_net), .I1(n9225[4]), .I2(n472), .I3(n36647), 
            .O(n9201[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_24_lut (.I0(GND_net), .I1(n282[22]), 
            .I2(n64[22]), .I3(n36982), .O(n66[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39195_4_lut (.I0(n33_adj_3692), .I1(n31_adj_3683), .I2(n29_adj_3682), 
            .I3(n47101), .O(n47097));
    defparam i39195_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_14_add_1214_7 (.CI(n36800), .I0(n1800[4]), .I1(n448_adj_3735), 
            .CO(n36801));
    SB_CARRY add_13_add_1_28678_add_1_24 (.CI(n36982), .I0(n282[22]), .I1(n64[22]), 
            .CO(n36983));
    SB_LUT4 add_4442_6_lut (.I0(GND_net), .I1(n8654[3]), .I2(n543), .I3(n36046), 
            .O(n8640[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40952_4_lut (.I0(n30_adj_3703), .I1(n10_adj_3701), .I2(n35_adj_7), 
            .I3(n47095), .O(n48855));   // verilog/motorControl.v(47[21:37])
    defparam i40952_4_lut.LUT_INIT = 16'haaac;
    SB_DFFE \PID_CONTROLLER.integral_1192__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[0]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 i39827_3_lut (.I0(n48410), .I1(n67[15]), .I2(n31_adj_3683), 
            .I3(GND_net), .O(n47730));   // verilog/motorControl.v(47[21:37])
    defparam i39827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_28678_14_lut (.I0(GND_net), .I1(n66[12]), .I2(n191[12]), 
            .I3(n34879), .O(\PID_CONTROLLER.result_31__N_3353 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41109_4_lut (.I0(n47730), .I1(n48855), .I2(n35_adj_7), .I3(n47097), 
            .O(n49012));   // verilog/motorControl.v(47[21:37])
    defparam i41109_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41110_3_lut (.I0(n49012), .I1(n67[18]), .I2(n37_adj_3681), 
            .I3(GND_net), .O(n49013));   // verilog/motorControl.v(47[21:37])
    defparam i41110_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4442_6 (.CI(n36046), .I0(n8654[3]), .I1(n543), .CO(n36047));
    SB_LUT4 mult_14_add_1214_6_lut (.I0(GND_net), .I1(n1800[3]), .I2(n375), 
            .I3(n36799), .O(n1799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_23_lut (.I0(GND_net), .I1(n282[21]), 
            .I2(n64[21]), .I3(n36981), .O(n66[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_6 (.CI(n36799), .I0(n1800[3]), .I1(n375), 
            .CO(n36800));
    SB_LUT4 mult_14_add_1218_18_lut (.I0(GND_net), .I1(n1804[15]), .I2(GND_net), 
            .I3(n36903), .O(n1803[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_5_lut (.I0(GND_net), .I1(n8654[2]), .I2(n446), .I3(n36045), 
            .O(n8640[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[18] ), 
            .I2(n60[18]), .I3(n34617), .O(n58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41063_3_lut (.I0(n49013), .I1(n401), .I2(n39_adj_10), .I3(GND_net), 
            .O(n48966));   // verilog/motorControl.v(47[21:37])
    defparam i41063_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28678_14 (.CI(n34879), .I0(n66[12]), .I1(n191[12]), .CO(n34880));
    SB_LUT4 mult_14_add_1214_5_lut (.I0(GND_net), .I1(n1800[2]), .I2(n302), 
            .I3(n36798), .O(n1799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_7 (.CI(n36647), .I0(n9225[4]), .I1(n472), .CO(n36648));
    SB_CARRY add_4454_23 (.CI(n36402), .I0(n8912[20]), .I1(GND_net), .CO(n36403));
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n61[17]), 
            .I3(n34712), .O(n403)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_22_lut (.I0(GND_net), .I1(n8912[19]), .I2(GND_net), 
            .I3(n36401), .O(n8886[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_5 (.CI(n36045), .I0(n8654[2]), .I1(n446), .CO(n36046));
    SB_LUT4 add_4442_4_lut (.I0(GND_net), .I1(n8654[1]), .I2(n349), .I3(n36044), 
            .O(n8640[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39187_4_lut (.I0(n43_adj_3680), .I1(n41_adj_3676), .I2(n39_adj_10), 
            .I3(n48912), .O(n47089));
    defparam i39187_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_28678_13_lut (.I0(GND_net), .I1(n66[11]), .I2(n191[11]), 
            .I3(n34878), .O(\PID_CONTROLLER.result_31__N_3353 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41147_4_lut (.I0(n47728), .I1(n48928), .I2(n45_adj_3678), 
            .I3(n47087), .O(n49050));   // verilog/motorControl.v(47[21:37])
    defparam i41147_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[6]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39833_3_lut (.I0(n48966), .I1(n67[20]), .I2(n41_adj_3676), 
            .I3(GND_net), .O(n47736));   // verilog/motorControl.v(47[21:37])
    defparam i39833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41165_4_lut (.I0(n47736), .I1(n49050), .I2(n45_adj_3678), 
            .I3(n47089), .O(n49068));   // verilog/motorControl.v(47[21:37])
    defparam i41165_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n34712), .I0(GND_net), .I1(n61[17]), 
            .CO(n34713));
    SB_CARRY add_4454_22 (.CI(n36401), .I0(n8912[19]), .I1(GND_net), .CO(n36402));
    SB_CARRY mult_14_add_1218_18 (.CI(n36903), .I0(n1804[15]), .I1(GND_net), 
            .CO(n36904));
    SB_LUT4 add_4454_21_lut (.I0(GND_net), .I1(n8912[18]), .I2(GND_net), 
            .I3(n36400), .O(n8886[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4442_4 (.CI(n36044), .I0(n8654[1]), .I1(n349), .CO(n36045));
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[7]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4472_6_lut (.I0(GND_net), .I1(n9225[3]), .I2(n399), .I3(n36646), 
            .O(n9201[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_23 (.CI(n36981), .I0(n282[21]), .I1(n64[21]), 
            .CO(n36982));
    SB_LUT4 i6_4_lut_adj_844 (.I0(\PID_CONTROLLER.result [29]), .I1(n12_adj_3730), 
            .I2(n8_adj_3728), .I3(n67[24]), .O(n43824));   // verilog/motorControl.v(47[21:37])
    defparam i6_4_lut_adj_844.LUT_INIT = 16'hfdfe;
    SB_CARRY mult_14_add_1214_5 (.CI(n36798), .I0(n1800[2]), .I1(n302), 
            .CO(n36799));
    SB_CARRY add_4454_21 (.CI(n36400), .I0(n8912[18]), .I1(GND_net), .CO(n36401));
    SB_LUT4 i41166_3_lut (.I0(n49068), .I1(n67[23]), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n49069));   // verilog/motorControl.v(47[21:37])
    defparam i41166_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i41884_4_lut (.I0(n49069), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n67[24]), .I3(n43824), .O(n49785));   // verilog/motorControl.v(47[21:37])
    defparam i41884_4_lut.LUT_INIT = 16'h3371;
    SB_LUT4 add_4442_3_lut (.I0(GND_net), .I1(n8654[0]), .I2(n252), .I3(n36043), 
            .O(n8640[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4442_3 (.CI(n36043), .I0(n8654[0]), .I1(n252), .CO(n36044));
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[8]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i154_2_lut (.I0(\Kd[2] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n228_adj_3613));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i154_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4472_6 (.CI(n36646), .I0(n9225[3]), .I1(n399), .CO(n36647));
    SB_LUT4 add_4472_5_lut (.I0(GND_net), .I1(n9225[2]), .I2(n326), .I3(n36645), 
            .O(n9201[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4442_2_lut (.I0(GND_net), .I1(n62), .I2(n155_adj_3741), 
            .I3(GND_net), .O(n8640[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4442_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_20_lut (.I0(GND_net), .I1(n8912[17]), .I2(GND_net), 
            .I3(n36399), .O(n8886[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_20 (.CI(n36399), .I0(n8912[17]), .I1(GND_net), .CO(n36400));
    SB_CARRY add_4442_2 (.CI(GND_net), .I0(n62), .I1(n155_adj_3741), .CO(n36043));
    SB_CARRY add_28678_13 (.CI(n34878), .I0(n66[11]), .I1(n191[11]), .CO(n34879));
    SB_CARRY sub_11_add_2_20 (.CI(n34617), .I0(\PID_CONTROLLER.err_prev[18] ), 
            .I1(n60[18]), .CO(n34618));
    SB_LUT4 add_4454_19_lut (.I0(GND_net), .I1(n8912[16]), .I2(GND_net), 
            .I3(n36398), .O(n8886[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_17_lut (.I0(GND_net), .I1(n1804[14]), .I2(GND_net), 
            .I3(n36902), .O(n1803[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_4_lut (.I0(GND_net), .I1(n1800[1]), .I2(n229_adj_3743), 
            .I3(n36797), .O(n1799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_5 (.CI(n36645), .I0(n9225[2]), .I1(n326), .CO(n36646));
    SB_CARRY add_4454_19 (.CI(n36398), .I0(n8912[16]), .I1(GND_net), .CO(n36399));
    SB_LUT4 mult_12_i67_2_lut (.I0(\Kd[1] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_28678_12_lut (.I0(GND_net), .I1(n66[10]), .I2(n191[10]), 
            .I3(n34877), .O(\PID_CONTROLLER.result_31__N_3353 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_12 (.CI(n34877), .I0(n66[10]), .I1(n191[10]), .CO(n34878));
    SB_LUT4 add_4454_18_lut (.I0(GND_net), .I1(n8912[15]), .I2(GND_net), 
            .I3(n36397), .O(n8886[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i219_2_lut (.I0(\Kd[3] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n325));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i4_2_lut (.I0(\Kd[0] ), .I1(n58[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3483));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[17] ), 
            .I2(n60[17]), .I3(n34616), .O(n58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_11_lut (.I0(GND_net), .I1(n66[9]), .I2(n191[9]), 
            .I3(n34876), .O(\PID_CONTROLLER.result_31__N_3353 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[9]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n61[16]), 
            .I3(n34711), .O(n67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i284_2_lut (.I0(\Kd[4] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n422));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i132_2_lut (.I0(\Kd[2] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i132_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_21_add_3_18 (.CI(n34711), .I0(GND_net), .I1(n61[16]), 
            .CO(n34712));
    SB_LUT4 add_4441_14_lut (.I0(GND_net), .I1(n8640[11]), .I2(GND_net), 
            .I3(n36042), .O(n8625[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_11 (.CI(n34876), .I0(n66[9]), .I1(n191[9]), .CO(n34877));
    SB_LUT4 add_28678_10_lut (.I0(GND_net), .I1(n66[8]), .I2(n191[8]), 
            .I3(n34875), .O(\PID_CONTROLLER.result_31__N_3353 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n61[15]), 
            .I3(n34710), .O(n67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n34710), .I0(GND_net), .I1(n61[15]), 
            .CO(n34711));
    SB_CARRY add_28678_10 (.CI(n34875), .I0(n66[8]), .I1(n191[8]), .CO(n34876));
    SB_LUT4 mult_12_i349_2_lut (.I0(\Kd[5] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n519));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4472_4_lut (.I0(GND_net), .I1(n9225[1]), .I2(n253), .I3(n36644), 
            .O(n9201[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_18 (.CI(n36397), .I0(n8912[15]), .I1(GND_net), .CO(n36398));
    SB_LUT4 add_4454_17_lut (.I0(GND_net), .I1(n8912[14]), .I2(GND_net), 
            .I3(n36396), .O(n8886[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_13_lut (.I0(GND_net), .I1(n8640[10]), .I2(GND_net), 
            .I3(n36041), .O(n8625[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[10]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4441_13 (.CI(n36041), .I0(n8640[10]), .I1(GND_net), .CO(n36042));
    SB_LUT4 mult_12_i414_2_lut (.I0(\Kd[6] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n616));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i197_2_lut (.I0(\Kd[3] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n292));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_28678_9_lut (.I0(GND_net), .I1(n66[7]), .I2(n191[7]), 
            .I3(n34874), .O(\PID_CONTROLLER.result_31__N_3353 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28678_9 (.CI(n34874), .I0(n66[7]), .I1(n191[7]), .CO(n34875));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n61[14]), 
            .I3(n34709), .O(n67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_12_lut (.I0(GND_net), .I1(n8640[9]), .I2(GND_net), 
            .I3(n36040), .O(n8625[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_8_lut (.I0(GND_net), .I1(n66[6]), .I2(n191[6]), 
            .I3(n34873), .O(\PID_CONTROLLER.result_31__N_3353 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_17 (.CI(n36396), .I0(n8912[14]), .I1(GND_net), .CO(n36397));
    SB_CARRY add_28678_8 (.CI(n34873), .I0(n66[6]), .I1(n191[6]), .CO(n34874));
    SB_LUT4 add_28678_7_lut (.I0(GND_net), .I1(n66[5]), .I2(n191[5]), 
            .I3(n34872), .O(\PID_CONTROLLER.result_31__N_3353 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_19 (.CI(n34616), .I0(\PID_CONTROLLER.err_prev[17] ), 
            .I1(n60[17]), .CO(n34617));
    SB_CARRY add_28678_7 (.CI(n34872), .I0(n66[5]), .I1(n191[5]), .CO(n34873));
    SB_CARRY unary_minus_21_add_3_16 (.CI(n34709), .I0(GND_net), .I1(n61[14]), 
            .CO(n34710));
    SB_LUT4 sub_11_add_2_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[16] ), 
            .I2(n60[16]), .I3(n34615), .O(n58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_18 (.CI(n34615), .I0(\PID_CONTROLLER.err_prev[16] ), 
            .I1(n60[16]), .CO(n34616));
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n61[13]), 
            .I3(n34708), .O(n407)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28678_6_lut (.I0(GND_net), .I1(n66[4]), .I2(n191[4]), 
            .I3(n34871), .O(\PID_CONTROLLER.result_31__N_3353 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_4 (.CI(n36797), .I0(n1800[1]), .I1(n229_adj_3743), 
            .CO(n36798));
    SB_LUT4 mult_10_i144_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n213));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i144_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4472_4 (.CI(n36644), .I0(n9225[1]), .I1(n253), .CO(n36645));
    SB_LUT4 i20698_1_lut (.I0(pwm_count[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25958));   // verilog/motorControl.v(110[18:29])
    defparam i20698_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i1_1_lut (.I0(pwm[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[0]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[11]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4472_3_lut (.I0(GND_net), .I1(n9225[0]), .I2(n180_adj_3549), 
            .I3(n36643), .O(n9201[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_16_lut (.I0(GND_net), .I1(n8912[13]), .I2(GND_net), 
            .I3(n36395), .O(n8886[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_3_lut (.I0(GND_net), .I1(n1800[0]), .I2(n156_adj_3746), 
            .I3(n36796), .O(n1799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i479_2_lut (.I0(\Kd[7] ), .I1(n58[11]), .I2(GND_net), 
            .I3(GND_net), .O(n713));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i479_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_28678_6 (.CI(n34871), .I0(n66[4]), .I1(n191[4]), .CO(n34872));
    SB_LUT4 unary_minus_70_inv_0_i2_1_lut (.I0(pwm[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[1]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4454_16 (.CI(n36395), .I0(n8912[13]), .I1(GND_net), .CO(n36396));
    SB_LUT4 mult_10_i209_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n310_adj_3480));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i262_2_lut (.I0(\Kd[4] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n389));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i262_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n34708), .I0(GND_net), .I1(n61[13]), 
            .CO(n34709));
    SB_CARRY mult_14_add_1218_17 (.CI(n36902), .I0(n1804[14]), .I1(GND_net), 
            .CO(n36903));
    SB_LUT4 unary_minus_70_inv_0_i3_1_lut (.I0(pwm[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[2]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i274_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n407_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i4_1_lut (.I0(pwm[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[3]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[12]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4441_12 (.CI(n36040), .I0(n8640[9]), .I1(GND_net), .CO(n36041));
    SB_LUT4 add_4454_15_lut (.I0(GND_net), .I1(n8912[12]), .I2(GND_net), 
            .I3(n36394), .O(n8886[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_3 (.CI(n36643), .I0(n9225[0]), .I1(n180_adj_3549), 
            .CO(n36644));
    SB_LUT4 add_28678_5_lut (.I0(GND_net), .I1(n66[3]), .I2(n191[3]), 
            .I3(n34870), .O(\PID_CONTROLLER.result_31__N_3353 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_inv_0_i5_1_lut (.I0(pwm[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[4]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4454_15 (.CI(n36394), .I0(n8912[12]), .I1(GND_net), .CO(n36395));
    SB_LUT4 add_4454_14_lut (.I0(GND_net), .I1(n8912[11]), .I2(GND_net), 
            .I3(n36393), .O(n8886[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i339_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n504));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i6_1_lut (.I0(pwm[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[5]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i327_2_lut (.I0(\Kd[5] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n486));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n601_adj_3478));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i7_1_lut (.I0(pwm[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[6]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i8_1_lut (.I0(pwm[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[7]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1214_3 (.CI(n36796), .I0(n1800[0]), .I1(n156_adj_3746), 
            .CO(n36797));
    SB_LUT4 add_13_add_1_28678_add_1_22_lut (.I0(GND_net), .I1(n282[20]), 
            .I2(n64[20]), .I3(n36980), .O(n66[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_11_lut (.I0(GND_net), .I1(n8640[8]), .I2(GND_net), 
            .I3(n36039), .O(n8625[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_2_lut (.I0(GND_net), .I1(n14_adj_3747), .I2(n83_adj_3748), 
            .I3(GND_net), .O(n1799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_11 (.CI(n36039), .I0(n8640[8]), .I1(GND_net), .CO(n36040));
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n698));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4472_2_lut (.I0(GND_net), .I1(n35_adj_3550), .I2(n107), 
            .I3(GND_net), .O(n9201[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_inv_0_i9_1_lut (.I0(pwm[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[8]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4441_10_lut (.I0(GND_net), .I1(n8640[7]), .I2(GND_net), 
            .I3(n36038), .O(n8625[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_16_lut (.I0(GND_net), .I1(n1804[13]), .I2(GND_net), 
            .I3(n36901), .O(n1803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n61[12]), 
            .I3(n34707), .O(n67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_14 (.CI(n34707), .I0(GND_net), .I1(n61[12]), 
            .CO(n34708));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n61[11]), 
            .I3(n34706), .O(n67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_22 (.CI(n36980), .I0(n282[20]), .I1(n64[20]), 
            .CO(n36981));
    SB_CARRY add_28678_5 (.CI(n34870), .I0(n66[3]), .I1(n191[3]), .CO(n34871));
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3593));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i392_2_lut (.I0(\Kd[6] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n583));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_28678_4_lut (.I0(GND_net), .I1(n66[2]), .I2(n191[2]), 
            .I3(n34869), .O(\PID_CONTROLLER.result_31__N_3353 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3592));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i136_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_3591));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i95_2_lut (.I0(\Kd[1] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n140));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i32_2_lut (.I0(\Kd[0] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4441_10 (.CI(n36038), .I0(n8640[7]), .I1(GND_net), .CO(n36039));
    SB_LUT4 unary_minus_70_inv_0_i10_1_lut (.I0(pwm[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n63[9]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4441_9_lut (.I0(GND_net), .I1(n8640[6]), .I2(GND_net), 
            .I3(n36037), .O(n8625[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_21_lut (.I0(GND_net), .I1(n282[19]), 
            .I2(n64[19]), .I3(n36979), .O(n66[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i201_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_3589));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i201_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4472_2 (.CI(GND_net), .I0(n35_adj_3550), .I1(n107), .CO(n36643));
    SB_CARRY add_4454_14 (.CI(n36393), .I0(n8912[11]), .I1(GND_net), .CO(n36394));
    SB_CARRY add_28678_4 (.CI(n34869), .I0(n66[2]), .I1(n191[2]), .CO(n34870));
    SB_LUT4 unary_minus_17_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[13]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4441_9 (.CI(n36037), .I0(n8640[6]), .I1(GND_net), .CO(n36038));
    SB_CARRY unary_minus_21_add_3_13 (.CI(n34706), .I0(GND_net), .I1(n61[11]), 
            .CO(n34707));
    SB_CARRY mult_14_add_1218_16 (.CI(n36901), .I0(n1804[13]), .I1(GND_net), 
            .CO(n36902));
    SB_LUT4 add_28678_3_lut (.I0(GND_net), .I1(n66[1]), .I2(n191[1]), 
            .I3(n34868), .O(\PID_CONTROLLER.result_31__N_3353 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i266_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n395_adj_3588));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4441_8_lut (.I0(GND_net), .I1(n8640[5]), .I2(n734), .I3(n36036), 
            .O(n8625[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_21 (.CI(n36979), .I0(n282[19]), .I1(n64[19]), 
            .CO(n36980));
    SB_LUT4 add_4454_13_lut (.I0(GND_net), .I1(n8912[10]), .I2(GND_net), 
            .I3(n36392), .O(n8886[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i331_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n492_adj_3587));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i11_1_lut (.I0(pwm[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[10]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4441_8 (.CI(n36036), .I0(n8640[5]), .I1(n734), .CO(n36037));
    SB_LUT4 add_13_add_1_28678_add_1_20_lut (.I0(GND_net), .I1(n282[18]), 
            .I2(n64[18]), .I3(n36978), .O(n66[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_20 (.CI(n36978), .I0(n282[18]), .I1(n64[18]), 
            .CO(n36979));
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n589_adj_3585));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1218_15_lut (.I0(GND_net), .I1(n1804[12]), .I2(GND_net), 
            .I3(n36900), .O(n1803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_2 (.CI(GND_net), .I0(n14_adj_3747), .I1(n83_adj_3748), 
            .CO(n36796));
    SB_LUT4 add_4441_7_lut (.I0(GND_net), .I1(n8640[4]), .I2(n637), .I3(n36035), 
            .O(n8625[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_13 (.CI(n36392), .I0(n8912[10]), .I1(GND_net), .CO(n36393));
    SB_CARRY add_4441_7 (.CI(n36035), .I0(n8640[4]), .I1(n637), .CO(n36036));
    SB_LUT4 add_4471_8_lut (.I0(GND_net), .I1(n9547[5]), .I2(n752_adj_3752), 
            .I3(n36642), .O(n9192[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n686_adj_3584));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_28678_3 (.CI(n34868), .I0(n66[1]), .I1(n191[1]), .CO(n34869));
    SB_LUT4 add_28678_2_lut (.I0(GND_net), .I1(n66[0]), .I2(n191[0]), 
            .I3(GND_net), .O(\PID_CONTROLLER.result_31__N_3353 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_28678_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_12_lut (.I0(GND_net), .I1(n8912[9]), .I2(GND_net), 
            .I3(n36391), .O(n8886[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4441_6_lut (.I0(GND_net), .I1(n8640[3]), .I2(n540), .I3(n36034), 
            .O(n8625[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_12 (.CI(n36391), .I0(n8912[9]), .I1(GND_net), .CO(n36392));
    SB_LUT4 mult_12_i91_2_lut (.I0(\Kd[1] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n134));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i91_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_15 (.CI(n36900), .I0(n1804[12]), .I1(GND_net), 
            .CO(n36901));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n61[10]), 
            .I3(n34705), .O(n410)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n34705), .I0(GND_net), .I1(n61[10]), 
            .CO(n34706));
    SB_LUT4 sub_11_add_2_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[15] ), 
            .I2(n60[15]), .I3(n34614), .O(n58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_24_lut (.I0(GND_net), .I1(n1799[21]), .I2(GND_net), 
            .I3(n36794), .O(n1798[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4471_7_lut (.I0(GND_net), .I1(n9547[4]), .I2(n655_adj_3754), 
            .I3(n36641), .O(n9192[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4471_7 (.CI(n36641), .I0(n9547[4]), .I1(n655_adj_3754), 
            .CO(n36642));
    SB_CARRY add_4441_6 (.CI(n36034), .I0(n8640[3]), .I1(n540), .CO(n36035));
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n61[9]), 
            .I3(n34704), .O(n67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i28_2_lut (.I0(\Kd[0] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3583));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i12_1_lut (.I0(pwm[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[11]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_28678_2 (.CI(GND_net), .I0(n66[0]), .I1(n191[0]), .CO(n34868));
    SB_LUT4 mult_12_i156_2_lut (.I0(\Kd[2] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n231_adj_3581));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i13_1_lut (.I0(pwm[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[12]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i221_2_lut (.I0(\Kd[3] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n328));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i14_1_lut (.I0(pwm[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[13]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n34704), .I0(GND_net), .I1(n61[9]), 
            .CO(n34705));
    SB_LUT4 add_4441_5_lut (.I0(GND_net), .I1(n8640[2]), .I2(n443_adj_3755), 
            .I3(n36033), .O(n8625[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n61[8]), 
            .I3(n34703), .O(n67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_5 (.CI(n36033), .I0(n8640[2]), .I1(n443_adj_3755), 
            .CO(n36034));
    SB_LUT4 mult_12_i286_2_lut (.I0(\Kd[4] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n425));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i15_1_lut (.I0(pwm[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[14]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i16_1_lut (.I0(pwm[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[15]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i457_2_lut (.I0(\Kd[7] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n680));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n35519), .O(n73[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n35518), .O(n73[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_11_lut (.I0(GND_net), .I1(n8912[8]), .I2(GND_net), 
            .I3(n36390), .O(n8886[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n34703), .I0(GND_net), .I1(n61[8]), 
            .CO(n34704));
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_10  (.CI(n35518), .I0(\PID_CONTROLLER.err[8] ), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n35519));
    SB_LUT4 add_13_add_1_28678_add_1_19_lut (.I0(GND_net), .I1(n282[17]), 
            .I2(n64[17]), .I3(n36977), .O(n66[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i351_2_lut (.I0(\Kd[5] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n522));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i17_1_lut (.I0(pwm[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[16]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_13_add_1_28678_add_1_19 (.CI(n36977), .I0(n282[17]), .I1(n64[17]), 
            .CO(n36978));
    SB_LUT4 add_4441_4_lut (.I0(GND_net), .I1(n8640[1]), .I2(n346), .I3(n36032), 
            .O(n8625[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_11 (.CI(n36390), .I0(n8912[8]), .I1(GND_net), .CO(n36391));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n35517), .O(n73[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_4 (.CI(n36032), .I0(n8640[1]), .I1(n346), .CO(n36033));
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_9  (.CI(n35517), .I0(\PID_CONTROLLER.err[7] ), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n35518));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n35516), .O(n73[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_18_lut (.I0(GND_net), .I1(n282[16]), 
            .I2(n64[16]), .I3(n36976), .O(n66[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_14_lut (.I0(GND_net), .I1(n1804[11]), .I2(GND_net), 
            .I3(n36899), .O(n1803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_18 (.CI(n36976), .I0(n282[16]), .I1(n64[16]), 
            .CO(n36977));
    SB_LUT4 add_4441_3_lut (.I0(GND_net), .I1(n8640[0]), .I2(n249), .I3(n36031), 
            .O(n8625[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i160_2_lut (.I0(\Kd[2] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n237_adj_3476));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[14]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_8  (.CI(n35516), .I0(\PID_CONTROLLER.err[6] ), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n35517));
    SB_LUT4 mult_12_i225_2_lut (.I0(\Kd[3] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n334));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i225_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_14 (.CI(n36899), .I0(n1804[11]), .I1(GND_net), 
            .CO(n36900));
    SB_LUT4 unary_minus_17_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[15]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i290_2_lut (.I0(\Kd[4] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n431));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i389_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n35515), .O(n73[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_3 (.CI(n36031), .I0(n8640[0]), .I1(n249), .CO(n36032));
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_7  (.CI(n35515), .I0(\PID_CONTROLLER.err[5] ), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n35516));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n35514), .O(n73[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_13_lut (.I0(GND_net), .I1(n1804[10]), .I2(GND_net), 
            .I3(n36898), .O(n1803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i355_2_lut (.I0(\Kd[5] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n528));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_24 (.CI(n36794), .I0(n1799[21]), .I1(GND_net), 
            .CO(n1691));
    SB_LUT4 mult_14_add_1213_23_lut (.I0(GND_net), .I1(n1799[20]), .I2(GND_net), 
            .I3(n36793), .O(n1798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_6  (.CI(n35514), .I0(\PID_CONTROLLER.err[4] ), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n35515));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n35513), .O(n73[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4471_6_lut (.I0(GND_net), .I1(n9547[3]), .I2(n558), .I3(n36640), 
            .O(n9192[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_10_lut (.I0(GND_net), .I1(n8912[7]), .I2(GND_net), 
            .I3(n36389), .O(n8886[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_10 (.CI(n36389), .I0(n8912[7]), .I1(GND_net), .CO(n36390));
    SB_CARRY sub_11_add_2_17 (.CI(n34614), .I0(\PID_CONTROLLER.err_prev[15] ), 
            .I1(n60[15]), .CO(n34615));
    SB_LUT4 mult_10_i146_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n216));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i211_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n313_adj_3473));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i18_1_lut (.I0(pwm[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[17]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i420_2_lut (.I0(\Kd[6] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n625));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i416_2_lut (.I0(\Kd[6] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n619));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i276_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n410_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4441_2_lut (.I0(GND_net), .I1(n59), .I2(n152_adj_3759), 
            .I3(GND_net), .O(n8625[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4441_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_17_lut (.I0(GND_net), .I1(n282[15]), 
            .I2(n64[15]), .I3(n36975), .O(n66[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i341_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n507));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i341_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_5  (.CI(n35513), .I0(\PID_CONTROLLER.err[3] ), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n35514));
    SB_CARRY mult_14_add_1218_13 (.CI(n36898), .I0(n1804[10]), .I1(GND_net), 
            .CO(n36899));
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n604));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[14] ), 
            .I2(n60[14]), .I3(n34613), .O(n58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_16 (.CI(n34613), .I0(\PID_CONTROLLER.err_prev[14] ), 
            .I1(n60[14]), .CO(n34614));
    SB_CARRY mult_14_add_1213_23 (.CI(n36793), .I0(n1799[20]), .I1(GND_net), 
            .CO(n36794));
    SB_CARRY add_4471_6 (.CI(n36640), .I0(n9547[3]), .I1(n558), .CO(n36641));
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n701));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n35512), .O(n73[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_9_lut (.I0(GND_net), .I1(n8912[6]), .I2(GND_net), 
            .I3(n36388), .O(n8886[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_22_lut (.I0(GND_net), .I1(n1799[19]), .I2(GND_net), 
            .I3(n36792), .O(n1798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4441_2 (.CI(GND_net), .I0(n59), .I1(n152_adj_3759), .CO(n36031));
    SB_LUT4 add_4440_15_lut (.I0(GND_net), .I1(n8625[12]), .I2(GND_net), 
            .I3(n36030), .O(n8609[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i485_2_lut (.I0(\Kd[7] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n722));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i485_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_4  (.CI(n35512), .I0(\PID_CONTROLLER.err[2] ), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n35513));
    SB_LUT4 unary_minus_70_inv_0_i19_1_lut (.I0(pwm[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[18]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4471_5_lut (.I0(GND_net), .I1(n9547[2]), .I2(n461), .I3(n36639), 
            .O(n9192[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4471_5 (.CI(n36639), .I0(n9547[2]), .I1(n461), .CO(n36640));
    SB_LUT4 mult_14_add_1218_12_lut (.I0(GND_net), .I1(n1804[9]), .I2(GND_net), 
            .I3(n36897), .O(n1803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4471_4_lut (.I0(GND_net), .I1(n9547[1]), .I2(n364_adj_3762), 
            .I3(n36638), .O(n9192[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[13] ), 
            .I2(n60[13]), .I3(n34612), .O(n58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_15 (.CI(n34612), .I0(\PID_CONTROLLER.err_prev[13] ), 
            .I1(n60[13]), .CO(n34613));
    SB_CARRY mult_14_add_1213_22 (.CI(n36792), .I0(n1799[19]), .I1(GND_net), 
            .CO(n36793));
    SB_LUT4 mult_14_add_1213_21_lut (.I0(GND_net), .I1(n1799[18]), .I2(GND_net), 
            .I3(n36791), .O(n1798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_21 (.CI(n36791), .I0(n1799[18]), .I1(GND_net), 
            .CO(n36792));
    SB_CARRY add_4471_4 (.CI(n36638), .I0(n9547[1]), .I1(n364_adj_3762), 
            .CO(n36639));
    SB_LUT4 add_4471_3_lut (.I0(GND_net), .I1(n9547[0]), .I2(n267), .I3(n36637), 
            .O(n9192[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_9 (.CI(n36388), .I0(n8912[6]), .I1(GND_net), .CO(n36389));
    SB_LUT4 add_4440_14_lut (.I0(GND_net), .I1(n8625[11]), .I2(GND_net), 
            .I3(n36029), .O(n8609[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4454_8_lut (.I0(GND_net), .I1(n8912[5]), .I2(n701_adj_3764), 
            .I3(n36387), .O(n8886[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_14 (.CI(n36029), .I0(n8625[11]), .I1(GND_net), .CO(n36030));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n35511), .O(n73[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_8 (.CI(n36387), .I0(n8912[5]), .I1(n701_adj_3764), 
            .CO(n36388));
    SB_LUT4 mult_12_i481_2_lut (.I0(\Kd[7] ), .I1(n58[12]), .I2(GND_net), 
            .I3(GND_net), .O(n716));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i20_1_lut (.I0(pwm[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[19]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4454_7_lut (.I0(GND_net), .I1(n8912[4]), .I2(n604_adj_3766), 
            .I3(n36386), .O(n8886[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_20_lut (.I0(GND_net), .I1(n1799[17]), .I2(GND_net), 
            .I3(n36790), .O(n1798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_12 (.CI(n36897), .I0(n1804[9]), .I1(GND_net), 
            .CO(n36898));
    SB_LUT4 add_4440_13_lut (.I0(GND_net), .I1(n8625[10]), .I2(GND_net), 
            .I3(n36028), .O(n8609[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_3  (.CI(n35511), .I0(\PID_CONTROLLER.err[1] ), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n35512));
    SB_CARRY add_4471_3 (.CI(n36637), .I0(n9547[0]), .I1(n267), .CO(n36638));
    SB_CARRY add_4454_7 (.CI(n36386), .I0(n8912[4]), .I1(n604_adj_3766), 
            .CO(n36387));
    SB_LUT4 add_4471_2_lut (.I0(GND_net), .I1(n83), .I2(n170_adj_3767), 
            .I3(GND_net), .O(n9192[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4471_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_17 (.CI(n36975), .I0(n282[15]), .I1(n64[15]), 
            .CO(n36976));
    SB_LUT4 \PID_CONTROLLER.integral_1192_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n73[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1192_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_13 (.CI(n36028), .I0(n8625[10]), .I1(GND_net), .CO(n36029));
    SB_LUT4 mult_14_add_1218_11_lut (.I0(GND_net), .I1(n1804[8]), .I2(GND_net), 
            .I3(n36896), .O(n1803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1192_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err[0] ), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n35511));
    SB_LUT4 sub_11_add_2_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[12] ), 
            .I2(n60[12]), .I3(n34611), .O(n58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4471_2 (.CI(GND_net), .I0(n83), .I1(n170_adj_3767), .CO(n36637));
    SB_LUT4 add_4454_6_lut (.I0(GND_net), .I1(n8912[3]), .I2(n507_adj_3769), 
            .I3(n36385), .O(n8886[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_20 (.CI(n36790), .I0(n1799[17]), .I1(GND_net), 
            .CO(n36791));
    SB_LUT4 add_4440_12_lut (.I0(GND_net), .I1(n8625[9]), .I2(GND_net), 
            .I3(n36027), .O(n8609[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_12 (.CI(n36027), .I0(n8625[9]), .I1(GND_net), .CO(n36028));
    SB_LUT4 add_4470_9_lut (.I0(GND_net), .I1(n9192[6]), .I2(GND_net), 
            .I3(n36636), .O(n9182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4454_6 (.CI(n36385), .I0(n8912[3]), .I1(n507_adj_3769), 
            .CO(n36386));
    SB_LUT4 add_4470_8_lut (.I0(GND_net), .I1(n9192[5]), .I2(n749_adj_3770), 
            .I3(n36635), .O(n9182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4454_5_lut (.I0(GND_net), .I1(n8912[2]), .I2(n410_adj_3771), 
            .I3(n36384), .O(n8886[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4440_11_lut (.I0(GND_net), .I1(n8625[8]), .I2(GND_net), 
            .I3(n36026), .O(n8609[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3571));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i21_1_lut (.I0(pwm[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[20]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i22_1_lut (.I0(pwm[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[21]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i23_1_lut (.I0(pwm[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[22]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1213_19_lut (.I0(GND_net), .I1(n1799[16]), .I2(GND_net), 
            .I3(n36789), .O(n1798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_11 (.CI(n36026), .I0(n8625[8]), .I1(GND_net), .CO(n36027));
    SB_CARRY add_4470_8 (.CI(n36635), .I0(n9192[5]), .I1(n749_adj_3770), 
            .CO(n36636));
    SB_CARRY add_4454_5 (.CI(n36384), .I0(n8912[2]), .I1(n410_adj_3771), 
            .CO(n36385));
    SB_CARRY sub_11_add_2_14 (.CI(n34611), .I0(\PID_CONTROLLER.err_prev[12] ), 
            .I1(n60[12]), .CO(n34612));
    SB_LUT4 add_4440_10_lut (.I0(GND_net), .I1(n8625[7]), .I2(GND_net), 
            .I3(n36025), .O(n8609[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_10 (.CI(n36025), .I0(n8625[7]), .I1(GND_net), .CO(n36026));
    SB_LUT4 sub_11_add_2_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[11] ), 
            .I2(n60[11]), .I3(n34610), .O(n58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_13 (.CI(n34610), .I0(\PID_CONTROLLER.err_prev[11] ), 
            .I1(n60[11]), .CO(n34611));
    SB_LUT4 add_4440_9_lut (.I0(GND_net), .I1(n8625[6]), .I2(GND_net), 
            .I3(n36024), .O(n8609[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20697_1_lut (.I0(\PID_CONTROLLER.result [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25957));   // verilog/motorControl.v(38[14] 59[8])
    defparam i20697_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4454_4_lut (.I0(GND_net), .I1(n8912[1]), .I2(n313_adj_3773), 
            .I3(n36383), .O(n8886[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_9 (.CI(n36024), .I0(n8625[6]), .I1(GND_net), .CO(n36025));
    SB_LUT4 add_4440_8_lut (.I0(GND_net), .I1(n8625[5]), .I2(n731), .I3(n36023), 
            .O(n8609[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_16_lut (.I0(GND_net), .I1(n282[14]), 
            .I2(n64[14]), .I3(n36974), .O(n66[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3468));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4454_4 (.CI(n36383), .I0(n8912[1]), .I1(n313_adj_3773), 
            .CO(n36384));
    SB_CARRY mult_14_add_1218_11 (.CI(n36896), .I0(n1804[8]), .I1(GND_net), 
            .CO(n36897));
    SB_LUT4 mult_14_add_1218_10_lut (.I0(GND_net), .I1(n1804[7]), .I2(GND_net), 
            .I3(n36895), .O(n1803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[0]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_13_add_1_28678_add_1_16 (.CI(n36974), .I0(n282[14]), .I1(n64[14]), 
            .CO(n36975));
    SB_LUT4 mult_10_i148_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n219_adj_3466));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i213_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n316));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i213_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4440_8 (.CI(n36023), .I0(n8625[5]), .I1(n731), .CO(n36024));
    SB_LUT4 add_4470_7_lut (.I0(GND_net), .I1(n9192[4]), .I2(n652_adj_3776), 
            .I3(n36634), .O(n9182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4440_7_lut (.I0(GND_net), .I1(n8625[4]), .I2(n634), .I3(n36022), 
            .O(n8609[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3567));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i278_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n413));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i203_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n301));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i343_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n510));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i268_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n398));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i333_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n495));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n592));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n689));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3565));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[1]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n607));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3559));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i473_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n704));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i71_2_lut (.I0(\Kd[1] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i8_2_lut (.I0(\Kd[0] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n207));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i136_2_lut (.I0(\Kd[2] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n201));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i93_2_lut (.I0(\Kd[1] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n137));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i30_2_lut (.I0(\Kd[0] ), .I1(n58[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i205_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n304));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i270_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n401_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i201_2_lut (.I0(\Kd[3] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n298));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i266_2_lut (.I0(\Kd[4] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n395));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i335_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n498));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n595));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i158_2_lut (.I0(\Kd[2] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n234_adj_3556));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n692));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3555));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i223_2_lut (.I0(\Kd[3] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n331));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i223_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_10 (.CI(n36895), .I0(n1804[7]), .I1(GND_net), 
            .CO(n36896));
    SB_LUT4 mult_14_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n61[7]), 
            .I3(n34702), .O(n67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3550));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4454_3_lut (.I0(GND_net), .I1(n8912[0]), .I2(n216_adj_3777), 
            .I3(n36382), .O(n8886[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_7 (.CI(n36022), .I0(n8625[4]), .I1(n634), .CO(n36023));
    SB_LUT4 mult_12_i288_2_lut (.I0(\Kd[4] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n428));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[10] ), 
            .I2(n60[10]), .I3(n34609), .O(n58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_12 (.CI(n34609), .I0(\PID_CONTROLLER.err_prev[10] ), 
            .I1(n60[10]), .CO(n34610));
    SB_LUT4 add_4440_6_lut (.I0(GND_net), .I1(n8625[3]), .I2(n537_adj_3779), 
            .I3(n36021), .O(n8609[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_6 (.CI(n36021), .I0(n8625[3]), .I1(n537_adj_3779), 
            .CO(n36022));
    SB_CARRY unary_minus_21_add_3_9 (.CI(n34702), .I0(GND_net), .I1(n61[7]), 
            .CO(n34703));
    SB_LUT4 sub_11_add_2_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[9] ), 
            .I2(n60[9]), .I3(n34608), .O(n58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i78_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(\GATES_5__N_3398[5] ));   // verilog/motorControl.v(91[19:34])
    defparam i78_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_4454_3 (.CI(n36382), .I0(n8912[0]), .I1(n216_adj_3777), 
            .CO(n36383));
    SB_LUT4 add_4454_2_lut (.I0(GND_net), .I1(n26_adj_3781), .I2(n119_adj_3782), 
            .I3(GND_net), .O(n8886[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4454_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_15_lut (.I0(GND_net), .I1(n282[13]), 
            .I2(n64[13]), .I3(n36973), .O(n66[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_9_lut (.I0(GND_net), .I1(n1804[6]), .I2(GND_net), 
            .I3(n36894), .O(n1803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_19 (.CI(n36789), .I0(n1799[16]), .I1(GND_net), 
            .CO(n36790));
    SB_CARRY add_4470_7 (.CI(n36634), .I0(n9192[4]), .I1(n652_adj_3776), 
            .CO(n36635));
    SB_CARRY add_4454_2 (.CI(GND_net), .I0(n26_adj_3781), .I1(n119_adj_3782), 
            .CO(n36382));
    SB_LUT4 add_4440_5_lut (.I0(GND_net), .I1(n8625[2]), .I2(n440), .I3(n36020), 
            .O(n8609[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_5 (.CI(n36020), .I0(n8625[2]), .I1(n440), .CO(n36021));
    SB_LUT4 add_4453_26_lut (.I0(GND_net), .I1(n8886[23]), .I2(GND_net), 
            .I3(n36381), .O(n8859[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4440_4_lut (.I0(GND_net), .I1(n8625[1]), .I2(n343), .I3(n36019), 
            .O(n8609[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_4 (.CI(n36019), .I0(n8625[1]), .I1(n343), .CO(n36020));
    SB_LUT4 add_4470_6_lut (.I0(GND_net), .I1(n9192[3]), .I2(n555_adj_3785), 
            .I3(n36633), .O(n9182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_25_lut (.I0(GND_net), .I1(n8886[22]), .I2(GND_net), 
            .I3(n36380), .O(n8859[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4440_3_lut (.I0(GND_net), .I1(n8625[0]), .I2(n246_adj_3786), 
            .I3(n36018), .O(n8609[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_3 (.CI(n36018), .I0(n8625[0]), .I1(n246_adj_3786), 
            .CO(n36019));
    SB_CARRY add_4453_25 (.CI(n36380), .I0(n8886[22]), .I1(GND_net), .CO(n36381));
    SB_LUT4 add_4440_2_lut (.I0(GND_net), .I1(n56_adj_3787), .I2(n149_adj_3788), 
            .I3(GND_net), .O(n8609[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4440_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4440_2 (.CI(GND_net), .I0(n56_adj_3787), .I1(n149_adj_3788), 
            .CO(n36018));
    SB_LUT4 mult_14_add_1213_18_lut (.I0(GND_net), .I1(n1799[15]), .I2(GND_net), 
            .I3(n36788), .O(n1798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4470_6 (.CI(n36633), .I0(n9192[3]), .I1(n555_adj_3785), 
            .CO(n36634));
    SB_LUT4 add_4453_24_lut (.I0(GND_net), .I1(n8886[21]), .I2(GND_net), 
            .I3(n36379), .O(n8859[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_16_lut (.I0(GND_net), .I1(n8609[13]), .I2(GND_net), 
            .I3(n36017), .O(n8592[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_15_lut (.I0(GND_net), .I1(n8609[12]), .I2(GND_net), 
            .I3(n36016), .O(n8592[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1191_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[8]), 
            .I3(n35497), .O(n70[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1191_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[7]), 
            .I3(n35496), .O(n70[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_24 (.CI(n36379), .I0(n8886[21]), .I1(GND_net), .CO(n36380));
    SB_CARRY add_4439_15 (.CI(n36016), .I0(n8609[12]), .I1(GND_net), .CO(n36017));
    SB_CARRY pwm_count_1191_add_4_9 (.CI(n35496), .I0(GND_net), .I1(pwm_count[7]), 
            .CO(n35497));
    SB_LUT4 pwm_count_1191_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[6]), 
            .I3(n35495), .O(n70[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_14_lut (.I0(GND_net), .I1(n8609[11]), .I2(GND_net), 
            .I3(n36015), .O(n8592[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1191_add_4_8 (.CI(n35495), .I0(GND_net), .I1(pwm_count[6]), 
            .CO(n35496));
    SB_LUT4 pwm_count_1191_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[5]), 
            .I3(n35494), .O(n70[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4470_5_lut (.I0(GND_net), .I1(n9192[2]), .I2(n458_adj_3792), 
            .I3(n36632), .O(n9182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_23_lut (.I0(GND_net), .I1(n8886[20]), .I2(GND_net), 
            .I3(n36378), .O(n8859[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_14 (.CI(n36015), .I0(n8609[11]), .I1(GND_net), .CO(n36016));
    SB_CARRY pwm_count_1191_add_4_7 (.CI(n35494), .I0(GND_net), .I1(pwm_count[5]), 
            .CO(n35495));
    SB_LUT4 pwm_count_1191_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[4]), 
            .I3(n35493), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_13_lut (.I0(GND_net), .I1(n8609[10]), .I2(GND_net), 
            .I3(n36014), .O(n8592[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1191_add_4_6 (.CI(n35493), .I0(GND_net), .I1(pwm_count[4]), 
            .CO(n35494));
    SB_LUT4 pwm_count_1191_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[3]), 
            .I3(n35492), .O(n70[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_23 (.CI(n36378), .I0(n8886[20]), .I1(GND_net), .CO(n36379));
    SB_CARRY add_4439_13 (.CI(n36014), .I0(n8609[10]), .I1(GND_net), .CO(n36015));
    SB_CARRY pwm_count_1191_add_4_5 (.CI(n35492), .I0(GND_net), .I1(pwm_count[3]), 
            .CO(n35493));
    SB_LUT4 pwm_count_1191_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[2]), 
            .I3(n35491), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_12_lut (.I0(GND_net), .I1(n8609[9]), .I2(GND_net), 
            .I3(n36013), .O(n8592[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1191_add_4_4 (.CI(n35491), .I0(GND_net), .I1(pwm_count[2]), 
            .CO(n35492));
    SB_LUT4 pwm_count_1191_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[1]), 
            .I3(n35490), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_9 (.CI(n36894), .I0(n1804[6]), .I1(GND_net), 
            .CO(n36895));
    SB_CARRY mult_14_add_1213_18 (.CI(n36788), .I0(n1799[15]), .I1(GND_net), 
            .CO(n36789));
    SB_CARRY add_4470_5 (.CI(n36632), .I0(n9192[2]), .I1(n458_adj_3792), 
            .CO(n36633));
    SB_LUT4 add_4453_22_lut (.I0(GND_net), .I1(n8886[19]), .I2(GND_net), 
            .I3(n36377), .O(n8859[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_12 (.CI(n36013), .I0(n8609[9]), .I1(GND_net), .CO(n36014));
    SB_CARRY pwm_count_1191_add_4_3 (.CI(n35490), .I0(GND_net), .I1(pwm_count[1]), 
            .CO(n35491));
    SB_LUT4 pwm_count_1191_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[0]), 
            .I3(VCC_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4439_11_lut (.I0(GND_net), .I1(n8609[8]), .I2(GND_net), 
            .I3(n36012), .O(n8592[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_count[0]), 
            .CO(n35490));
    SB_LUT4 Kd_delay_counter_1190_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[6]), .I3(n35489), .O(n69[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_22 (.CI(n36377), .I0(n8886[19]), .I1(GND_net), .CO(n36378));
    SB_CARRY add_4439_11 (.CI(n36012), .I0(n8609[8]), .I1(GND_net), .CO(n36013));
    SB_LUT4 Kd_delay_counter_1190_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[5]), .I3(n35488), .O(n69[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_7 (.CI(n35488), .I0(GND_net), .I1(Kd_delay_counter[5]), 
            .CO(n35489));
    SB_LUT4 add_4439_10_lut (.I0(GND_net), .I1(n8609[7]), .I2(GND_net), 
            .I3(n36011), .O(n8592[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1190_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[4]), .I3(n35487), .O(n69[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_6 (.CI(n35487), .I0(GND_net), .I1(Kd_delay_counter[4]), 
            .CO(n35488));
    SB_LUT4 add_4470_4_lut (.I0(GND_net), .I1(n9192[1]), .I2(n361_adj_3799), 
            .I3(n36631), .O(n9182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_21_lut (.I0(GND_net), .I1(n8886[18]), .I2(GND_net), 
            .I3(n36376), .O(n8859[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_10 (.CI(n36011), .I0(n8609[7]), .I1(GND_net), .CO(n36012));
    SB_LUT4 Kd_delay_counter_1190_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[3]), .I3(n35486), .O(n69[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_5 (.CI(n35486), .I0(GND_net), .I1(Kd_delay_counter[3]), 
            .CO(n35487));
    SB_LUT4 add_4439_9_lut (.I0(GND_net), .I1(n8609[6]), .I2(GND_net), 
            .I3(n36010), .O(n8592[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1190_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[2]), .I3(n35485), .O(n69[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_4 (.CI(n35485), .I0(GND_net), .I1(Kd_delay_counter[2]), 
            .CO(n35486));
    SB_CARRY add_4453_21 (.CI(n36376), .I0(n8886[18]), .I1(GND_net), .CO(n36377));
    SB_CARRY add_4439_9 (.CI(n36010), .I0(n8609[6]), .I1(GND_net), .CO(n36011));
    SB_LUT4 Kd_delay_counter_1190_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[1]), .I3(n35484), .O(n69[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_3 (.CI(n35484), .I0(GND_net), .I1(Kd_delay_counter[1]), 
            .CO(n35485));
    SB_LUT4 add_4439_8_lut (.I0(GND_net), .I1(n8609[5]), .I2(n728), .I3(n36009), 
            .O(n8592[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1190_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[0]), .I3(VCC_net), .O(n69[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1190_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1190_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(Kd_delay_counter[0]), .CO(n35484));
    SB_LUT4 mult_14_add_1213_17_lut (.I0(GND_net), .I1(n1799[14]), .I2(GND_net), 
            .I3(n36787), .O(n1798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4470_4 (.CI(n36631), .I0(n9192[1]), .I1(n361_adj_3799), 
            .CO(n36632));
    SB_LUT4 add_4453_20_lut (.I0(GND_net), .I1(n8886[17]), .I2(GND_net), 
            .I3(n36375), .O(n8859[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_8 (.CI(n36009), .I0(n8609[5]), .I1(n728), .CO(n36010));
    SB_LUT4 add_4439_7_lut (.I0(GND_net), .I1(n8609[4]), .I2(n631), .I3(n36008), 
            .O(n8592[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_20 (.CI(n36375), .I0(n8886[17]), .I1(GND_net), .CO(n36376));
    SB_CARRY add_4439_7 (.CI(n36008), .I0(n8609[4]), .I1(n631), .CO(n36009));
    SB_LUT4 add_4439_6_lut (.I0(GND_net), .I1(n8609[3]), .I2(n534), .I3(n36007), 
            .O(n8592[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4470_3_lut (.I0(GND_net), .I1(n9192[0]), .I2(n264_adj_3803), 
            .I3(n36630), .O(n9182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_19_lut (.I0(GND_net), .I1(n8886[16]), .I2(GND_net), 
            .I3(n36374), .O(n8859[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_6 (.CI(n36007), .I0(n8609[3]), .I1(n534), .CO(n36008));
    SB_LUT4 add_4439_5_lut (.I0(GND_net), .I1(n8609[2]), .I2(n437_adj_3804), 
            .I3(n36006), .O(n8592[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_19 (.CI(n36374), .I0(n8886[16]), .I1(GND_net), .CO(n36375));
    SB_CARRY add_4439_5 (.CI(n36006), .I0(n8609[2]), .I1(n437_adj_3804), 
            .CO(n36007));
    SB_LUT4 add_4439_4_lut (.I0(GND_net), .I1(n8609[1]), .I2(n340), .I3(n36005), 
            .O(n8592[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_15 (.CI(n36973), .I0(n282[13]), .I1(n64[13]), 
            .CO(n36974));
    SB_LUT4 mult_14_add_1218_8_lut (.I0(GND_net), .I1(n1804[5]), .I2(n533), 
            .I3(n36893), .O(n1803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_17 (.CI(n36787), .I0(n1799[14]), .I1(GND_net), 
            .CO(n36788));
    SB_CARRY add_4470_3 (.CI(n36630), .I0(n9192[0]), .I1(n264_adj_3803), 
            .CO(n36631));
    SB_LUT4 add_4453_18_lut (.I0(GND_net), .I1(n8886[15]), .I2(GND_net), 
            .I3(n36373), .O(n8859[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_4 (.CI(n36005), .I0(n8609[1]), .I1(n340), .CO(n36006));
    SB_LUT4 add_4439_3_lut (.I0(GND_net), .I1(n8609[0]), .I2(n243_adj_3806), 
            .I3(n36004), .O(n8592[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_18 (.CI(n36373), .I0(n8886[15]), .I1(GND_net), .CO(n36374));
    SB_CARRY add_4439_3 (.CI(n36004), .I0(n8609[0]), .I1(n243_adj_3806), 
            .CO(n36005));
    SB_LUT4 add_4439_2_lut (.I0(GND_net), .I1(n53_adj_3807), .I2(n146_adj_3808), 
            .I3(GND_net), .O(n8592[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4439_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4470_2_lut (.I0(GND_net), .I1(n74_adj_3809), .I2(n167_adj_3810), 
            .I3(GND_net), .O(n9182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4470_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_17_lut (.I0(GND_net), .I1(n8886[14]), .I2(GND_net), 
            .I3(n36372), .O(n8859[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4439_2 (.CI(GND_net), .I0(n53_adj_3807), .I1(n146_adj_3808), 
            .CO(n36004));
    SB_LUT4 add_4438_17_lut (.I0(GND_net), .I1(n8592[14]), .I2(GND_net), 
            .I3(n36003), .O(n8574[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_17 (.CI(n36372), .I0(n8886[14]), .I1(GND_net), .CO(n36373));
    SB_LUT4 add_4438_16_lut (.I0(GND_net), .I1(n8592[13]), .I2(GND_net), 
            .I3(n36002), .O(n8574[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_16 (.CI(n36002), .I0(n8592[13]), .I1(GND_net), .CO(n36003));
    SB_LUT4 mult_14_add_1213_16_lut (.I0(GND_net), .I1(n1799[13]), .I2(GND_net), 
            .I3(n36786), .O(n1798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4470_2 (.CI(GND_net), .I0(n74_adj_3809), .I1(n167_adj_3810), 
            .CO(n36630));
    SB_LUT4 add_4453_16_lut (.I0(GND_net), .I1(n8886[13]), .I2(GND_net), 
            .I3(n36371), .O(n8859[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_15_lut (.I0(GND_net), .I1(n8592[12]), .I2(GND_net), 
            .I3(n36001), .O(n8574[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_15 (.CI(n36001), .I0(n8592[12]), .I1(GND_net), .CO(n36002));
    SB_CARRY add_4453_16 (.CI(n36371), .I0(n8886[13]), .I1(GND_net), .CO(n36372));
    SB_LUT4 add_4438_14_lut (.I0(GND_net), .I1(n8592[11]), .I2(GND_net), 
            .I3(n36000), .O(n8574[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_14 (.CI(n36000), .I0(n8592[11]), .I1(GND_net), .CO(n36001));
    SB_LUT4 add_4469_10_lut (.I0(GND_net), .I1(n9182[7]), .I2(GND_net), 
            .I3(n36629), .O(n9171[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_15_lut (.I0(GND_net), .I1(n8886[12]), .I2(GND_net), 
            .I3(n36370), .O(n8859[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_13_lut (.I0(GND_net), .I1(n8592[10]), .I2(GND_net), 
            .I3(n35999), .O(n8574[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_13 (.CI(n35999), .I0(n8592[10]), .I1(GND_net), .CO(n36000));
    SB_CARRY add_4453_15 (.CI(n36370), .I0(n8886[12]), .I1(GND_net), .CO(n36371));
    SB_LUT4 add_4438_12_lut (.I0(GND_net), .I1(n8592[9]), .I2(GND_net), 
            .I3(n35998), .O(n8574[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_12 (.CI(n35998), .I0(n8592[9]), .I1(GND_net), .CO(n35999));
    SB_CARRY mult_14_add_1218_8 (.CI(n36893), .I0(n1804[5]), .I1(n533), 
            .CO(n36894));
    SB_CARRY mult_14_add_1213_16 (.CI(n36786), .I0(n1799[13]), .I1(GND_net), 
            .CO(n36787));
    SB_LUT4 add_4469_9_lut (.I0(GND_net), .I1(n9182[6]), .I2(GND_net), 
            .I3(n36628), .O(n9171[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_14_lut (.I0(GND_net), .I1(n8886[11]), .I2(GND_net), 
            .I3(n36369), .O(n8859[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_11_lut (.I0(GND_net), .I1(n8592[8]), .I2(GND_net), 
            .I3(n35997), .O(n8574[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_11 (.CI(n35997), .I0(n8592[8]), .I1(GND_net), .CO(n35998));
    SB_CARRY add_4453_14 (.CI(n36369), .I0(n8886[11]), .I1(GND_net), .CO(n36370));
    SB_LUT4 add_4438_10_lut (.I0(GND_net), .I1(n8592[7]), .I2(GND_net), 
            .I3(n35996), .O(n8574[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_10 (.CI(n35996), .I0(n8592[7]), .I1(GND_net), .CO(n35997));
    SB_CARRY add_4469_9 (.CI(n36628), .I0(n9182[6]), .I1(GND_net), .CO(n36629));
    SB_LUT4 add_4453_13_lut (.I0(GND_net), .I1(n8886[10]), .I2(GND_net), 
            .I3(n36368), .O(n8859[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_9_lut (.I0(GND_net), .I1(n8592[6]), .I2(GND_net), 
            .I3(n35995), .O(n8574[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_9 (.CI(n35995), .I0(n8592[6]), .I1(GND_net), .CO(n35996));
    SB_CARRY add_4453_13 (.CI(n36368), .I0(n8886[10]), .I1(GND_net), .CO(n36369));
    SB_LUT4 add_4438_8_lut (.I0(GND_net), .I1(n8592[5]), .I2(n725_adj_3811), 
            .I3(n35994), .O(n8574[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_8 (.CI(n35994), .I0(n8592[5]), .I1(n725_adj_3811), 
            .CO(n35995));
    SB_LUT4 mult_14_add_1213_15_lut (.I0(GND_net), .I1(n1799[12]), .I2(GND_net), 
            .I3(n36785), .O(n1798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4469_8_lut (.I0(GND_net), .I1(n9182[5]), .I2(n746_adj_3812), 
            .I3(n36627), .O(n9171[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_12_lut (.I0(GND_net), .I1(n8886[9]), .I2(GND_net), 
            .I3(n36367), .O(n8859[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_7_lut (.I0(GND_net), .I1(n8592[4]), .I2(n628_adj_3813), 
            .I3(n35993), .O(n8574[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_7 (.CI(n35993), .I0(n8592[4]), .I1(n628_adj_3813), 
            .CO(n35994));
    SB_CARRY add_4453_12 (.CI(n36367), .I0(n8886[9]), .I1(GND_net), .CO(n36368));
    SB_LUT4 add_4438_6_lut (.I0(GND_net), .I1(n8592[3]), .I2(n531_adj_3814), 
            .I3(n35992), .O(n8574[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_6 (.CI(n35992), .I0(n8592[3]), .I1(n531_adj_3814), 
            .CO(n35993));
    SB_CARRY add_4469_8 (.CI(n36627), .I0(n9182[5]), .I1(n746_adj_3812), 
            .CO(n36628));
    SB_LUT4 add_4453_11_lut (.I0(GND_net), .I1(n8886[8]), .I2(GND_net), 
            .I3(n36366), .O(n8859[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_5_lut (.I0(GND_net), .I1(n8592[2]), .I2(n434_adj_3815), 
            .I3(n35991), .O(n8574[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_5 (.CI(n35991), .I0(n8592[2]), .I1(n434_adj_3815), 
            .CO(n35992));
    SB_CARRY add_4453_11 (.CI(n36366), .I0(n8886[8]), .I1(GND_net), .CO(n36367));
    SB_LUT4 add_4438_4_lut (.I0(GND_net), .I1(n8592[1]), .I2(n337_adj_3816), 
            .I3(n35990), .O(n8574[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_4 (.CI(n35990), .I0(n8592[1]), .I1(n337_adj_3816), 
            .CO(n35991));
    SB_LUT4 add_13_add_1_28678_add_1_14_lut (.I0(GND_net), .I1(n282[12]), 
            .I2(n64[12]), .I3(n36972), .O(n66[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_7_lut (.I0(GND_net), .I1(n1804[4]), .I2(n460_adj_3819), 
            .I3(n36892), .O(n1803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_15 (.CI(n36785), .I0(n1799[12]), .I1(GND_net), 
            .CO(n36786));
    SB_LUT4 add_4469_7_lut (.I0(GND_net), .I1(n9182[4]), .I2(n649_adj_3820), 
            .I3(n36626), .O(n9171[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_10_lut (.I0(GND_net), .I1(n8886[7]), .I2(GND_net), 
            .I3(n36365), .O(n8859[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4438_3_lut (.I0(GND_net), .I1(n8592[0]), .I2(n240_adj_3821), 
            .I3(n35989), .O(n8574[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_3 (.CI(n35989), .I0(n8592[0]), .I1(n240_adj_3821), 
            .CO(n35990));
    SB_CARRY add_4453_10 (.CI(n36365), .I0(n8886[7]), .I1(GND_net), .CO(n36366));
    SB_LUT4 add_4438_2_lut (.I0(GND_net), .I1(n50_adj_3822), .I2(n143_adj_3823), 
            .I3(GND_net), .O(n8574[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4438_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4438_2 (.CI(GND_net), .I0(n50_adj_3822), .I1(n143_adj_3823), 
            .CO(n35989));
    SB_CARRY add_4469_7 (.CI(n36626), .I0(n9182[4]), .I1(n649_adj_3820), 
            .CO(n36627));
    SB_LUT4 add_4453_9_lut (.I0(GND_net), .I1(n8886[6]), .I2(GND_net), 
            .I3(n36364), .O(n8859[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_18_lut (.I0(GND_net), .I1(n8574[15]), .I2(GND_net), 
            .I3(n35988), .O(n8555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_17_lut (.I0(GND_net), .I1(n8574[14]), .I2(GND_net), 
            .I3(n35987), .O(n8555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_9 (.CI(n36364), .I0(n8886[6]), .I1(GND_net), .CO(n36365));
    SB_CARRY add_4437_17 (.CI(n35987), .I0(n8574[14]), .I1(GND_net), .CO(n35988));
    SB_LUT4 add_4437_16_lut (.I0(GND_net), .I1(n8574[13]), .I2(GND_net), 
            .I3(n35986), .O(n8555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_14_lut (.I0(GND_net), .I1(n1799[11]), .I2(GND_net), 
            .I3(n36784), .O(n1798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4469_6_lut (.I0(GND_net), .I1(n9182[3]), .I2(n552_adj_3824), 
            .I3(n36625), .O(n9171[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_8_lut (.I0(GND_net), .I1(n8886[5]), .I2(n698_adj_3825), 
            .I3(n36363), .O(n8859[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_16 (.CI(n35986), .I0(n8574[13]), .I1(GND_net), .CO(n35987));
    SB_LUT4 add_4437_15_lut (.I0(GND_net), .I1(n8574[12]), .I2(GND_net), 
            .I3(n35985), .O(n8555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_11 (.CI(n34608), .I0(\PID_CONTROLLER.err_prev[9] ), 
            .I1(n60[9]), .CO(n34609));
    SB_LUT4 sub_11_add_2_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[8] ), 
            .I2(n60[8]), .I3(n34607), .O(n58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4469_6 (.CI(n36625), .I0(n9182[3]), .I1(n552_adj_3824), 
            .CO(n36626));
    SB_CARRY add_4437_15 (.CI(n35985), .I0(n8574[12]), .I1(GND_net), .CO(n35986));
    SB_CARRY add_4453_8 (.CI(n36363), .I0(n8886[5]), .I1(n698_adj_3825), 
            .CO(n36364));
    SB_CARRY add_13_add_1_28678_add_1_14 (.CI(n36972), .I0(n282[12]), .I1(n64[12]), 
            .CO(n36973));
    SB_CARRY sub_11_add_2_10 (.CI(n34607), .I0(\PID_CONTROLLER.err_prev[8] ), 
            .I1(n60[8]), .CO(n34608));
    SB_LUT4 add_4469_5_lut (.I0(GND_net), .I1(n9182[2]), .I2(n455_adj_3827), 
            .I3(n36624), .O(n9171[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_14_lut (.I0(GND_net), .I1(n8574[11]), .I2(GND_net), 
            .I3(n35984), .O(n8555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_14 (.CI(n36784), .I0(n1799[11]), .I1(GND_net), 
            .CO(n36785));
    SB_CARRY add_4437_14 (.CI(n35984), .I0(n8574[11]), .I1(GND_net), .CO(n35985));
    SB_LUT4 sub_11_add_2_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[7] ), 
            .I2(n60[7]), .I3(n34606), .O(n58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_9 (.CI(n34606), .I0(\PID_CONTROLLER.err_prev[7] ), 
            .I1(n60[7]), .CO(n34607));
    SB_LUT4 mult_14_add_1213_13_lut (.I0(GND_net), .I1(n1799[10]), .I2(GND_net), 
            .I3(n36783), .O(n1798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[6] ), 
            .I2(n60[6]), .I3(n34605), .O(n58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n61[6]), 
            .I3(n34701), .O(n414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_7 (.CI(n36892), .I0(n1804[4]), .I1(n460_adj_3819), 
            .CO(n36893));
    SB_CARRY mult_14_add_1213_13 (.CI(n36783), .I0(n1799[10]), .I1(GND_net), 
            .CO(n36784));
    SB_CARRY add_4469_5 (.CI(n36624), .I0(n9182[2]), .I1(n455_adj_3827), 
            .CO(n36625));
    SB_CARRY sub_11_add_2_8 (.CI(n34605), .I0(\PID_CONTROLLER.err_prev[6] ), 
            .I1(n60[6]), .CO(n34606));
    SB_LUT4 add_4469_4_lut (.I0(GND_net), .I1(n9182[1]), .I2(n358_adj_3830), 
            .I3(n36623), .O(n9171[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_7_lut (.I0(GND_net), .I1(n8886[4]), .I2(n601_adj_3831), 
            .I3(n36362), .O(n8859[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4469_4 (.CI(n36623), .I0(n9182[1]), .I1(n358_adj_3830), 
            .CO(n36624));
    SB_CARRY unary_minus_21_add_3_8 (.CI(n34701), .I0(GND_net), .I1(n61[6]), 
            .CO(n34702));
    SB_LUT4 mult_14_add_1213_12_lut (.I0(GND_net), .I1(n1799[9]), .I2(GND_net), 
            .I3(n36782), .O(n1798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_13_lut (.I0(GND_net), .I1(n8574[10]), .I2(GND_net), 
            .I3(n35983), .O(n8555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n61[5]), 
            .I3(n34700), .O(n67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_13_lut (.I0(GND_net), .I1(n282[11]), 
            .I2(n64[11]), .I3(n36971), .O(n66[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_6_lut (.I0(GND_net), .I1(n1804[3]), .I2(n387_adj_3833), 
            .I3(n36891), .O(n1803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_13 (.CI(n35983), .I0(n8574[10]), .I1(GND_net), .CO(n35984));
    SB_LUT4 sub_11_add_2_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[5] ), 
            .I2(n60[5]), .I3(n34604), .O(n58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_13 (.CI(n36971), .I0(n282[11]), .I1(n64[11]), 
            .CO(n36972));
    SB_CARRY add_4453_7 (.CI(n36362), .I0(n8886[4]), .I1(n601_adj_3831), 
            .CO(n36363));
    SB_LUT4 add_4469_3_lut (.I0(GND_net), .I1(n9182[0]), .I2(n261_adj_3835), 
            .I3(n36622), .O(n9171[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_12_lut (.I0(GND_net), .I1(n8574[9]), .I2(GND_net), 
            .I3(n35982), .O(n8555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_7 (.CI(n34604), .I0(\PID_CONTROLLER.err_prev[5] ), 
            .I1(n60[5]), .CO(n34605));
    SB_CARRY mult_14_add_1218_6 (.CI(n36891), .I0(n1804[3]), .I1(n387_adj_3833), 
            .CO(n36892));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n34700), .I0(GND_net), .I1(n61[5]), 
            .CO(n34701));
    SB_CARRY mult_14_add_1213_12 (.CI(n36782), .I0(n1799[9]), .I1(GND_net), 
            .CO(n36783));
    SB_CARRY add_4469_3 (.CI(n36622), .I0(n9182[0]), .I1(n261_adj_3835), 
            .CO(n36623));
    SB_LUT4 add_4453_6_lut (.I0(GND_net), .I1(n8886[3]), .I2(n504_adj_3836), 
            .I3(n36361), .O(n8859[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_6 (.CI(n36361), .I0(n8886[3]), .I1(n504_adj_3836), 
            .CO(n36362));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n61[4]), 
            .I3(n34699), .O(n416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_12 (.CI(n35982), .I0(n8574[9]), .I1(GND_net), .CO(n35983));
    SB_LUT4 add_4453_5_lut (.I0(GND_net), .I1(n8886[2]), .I2(n407_adj_3837), 
            .I3(n36360), .O(n8859[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_5 (.CI(n36360), .I0(n8886[2]), .I1(n407_adj_3837), 
            .CO(n36361));
    SB_LUT4 add_4437_11_lut (.I0(GND_net), .I1(n8574[8]), .I2(GND_net), 
            .I3(n35981), .O(n8555[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_11 (.CI(n35981), .I0(n8574[8]), .I1(GND_net), .CO(n35982));
    SB_LUT4 add_4437_10_lut (.I0(GND_net), .I1(n8574[7]), .I2(GND_net), 
            .I3(n35980), .O(n8555[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4469_2_lut (.I0(GND_net), .I1(n71_adj_3838), .I2(n164_adj_3839), 
            .I3(GND_net), .O(n9171[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4469_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4453_4_lut (.I0(GND_net), .I1(n8886[1]), .I2(n310_adj_3840), 
            .I3(n36359), .O(n8859[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_10 (.CI(n35980), .I0(n8574[7]), .I1(GND_net), .CO(n35981));
    SB_LUT4 add_4437_9_lut (.I0(GND_net), .I1(n8574[6]), .I2(GND_net), 
            .I3(n35979), .O(n8555[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[4] ), 
            .I2(n60[4]), .I3(n34603), .O(n58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_6 (.CI(n34603), .I0(\PID_CONTROLLER.err_prev[4] ), 
            .I1(n60[4]), .CO(n34604));
    SB_CARRY unary_minus_21_add_3_6 (.CI(n34699), .I0(GND_net), .I1(n61[4]), 
            .CO(n34700));
    SB_CARRY add_4469_2 (.CI(GND_net), .I0(n71_adj_3838), .I1(n164_adj_3839), 
            .CO(n36622));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n61[3]), 
            .I3(n34698), .O(n67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_9 (.CI(n35979), .I0(n8574[6]), .I1(GND_net), .CO(n35980));
    SB_LUT4 add_4468_11_lut (.I0(GND_net), .I1(n9171[8]), .I2(GND_net), 
            .I3(n36621), .O(n9159[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(n41825));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_4437_8_lut (.I0(GND_net), .I1(n8574[5]), .I2(n722_adj_3842), 
            .I3(n35978), .O(n8555[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_4 (.CI(n36359), .I0(n8886[1]), .I1(n310_adj_3840), 
            .CO(n36360));
    SB_LUT4 sub_11_add_2_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[3] ), 
            .I2(n60[3]), .I3(n34602), .O(n58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_8 (.CI(n35978), .I0(n8574[5]), .I1(n722_adj_3842), 
            .CO(n35979));
    SB_LUT4 add_13_add_1_28678_add_1_12_lut (.I0(GND_net), .I1(n282[10]), 
            .I2(n64[10]), .I3(n36970), .O(n66[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_5 (.CI(n34602), .I0(\PID_CONTROLLER.err_prev[3] ), 
            .I1(n60[3]), .CO(n34603));
    SB_LUT4 mult_14_add_1218_5_lut (.I0(GND_net), .I1(n1804[2]), .I2(n314_adj_3845), 
            .I3(n36890), .O(n1803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_11_lut (.I0(GND_net), .I1(n1799[8]), .I2(GND_net), 
            .I3(n36781), .O(n1798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_12 (.CI(n36970), .I0(n282[10]), .I1(n64[10]), 
            .CO(n36971));
    SB_CARRY mult_14_add_1213_11 (.CI(n36781), .I0(n1799[8]), .I1(GND_net), 
            .CO(n36782));
    SB_LUT4 add_4468_10_lut (.I0(GND_net), .I1(n9171[7]), .I2(GND_net), 
            .I3(n36620), .O(n9159[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_10_lut (.I0(GND_net), .I1(n1799[7]), .I2(GND_net), 
            .I3(n36780), .O(n1798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n34698), .I0(GND_net), .I1(n61[3]), 
            .CO(n34699));
    SB_LUT4 add_4453_3_lut (.I0(GND_net), .I1(n8886[0]), .I2(n213_adj_3846), 
            .I3(n36358), .O(n8859[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4437_7_lut (.I0(GND_net), .I1(n8574[4]), .I2(n625_adj_3847), 
            .I3(n35977), .O(n8555[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n61[2]), 
            .I3(n34697), .O(n67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_11_lut (.I0(GND_net), .I1(n282[9]), 
            .I2(n64[9]), .I3(n36969), .O(n66[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_10 (.CI(n36620), .I0(n9171[7]), .I1(GND_net), .CO(n36621));
    SB_CARRY mult_14_add_1213_10 (.CI(n36780), .I0(n1799[7]), .I1(GND_net), 
            .CO(n36781));
    SB_LUT4 sub_11_add_2_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[2] ), 
            .I2(n60[2]), .I3(n34601), .O(n58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_7 (.CI(n35977), .I0(n8574[4]), .I1(n625_adj_3847), 
            .CO(n35978));
    SB_CARRY add_13_add_1_28678_add_1_11 (.CI(n36969), .I0(n282[9]), .I1(n64[9]), 
            .CO(n36970));
    SB_CARRY sub_11_add_2_4 (.CI(n34601), .I0(\PID_CONTROLLER.err_prev[2] ), 
            .I1(n60[2]), .CO(n34602));
    SB_LUT4 add_4437_6_lut (.I0(GND_net), .I1(n8574[3]), .I2(n528_adj_3849), 
            .I3(n35976), .O(n8555[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_5 (.CI(n36890), .I0(n1804[2]), .I1(n314_adj_3845), 
            .CO(n36891));
    SB_LUT4 mult_14_add_1218_4_lut (.I0(GND_net), .I1(n1804[1]), .I2(n241_adj_3851), 
            .I3(n36889), .O(n1803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_4 (.CI(n36889), .I0(n1804[1]), .I1(n241_adj_3851), 
            .CO(n36890));
    SB_LUT4 sub_11_add_2_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[1] ), 
            .I2(n60[1]), .I3(n34600), .O(n58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_10_lut (.I0(GND_net), .I1(n282[8]), 
            .I2(n64[8]), .I3(n36968), .O(n66[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_3 (.CI(n36358), .I0(n8886[0]), .I1(n213_adj_3846), 
            .CO(n36359));
    SB_CARRY add_4437_6 (.CI(n35976), .I0(n8574[3]), .I1(n528_adj_3849), 
            .CO(n35977));
    SB_LUT4 i5_4_lut_adj_845 (.I0(n48474), .I1(pwm[21]), .I2(pwm[8]), 
            .I3(pwm_count[8]), .O(n20_adj_3853));
    defparam i5_4_lut_adj_845.LUT_INIT = 16'hecfe;
    SB_LUT4 i11_4_lut (.I0(pwm[11]), .I1(pwm[17]), .I2(pwm[19]), .I3(pwm[12]), 
            .O(n26_adj_3854));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(pwm[14]), .I1(pwm[10]), .I2(pwm[16]), .I3(pwm[9]), 
            .O(n24_adj_3855));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(pwm[13]), .I1(n26_adj_3854), .I2(n20_adj_3853), 
            .I3(pwm[22]), .O(n28_adj_3856));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(pwm[15]), .I1(pwm[18]), .I2(pwm[20]), .I3(GND_net), 
            .O(n23_adj_3857));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mult_14_add_1218_3_lut (.I0(GND_net), .I1(n1804[0]), .I2(n168_adj_3859), 
            .I3(n36888), .O(n1803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_846 (.I0(pwm[23]), .I1(n23_adj_3857), .I2(n28_adj_3856), 
            .I3(n24_adj_3855), .O(n17_adj_3860));   // verilog/motorControl.v(65[9:32])
    defparam i1_4_lut_adj_846.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_21_add_3_4 (.CI(n34697), .I0(GND_net), .I1(n61[2]), 
            .CO(n34698));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n61[1]), 
            .I3(n34696), .O(n67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_3 (.CI(n34600), .I0(\PID_CONTROLLER.err_prev[1] ), 
            .I1(n60[1]), .CO(n34601));
    SB_LUT4 add_4453_2_lut (.I0(GND_net), .I1(n23_adj_3861), .I2(n116_adj_3862), 
            .I3(GND_net), .O(n8859[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4453_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_10 (.CI(n36968), .I0(n282[8]), .I1(n64[8]), 
            .CO(n36969));
    SB_CARRY mult_14_add_1218_3 (.CI(n36888), .I0(n1804[0]), .I1(n168_adj_3859), 
            .CO(n36889));
    SB_LUT4 mult_14_add_1218_2_lut (.I0(GND_net), .I1(n26_adj_3863), .I2(n95), 
            .I3(GND_net), .O(n1803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4453_2 (.CI(GND_net), .I0(n23_adj_3861), .I1(n116_adj_3862), 
            .CO(n36358));
    SB_LUT4 add_4437_5_lut (.I0(GND_net), .I1(n8574[2]), .I2(n431_adj_3864), 
            .I3(n35975), .O(n8555[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n34696), .I0(GND_net), .I1(n61[1]), 
            .CO(n34697));
    SB_CARRY mult_14_add_1218_2 (.CI(GND_net), .I0(n26_adj_3863), .I1(n95), 
            .CO(n36888));
    SB_LUT4 sub_11_add_2_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[0] ), 
            .I2(n60[0]), .I3(VCC_net), .O(n58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n25957), .I1(GND_net), .I2(n61[0]), 
            .I3(VCC_net), .O(n46522)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_14_add_1213_9_lut (.I0(GND_net), .I1(n1799[6]), .I2(GND_net), 
            .I3(n36779), .O(n1798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_24_lut (.I0(GND_net), .I1(n1803[21]), .I2(GND_net), 
            .I3(n36886), .O(n1802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_9_lut (.I0(GND_net), .I1(n282[7]), 
            .I2(n64[7]), .I3(n36967), .O(n66[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_5 (.CI(n35975), .I0(n8574[2]), .I1(n431_adj_3864), 
            .CO(n35976));
    SB_LUT4 add_4437_4_lut (.I0(GND_net), .I1(n8574[1]), .I2(n334_adj_3867), 
            .I3(n35974), .O(n8555[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_4 (.CI(n35974), .I0(n8574[1]), .I1(n334_adj_3867), 
            .CO(n35975));
    SB_CARRY add_13_add_1_28678_add_1_9 (.CI(n36967), .I0(n282[7]), .I1(n64[7]), 
            .CO(n36968));
    SB_CARRY sub_11_add_2_2 (.CI(VCC_net), .I0(\PID_CONTROLLER.err_prev[0] ), 
            .I1(n60[0]), .CO(n34600));
    SB_LUT4 add_13_add_1_28678_add_1_8_lut (.I0(GND_net), .I1(n282[6]), 
            .I2(n64[6]), .I3(n36966), .O(n66[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_8 (.CI(n36966), .I0(n282[6]), .I1(n64[6]), 
            .CO(n36967));
    SB_CARRY mult_14_add_1217_24 (.CI(n36886), .I0(n1803[21]), .I1(GND_net), 
            .CO(n1707));
    SB_CARRY mult_14_add_1213_9 (.CI(n36779), .I0(n1799[6]), .I1(GND_net), 
            .CO(n36780));
    SB_LUT4 mult_14_add_1213_8_lut (.I0(GND_net), .I1(n1799[5]), .I2(n518), 
            .I3(n36778), .O(n1798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_8 (.CI(n36778), .I0(n1799[5]), .I1(n518), 
            .CO(n36779));
    SB_LUT4 mult_14_add_1213_7_lut (.I0(GND_net), .I1(n1799[4]), .I2(n445), 
            .I3(n36777), .O(n1798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4468_9_lut (.I0(GND_net), .I1(n9171[6]), .I2(GND_net), 
            .I3(n36619), .O(n9159[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_7_lut (.I0(GND_net), .I1(n282[5]), 
            .I2(n64[5]), .I3(n36965), .O(n66[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n61[0]), 
            .CO(n34696));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n76[23]), 
            .I3(n34695), .O(n75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_9 (.CI(n36619), .I0(n9171[6]), .I1(GND_net), .CO(n36620));
    SB_CARRY add_13_add_1_28678_add_1_7 (.CI(n36965), .I0(n282[5]), .I1(n64[5]), 
            .CO(n36966));
    SB_LUT4 add_4437_3_lut (.I0(GND_net), .I1(n8574[0]), .I2(n237_adj_3872), 
            .I3(n35973), .O(n8555[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4468_8_lut (.I0(GND_net), .I1(n9171[5]), .I2(n743_adj_3873), 
            .I3(n36618), .O(n9159[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4437_3 (.CI(n35973), .I0(n8574[0]), .I1(n237_adj_3872), 
            .CO(n35974));
    SB_LUT4 add_4437_2_lut (.I0(GND_net), .I1(n47_adj_3874), .I2(n140_adj_3875), 
            .I3(GND_net), .O(n8555[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4437_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_23_lut (.I0(GND_net), .I1(n1803[20]), .I2(GND_net), 
            .I3(n36885), .O(n1802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_7 (.CI(n36777), .I0(n1799[4]), .I1(n445), 
            .CO(n36778));
    SB_LUT4 mult_14_add_1213_6_lut (.I0(GND_net), .I1(n1799[3]), .I2(n372), 
            .I3(n36776), .O(n1798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4452_27_lut (.I0(GND_net), .I1(n8859[24]), .I2(GND_net), 
            .I3(n36357), .O(n8831[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[22]), .I3(n34694), .O(n45_adj_3877)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4437_2 (.CI(GND_net), .I0(n47_adj_3874), .I1(n140_adj_3875), 
            .CO(n35973));
    SB_CARRY add_4468_8 (.CI(n36618), .I0(n9171[5]), .I1(n743_adj_3873), 
            .CO(n36619));
    SB_LUT4 add_4452_26_lut (.I0(GND_net), .I1(n8859[23]), .I2(GND_net), 
            .I3(n36356), .O(n8831[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_26 (.CI(n36356), .I0(n8859[23]), .I1(GND_net), .CO(n36357));
    SB_CARRY unary_minus_5_add_3_24 (.CI(n34694), .I0(GND_net), .I1(n76[22]), 
            .CO(n34695));
    SB_LUT4 add_4468_7_lut (.I0(GND_net), .I1(n9171[4]), .I2(n646_adj_3879), 
            .I3(n36617), .O(n9159[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i73_4_lut (.I0(pwm[23]), .I1(n25), .I2(n30), .I3(n26), .O(n878));   // verilog/motorControl.v(86[19:44])
    defparam i73_4_lut.LUT_INIT = 16'haaa8;
    SB_DFF \PID_CONTROLLER.result_i1  (.Q(\PID_CONTROLLER.result [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_4452_25_lut (.I0(GND_net), .I1(n8859[22]), .I2(GND_net), 
            .I3(n36355), .O(n8831[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_847 (.I0(hall3), .I1(n878), .I2(GND_net), .I3(GND_net), 
            .O(n41830));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h4444;
    SB_LUT4 add_4436_19_lut (.I0(GND_net), .I1(n8555[16]), .I2(GND_net), 
            .I3(n35972), .O(n8535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34686_2_lut (.I0(hall2), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n42569));
    defparam i34686_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i38786_3_lut (.I0(n41830), .I1(hall1), .I2(hall2), .I3(GND_net), 
            .O(n46668));   // verilog/motorControl.v(86[14] 109[8])
    defparam i38786_3_lut.LUT_INIT = 16'h8080;
    SB_DFF \PID_CONTROLLER.result_i2  (.Q(\PID_CONTROLLER.result [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i3  (.Q(\PID_CONTROLLER.result [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i4  (.Q(\PID_CONTROLLER.result[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i5  (.Q(\PID_CONTROLLER.result [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i6  (.Q(\PID_CONTROLLER.result[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i7  (.Q(\PID_CONTROLLER.result [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i8  (.Q(\PID_CONTROLLER.result [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i9  (.Q(\PID_CONTROLLER.result [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i10  (.Q(\PID_CONTROLLER.result[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i11  (.Q(\PID_CONTROLLER.result [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i12  (.Q(\PID_CONTROLLER.result [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i13  (.Q(\PID_CONTROLLER.result[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i14  (.Q(\PID_CONTROLLER.result [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i15  (.Q(\PID_CONTROLLER.result [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i16  (.Q(\PID_CONTROLLER.result [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i17  (.Q(\PID_CONTROLLER.result[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i18  (.Q(\PID_CONTROLLER.result [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i19  (.Q(\PID_CONTROLLER.result[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i20  (.Q(\PID_CONTROLLER.result [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i21  (.Q(\PID_CONTROLLER.result [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i22  (.Q(\PID_CONTROLLER.result [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i23  (.Q(\PID_CONTROLLER.result [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i24  (.Q(\PID_CONTROLLER.result [24]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i25  (.Q(\PID_CONTROLLER.result [25]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [25]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i26  (.Q(\PID_CONTROLLER.result [26]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [26]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i27  (.Q(\PID_CONTROLLER.result [27]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [27]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i28  (.Q(\PID_CONTROLLER.result [28]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [28]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i29  (.Q(\PID_CONTROLLER.result [29]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [29]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i30  (.Q(\PID_CONTROLLER.result [30]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [30]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i31  (.Q(\PID_CONTROLLER.result [31]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3353 [31]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err[1] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF GATES_i3 (.Q(PIN_8_c_2), .C(clk32MHz), .D(GATES_5__N_3138[2]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i4 (.Q(PIN_9_c_3), .C(clk32MHz), .D(GATES_5__N_3138[3]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i5 (.Q(PIN_10_c_4), .C(clk32MHz), .D(GATES_5__N_3138[4]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i6 (.Q(PIN_11_c_5), .C(clk32MHz), .D(GATES_5__N_3138[5]));   // verilog/motorControl.v(64[10] 111[6])
    SB_LUT4 add_4436_18_lut (.I0(GND_net), .I1(n8555[15]), .I2(GND_net), 
            .I3(n35971), .O(n8535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_6 (.CI(n36776), .I0(n1799[3]), .I1(n372), 
            .CO(n36777));
    SB_LUT4 i34_4_lut (.I0(n46668), .I1(n42569), .I2(n17_adj_3860), .I3(n41825), 
            .O(n18_adj_3883));   // verilog/motorControl.v(86[14] 109[8])
    defparam i34_4_lut.LUT_INIT = 16'ha3a0;
    SB_CARRY add_4436_18 (.CI(n35971), .I0(n8555[15]), .I1(GND_net), .CO(n35972));
    SB_LUT4 add_13_add_1_28678_add_1_6_lut (.I0(GND_net), .I1(n282[4]), 
            .I2(n64[4]), .I3(n36964), .O(n66[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_7 (.CI(n36617), .I0(n9171[4]), .I1(n646_adj_3879), 
            .CO(n36618));
    SB_LUT4 add_4468_6_lut (.I0(GND_net), .I1(n9171[3]), .I2(n549_adj_3884), 
            .I3(n36616), .O(n9159[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_5_lut (.I0(GND_net), .I1(n1799[2]), .I2(n299_adj_3886), 
            .I3(n36775), .O(n1798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_6 (.CI(n36616), .I0(n9171[3]), .I1(n549_adj_3884), 
            .CO(n36617));
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err[2] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_4452_25 (.CI(n36355), .I0(n8859[22]), .I1(GND_net), .CO(n36356));
    SB_CARRY mult_14_add_1213_5 (.CI(n36775), .I0(n1799[2]), .I1(n299_adj_3886), 
            .CO(n36776));
    SB_LUT4 add_4468_5_lut (.I0(GND_net), .I1(n9171[2]), .I2(n452_adj_3887), 
            .I3(n36615), .O(n9159[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_23 (.CI(n36885), .I0(n1803[20]), .I1(GND_net), 
            .CO(n36886));
    SB_LUT4 mult_14_add_1213_4_lut (.I0(GND_net), .I1(n1799[1]), .I2(n226_adj_3889), 
            .I3(n36774), .O(n1798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_24_lut (.I0(GND_net), .I1(n8859[21]), .I2(GND_net), 
            .I3(n36354), .O(n8831[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_4 (.CI(n36774), .I0(n1799[1]), .I1(n226_adj_3889), 
            .CO(n36775));
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err[3] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err[8] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err[9] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err[11] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err[12] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err[15] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err[16] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err[18] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err[22] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i24  (.Q(\PID_CONTROLLER.err[23] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i25  (.Q(\PID_CONTROLLER.err[31] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_3175 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 i33_4_lut (.I0(n18_adj_3883), .I1(n17_adj_3860), .I2(\GATES_5__N_3398[5] ), 
            .I3(n41830), .O(GATES_5__N_3138[1]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i33_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_4468_5 (.CI(n36615), .I0(n9171[2]), .I1(n452_adj_3887), 
            .CO(n36616));
    SB_LUT4 add_4436_17_lut (.I0(GND_net), .I1(n8555[14]), .I2(GND_net), 
            .I3(n35970), .O(n8535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_6 (.CI(n36964), .I0(n282[4]), .I1(n64[4]), 
            .CO(n36965));
    SB_LUT4 mult_14_add_1217_22_lut (.I0(GND_net), .I1(n1803[19]), .I2(GND_net), 
            .I3(n36884), .O(n1802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_22 (.CI(n36884), .I0(n1803[19]), .I1(GND_net), 
            .CO(n36885));
    SB_LUT4 mult_14_i144_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3549));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_28678_add_1_5_lut (.I0(GND_net), .I1(n282[3]), 
            .I2(n64[3]), .I3(n36963), .O(n66[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[21]), .I3(n34693), .O(n43_adj_3890)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1217_21_lut (.I0(GND_net), .I1(n1803[18]), .I2(GND_net), 
            .I3(n36883), .O(n1802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_3_lut (.I0(GND_net), .I1(n1799[0]), .I2(n153_adj_3893), 
            .I3(n36773), .O(n1798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4468_4_lut (.I0(GND_net), .I1(n9171[1]), .I2(n355_adj_3894), 
            .I3(n36614), .O(n9159[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_3 (.CI(n36773), .I0(n1799[0]), .I1(n153_adj_3893), 
            .CO(n36774));
    SB_CARRY add_4452_24 (.CI(n36354), .I0(n8859[21]), .I1(GND_net), .CO(n36355));
    SB_LUT4 add_4452_23_lut (.I0(GND_net), .I1(n8859[20]), .I2(GND_net), 
            .I3(n36353), .O(n8831[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_4 (.CI(n36614), .I0(n9171[1]), .I1(n355_adj_3894), 
            .CO(n36615));
    SB_CARRY add_4452_23 (.CI(n36353), .I0(n8859[20]), .I1(GND_net), .CO(n36354));
    SB_LUT4 add_4452_22_lut (.I0(GND_net), .I1(n8859[19]), .I2(GND_net), 
            .I3(n36352), .O(n8831[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_21 (.CI(n36883), .I0(n1803[18]), .I1(GND_net), 
            .CO(n36884));
    SB_LUT4 mult_14_add_1213_2_lut (.I0(GND_net), .I1(n11_adj_3895), .I2(n80_adj_3896), 
            .I3(GND_net), .O(n1798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4468_3_lut (.I0(GND_net), .I1(n9171[0]), .I2(n258_adj_3897), 
            .I3(n36613), .O(n9159[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_22 (.CI(n36352), .I0(n8859[19]), .I1(GND_net), .CO(n36353));
    SB_LUT4 add_4452_21_lut (.I0(GND_net), .I1(n8859[18]), .I2(GND_net), 
            .I3(n36351), .O(n8831[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_3 (.CI(n36613), .I0(n9171[0]), .I1(n258_adj_3897), 
            .CO(n36614));
    SB_LUT4 mult_12_i353_2_lut (.I0(\Kd[5] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n525));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4452_21 (.CI(n36351), .I0(n8859[18]), .I1(GND_net), .CO(n36352));
    SB_LUT4 add_4452_20_lut (.I0(GND_net), .I1(n8859[17]), .I2(GND_net), 
            .I3(n36350), .O(n8831[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_5 (.CI(n36963), .I0(n282[3]), .I1(n64[3]), 
            .CO(n36964));
    SB_LUT4 mult_14_add_1217_20_lut (.I0(GND_net), .I1(n1803[17]), .I2(GND_net), 
            .I3(n36882), .O(n1802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_2 (.CI(GND_net), .I0(n11_adj_3895), .I1(n80_adj_3896), 
            .CO(n36773));
    SB_LUT4 add_4468_2_lut (.I0(GND_net), .I1(n68_adj_3898), .I2(n161_adj_3899), 
            .I3(GND_net), .O(n9159[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4468_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_20 (.CI(n36350), .I0(n8859[17]), .I1(GND_net), .CO(n36351));
    SB_LUT4 add_4452_19_lut (.I0(GND_net), .I1(n8859[16]), .I2(GND_net), 
            .I3(n36349), .O(n8831[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4468_2 (.CI(GND_net), .I0(n68_adj_3898), .I1(n161_adj_3899), 
            .CO(n36613));
    SB_CARRY add_4452_19 (.CI(n36349), .I0(n8859[16]), .I1(GND_net), .CO(n36350));
    SB_LUT4 add_4452_18_lut (.I0(GND_net), .I1(n8859[15]), .I2(GND_net), 
            .I3(n36348), .O(n8831[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_20 (.CI(n36882), .I0(n1803[17]), .I1(GND_net), 
            .CO(n36883));
    SB_LUT4 mult_14_add_1212_24_lut (.I0(GND_net), .I1(n1798[21]), .I2(GND_net), 
            .I3(n36771), .O(n1797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i193_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i193_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i418_2_lut (.I0(\Kd[6] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n622));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n34693), .I0(GND_net), .I1(n76[21]), 
            .CO(n34694));
    SB_CARRY mult_14_add_1212_24 (.CI(n36771), .I0(n1798[21]), .I1(GND_net), 
            .CO(n1687));
    SB_LUT4 mult_14_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4436_17 (.CI(n35970), .I0(n8555[14]), .I1(GND_net), .CO(n35971));
    SB_LUT4 add_4436_16_lut (.I0(GND_net), .I1(n8555[13]), .I2(GND_net), 
            .I3(n35969), .O(n8535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_16 (.CI(n35969), .I0(n8555[13]), .I1(GND_net), .CO(n35970));
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[2]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_13_add_1_28678_add_1_4_lut (.I0(GND_net), .I1(n282[2]), 
            .I2(n64[2]), .I3(n36962), .O(n66[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4467_12_lut (.I0(GND_net), .I1(n9159[9]), .I2(GND_net), 
            .I3(n36612), .O(n9146[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_18 (.CI(n36348), .I0(n8859[15]), .I1(GND_net), .CO(n36349));
    SB_LUT4 add_4452_17_lut (.I0(GND_net), .I1(n8859[14]), .I2(GND_net), 
            .I3(n36347), .O(n8831[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4467_11_lut (.I0(GND_net), .I1(n9159[8]), .I2(GND_net), 
            .I3(n36611), .O(n9146[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_17 (.CI(n36347), .I0(n8859[14]), .I1(GND_net), .CO(n36348));
    SB_CARRY add_13_add_1_28678_add_1_4 (.CI(n36962), .I0(n282[2]), .I1(n64[2]), 
            .CO(n36963));
    SB_LUT4 mult_14_add_1217_19_lut (.I0(GND_net), .I1(n1803[16]), .I2(GND_net), 
            .I3(n36881), .O(n1802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_23_lut (.I0(GND_net), .I1(n1798[20]), .I2(GND_net), 
            .I3(n36770), .O(n1797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_11 (.CI(n36611), .I0(n9159[8]), .I1(GND_net), .CO(n36612));
    SB_LUT4 add_4467_10_lut (.I0(GND_net), .I1(n9159[7]), .I2(GND_net), 
            .I3(n36610), .O(n9146[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_19 (.CI(n36881), .I0(n1803[16]), .I1(GND_net), 
            .CO(n36882));
    SB_LUT4 mult_12_i483_2_lut (.I0(\Kd[7] ), .I1(n58[13]), .I2(GND_net), 
            .I3(GND_net), .O(n719));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i483_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1212_23 (.CI(n36770), .I0(n1798[20]), .I1(GND_net), 
            .CO(n36771));
    SB_CARRY add_4467_10 (.CI(n36610), .I0(n9159[7]), .I1(GND_net), .CO(n36611));
    SB_LUT4 add_4467_9_lut (.I0(GND_net), .I1(n9159[6]), .I2(GND_net), 
            .I3(n36609), .O(n9146[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_3_lut (.I0(GND_net), .I1(n282[1]), 
            .I2(n64[1]), .I3(n36961), .O(n66[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_18_lut (.I0(GND_net), .I1(n1803[15]), .I2(GND_net), 
            .I3(n36880), .O(n1802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_22_lut (.I0(GND_net), .I1(n1798[19]), .I2(GND_net), 
            .I3(n36769), .O(n1797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_9 (.CI(n36609), .I0(n9159[6]), .I1(GND_net), .CO(n36610));
    SB_LUT4 add_4467_8_lut (.I0(GND_net), .I1(n9159[5]), .I2(n740_adj_3900), 
            .I3(n36608), .O(n9146[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_18 (.CI(n36880), .I0(n1803[15]), .I1(GND_net), 
            .CO(n36881));
    SB_CARRY mult_14_add_1212_22 (.CI(n36769), .I0(n1798[19]), .I1(GND_net), 
            .CO(n36770));
    SB_CARRY add_4467_8 (.CI(n36608), .I0(n9159[5]), .I1(n740_adj_3900), 
            .CO(n36609));
    SB_LUT4 add_4467_7_lut (.I0(GND_net), .I1(n9159[4]), .I2(n643_adj_3901), 
            .I3(n36607), .O(n9146[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_3 (.CI(n36961), .I0(n282[1]), .I1(n64[1]), 
            .CO(n36962));
    SB_LUT4 mult_14_add_1217_17_lut (.I0(GND_net), .I1(n1803[14]), .I2(GND_net), 
            .I3(n36879), .O(n1802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_21_lut (.I0(GND_net), .I1(n1798[18]), .I2(GND_net), 
            .I3(n36768), .O(n1797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_15_lut (.I0(GND_net), .I1(n8555[12]), .I2(GND_net), 
            .I3(n35968), .O(n8535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_7 (.CI(n36607), .I0(n9159[4]), .I1(n643_adj_3901), 
            .CO(n36608));
    SB_LUT4 add_4467_6_lut (.I0(GND_net), .I1(n9159[3]), .I2(n546_adj_3902), 
            .I3(n36606), .O(n9146[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_16_lut (.I0(GND_net), .I1(n8859[13]), .I2(GND_net), 
            .I3(n36346), .O(n8831[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_21 (.CI(n36768), .I0(n1798[18]), .I1(GND_net), 
            .CO(n36769));
    SB_CARRY add_4467_6 (.CI(n36606), .I0(n9159[3]), .I1(n546_adj_3902), 
            .CO(n36607));
    SB_LUT4 mult_14_i242_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i242_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3520));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4467_5_lut (.I0(GND_net), .I1(n9159[2]), .I2(n449_adj_3903), 
            .I3(n36605), .O(n9146[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_16 (.CI(n36346), .I0(n8859[13]), .I1(GND_net), .CO(n36347));
    SB_LUT4 add_4452_15_lut (.I0(GND_net), .I1(n8859[12]), .I2(GND_net), 
            .I3(n36345), .O(n8831[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_15 (.CI(n35968), .I0(n8555[12]), .I1(GND_net), .CO(n35969));
    SB_CARRY add_4452_15 (.CI(n36345), .I0(n8859[12]), .I1(GND_net), .CO(n36346));
    SB_LUT4 mult_14_add_1212_20_lut (.I0(GND_net), .I1(n1798[17]), .I2(GND_net), 
            .I3(n36767), .O(n1797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_5 (.CI(n36605), .I0(n9159[2]), .I1(n449_adj_3903), 
            .CO(n36606));
    SB_LUT4 add_4467_4_lut (.I0(GND_net), .I1(n9159[1]), .I2(n352_adj_3904), 
            .I3(n36604), .O(n9146[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_14_lut (.I0(GND_net), .I1(n8859[11]), .I2(GND_net), 
            .I3(n36344), .O(n8831[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[20]), .I3(n34692), .O(n41_adj_3905)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4452_14 (.CI(n36344), .I0(n8859[11]), .I1(GND_net), .CO(n36345));
    SB_LUT4 add_4436_14_lut (.I0(GND_net), .I1(n8555[11]), .I2(GND_net), 
            .I3(n35967), .O(n8535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_13_lut (.I0(GND_net), .I1(n8859[10]), .I2(GND_net), 
            .I3(n36343), .O(n8831[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_28678_add_1_2_lut (.I0(GND_net), .I1(n282[0]), 
            .I2(n64[0]), .I3(GND_net), .O(n66[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_28678_add_1_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_17 (.CI(n36879), .I0(n1803[14]), .I1(GND_net), 
            .CO(n36880));
    SB_CARRY add_4436_14 (.CI(n35967), .I0(n8555[11]), .I1(GND_net), .CO(n35968));
    SB_LUT4 add_4436_13_lut (.I0(GND_net), .I1(n8555[10]), .I2(GND_net), 
            .I3(n35966), .O(n8535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_16_lut (.I0(GND_net), .I1(n1803[13]), .I2(GND_net), 
            .I3(n36878), .O(n1802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_4 (.CI(n36604), .I0(n9159[1]), .I1(n352_adj_3904), 
            .CO(n36605));
    SB_CARRY add_4452_13 (.CI(n36343), .I0(n8859[10]), .I1(GND_net), .CO(n36344));
    SB_LUT4 add_4452_12_lut (.I0(GND_net), .I1(n8859[9]), .I2(GND_net), 
            .I3(n36342), .O(n8831[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_20 (.CI(n36767), .I0(n1798[17]), .I1(GND_net), 
            .CO(n36768));
    SB_CARRY add_4436_13 (.CI(n35966), .I0(n8555[10]), .I1(GND_net), .CO(n35967));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n34692), .I0(GND_net), .I1(n76[20]), 
            .CO(n34693));
    SB_LUT4 add_4436_12_lut (.I0(GND_net), .I1(n8555[9]), .I2(GND_net), 
            .I3(n35965), .O(n8535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_28678_add_1_2 (.CI(GND_net), .I0(n282[0]), .I1(n64[0]), 
            .CO(n36961));
    SB_LUT4 add_4467_3_lut (.I0(GND_net), .I1(n9159[0]), .I2(n255_adj_3909), 
            .I3(n36603), .O(n9146[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_12 (.CI(n36342), .I0(n8859[9]), .I1(GND_net), .CO(n36343));
    SB_CARRY add_4436_12 (.CI(n35965), .I0(n8555[9]), .I1(GND_net), .CO(n35966));
    SB_LUT4 add_4436_11_lut (.I0(GND_net), .I1(n8555[8]), .I2(GND_net), 
            .I3(n35964), .O(n8535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_11 (.CI(n35964), .I0(n8555[8]), .I1(GND_net), .CO(n35965));
    SB_LUT4 add_4436_10_lut (.I0(GND_net), .I1(n8555[7]), .I2(GND_net), 
            .I3(n35963), .O(n8535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_16 (.CI(n36878), .I0(n1803[13]), .I1(GND_net), 
            .CO(n36879));
    SB_LUT4 mult_14_add_1212_19_lut (.I0(GND_net), .I1(n1798[16]), .I2(GND_net), 
            .I3(n36766), .O(n1797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_15_lut (.I0(GND_net), .I1(n1803[12]), .I2(GND_net), 
            .I3(n36877), .O(n1802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4467_3 (.CI(n36603), .I0(n9159[0]), .I1(n255_adj_3909), 
            .CO(n36604));
    SB_LUT4 add_4452_11_lut (.I0(GND_net), .I1(n8859[8]), .I2(GND_net), 
            .I3(n36341), .O(n8831[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_11 (.CI(n36341), .I0(n8859[8]), .I1(GND_net), .CO(n36342));
    SB_LUT4 add_4467_2_lut (.I0(GND_net), .I1(n65_adj_3910), .I2(n158_adj_3911), 
            .I3(GND_net), .O(n9146[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4467_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_10_lut (.I0(GND_net), .I1(n8859[7]), .I2(GND_net), 
            .I3(n36340), .O(n8831[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_10 (.CI(n36340), .I0(n8859[7]), .I1(GND_net), .CO(n36341));
    SB_CARRY mult_14_add_1212_19 (.CI(n36766), .I0(n1798[16]), .I1(GND_net), 
            .CO(n36767));
    SB_CARRY add_4467_2 (.CI(GND_net), .I0(n65_adj_3910), .I1(n158_adj_3911), 
            .CO(n36603));
    SB_LUT4 add_4452_9_lut (.I0(GND_net), .I1(n8859[6]), .I2(GND_net), 
            .I3(n36339), .O(n8831[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_10 (.CI(n35963), .I0(n8555[7]), .I1(GND_net), .CO(n35964));
    SB_LUT4 add_4436_9_lut (.I0(GND_net), .I1(n8555[6]), .I2(GND_net), 
            .I3(n35962), .O(n8535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_9 (.CI(n36339), .I0(n8859[6]), .I1(GND_net), .CO(n36340));
    SB_LUT4 add_3176_10_lut (.I0(GND_net), .I1(n1804[22]), .I2(n1711), 
            .I3(n36960), .O(n6821[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_9 (.CI(n35962), .I0(n8555[6]), .I1(GND_net), .CO(n35963));
    SB_LUT4 add_4436_8_lut (.I0(GND_net), .I1(n8555[5]), .I2(n719_adj_3912), 
            .I3(n35961), .O(n8535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_13_lut (.I0(GND_net), .I1(n9146[10]), .I2(GND_net), 
            .I3(n36602), .O(n9132[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_8_lut (.I0(GND_net), .I1(n8859[5]), .I2(n695_adj_3913), 
            .I3(n36338), .O(n8831[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_8 (.CI(n35961), .I0(n8555[5]), .I1(n719_adj_3912), 
            .CO(n35962));
    SB_LUT4 add_4436_7_lut (.I0(GND_net), .I1(n8555[4]), .I2(n622_adj_3914), 
            .I3(n35960), .O(n8535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_7 (.CI(n35960), .I0(n8555[4]), .I1(n622_adj_3914), 
            .CO(n35961));
    SB_CARRY add_4452_8 (.CI(n36338), .I0(n8859[5]), .I1(n695_adj_3913), 
            .CO(n36339));
    SB_LUT4 add_4452_7_lut (.I0(GND_net), .I1(n8859[4]), .I2(n598_adj_3915), 
            .I3(n36337), .O(n8831[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_6_lut (.I0(GND_net), .I1(n8555[3]), .I2(n525_adj_3916), 
            .I3(n35959), .O(n8535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_15 (.CI(n36877), .I0(n1803[12]), .I1(GND_net), 
            .CO(n36878));
    SB_CARRY add_4436_6 (.CI(n35959), .I0(n8555[3]), .I1(n525_adj_3916), 
            .CO(n35960));
    SB_CARRY add_4452_7 (.CI(n36337), .I0(n8859[4]), .I1(n598_adj_3915), 
            .CO(n36338));
    SB_LUT4 add_3176_9_lut (.I0(GND_net), .I1(n1803[22]), .I2(n1707), 
            .I3(n36959), .O(n6821[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_14_lut (.I0(GND_net), .I1(n1803[11]), .I2(GND_net), 
            .I3(n36876), .O(n1802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i142_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n210));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_18_lut (.I0(GND_net), .I1(n1798[15]), .I2(GND_net), 
            .I3(n36765), .O(n1797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_12_lut (.I0(GND_net), .I1(n9146[9]), .I2(GND_net), 
            .I3(n36601), .O(n9132[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_6_lut (.I0(GND_net), .I1(n8859[3]), .I2(n501_adj_3917), 
            .I3(n36336), .O(n8831[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_6 (.CI(n36336), .I0(n8859[3]), .I1(n501_adj_3917), 
            .CO(n36337));
    SB_CARRY add_4466_12 (.CI(n36601), .I0(n9146[9]), .I1(GND_net), .CO(n36602));
    SB_LUT4 add_4452_5_lut (.I0(GND_net), .I1(n8859[2]), .I2(n404_adj_3918), 
            .I3(n36335), .O(n8831[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_5 (.CI(n36335), .I0(n8859[2]), .I1(n404_adj_3918), 
            .CO(n36336));
    SB_CARRY mult_14_add_1212_18 (.CI(n36765), .I0(n1798[15]), .I1(GND_net), 
            .CO(n36766));
    SB_LUT4 add_4466_11_lut (.I0(GND_net), .I1(n9146[8]), .I2(GND_net), 
            .I3(n36600), .O(n9132[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_4_lut (.I0(GND_net), .I1(n8859[1]), .I2(n307_adj_3919), 
            .I3(n36334), .O(n8831[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4452_4 (.CI(n36334), .I0(n8859[1]), .I1(n307_adj_3919), 
            .CO(n36335));
    SB_LUT4 add_4436_5_lut (.I0(GND_net), .I1(n8555[2]), .I2(n428_adj_3920), 
            .I3(n35958), .O(n8535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_5 (.CI(n35958), .I0(n8555[2]), .I1(n428_adj_3920), 
            .CO(n35959));
    SB_LUT4 add_4452_3_lut (.I0(GND_net), .I1(n8859[0]), .I2(n210_adj_3921), 
            .I3(n36333), .O(n8831[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_4_lut (.I0(GND_net), .I1(n8555[1]), .I2(n331_adj_3922), 
            .I3(n35957), .O(n8535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_9 (.CI(n36959), .I0(n1803[22]), .I1(n1707), .CO(n36960));
    SB_CARRY add_4452_3 (.CI(n36333), .I0(n8859[0]), .I1(n210_adj_3921), 
            .CO(n36334));
    SB_CARRY add_4436_4 (.CI(n35957), .I0(n8555[1]), .I1(n331_adj_3922), 
            .CO(n35958));
    SB_LUT4 add_4436_3_lut (.I0(GND_net), .I1(n8555[0]), .I2(n234_adj_3923), 
            .I3(n35956), .O(n8535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_3 (.CI(n35956), .I0(n8555[0]), .I1(n234_adj_3923), 
            .CO(n35957));
    SB_LUT4 mult_14_add_1212_17_lut (.I0(GND_net), .I1(n1798[14]), .I2(GND_net), 
            .I3(n36764), .O(n1797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_11 (.CI(n36600), .I0(n9146[8]), .I1(GND_net), .CO(n36601));
    SB_LUT4 add_3176_8_lut (.I0(GND_net), .I1(n1802[22]), .I2(n1703), 
            .I3(n36958), .O(n6821[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4452_2_lut (.I0(GND_net), .I1(n20_adj_3924), .I2(n113_adj_3925), 
            .I3(GND_net), .O(n8831[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4452_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4436_2_lut (.I0(GND_net), .I1(n44_adj_3926), .I2(n137_adj_3927), 
            .I3(GND_net), .O(n8535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4436_2 (.CI(GND_net), .I0(n44_adj_3926), .I1(n137_adj_3927), 
            .CO(n35956));
    SB_CARRY mult_14_add_1212_17 (.CI(n36764), .I0(n1798[14]), .I1(GND_net), 
            .CO(n36765));
    SB_CARRY add_4452_2 (.CI(GND_net), .I0(n20_adj_3924), .I1(n113_adj_3925), 
            .CO(n36333));
    SB_LUT4 add_4435_20_lut (.I0(GND_net), .I1(n8535[17]), .I2(GND_net), 
            .I3(n35955), .O(n8514[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_19_lut (.I0(GND_net), .I1(n8535[16]), .I2(GND_net), 
            .I3(n35954), .O(n8514[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_14 (.CI(n36876), .I0(n1803[11]), .I1(GND_net), 
            .CO(n36877));
    SB_LUT4 mult_14_add_1212_16_lut (.I0(GND_net), .I1(n1798[13]), .I2(GND_net), 
            .I3(n36763), .O(n1797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_10_lut (.I0(GND_net), .I1(n9146[7]), .I2(GND_net), 
            .I3(n36599), .O(n9132[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_28_lut (.I0(GND_net), .I1(n8831[25]), .I2(GND_net), 
            .I3(n36332), .O(n8802[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_27_lut (.I0(GND_net), .I1(n8831[24]), .I2(GND_net), 
            .I3(n36331), .O(n8802[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_10 (.CI(n36599), .I0(n9146[7]), .I1(GND_net), .CO(n36600));
    SB_CARRY add_4451_27 (.CI(n36331), .I0(n8831[24]), .I1(GND_net), .CO(n36332));
    SB_LUT4 add_4451_26_lut (.I0(GND_net), .I1(n8831[23]), .I2(GND_net), 
            .I3(n36330), .O(n8802[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_16 (.CI(n36763), .I0(n1798[13]), .I1(GND_net), 
            .CO(n36764));
    SB_LUT4 add_4466_9_lut (.I0(GND_net), .I1(n9146[6]), .I2(GND_net), 
            .I3(n36598), .O(n9132[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_26 (.CI(n36330), .I0(n8831[23]), .I1(GND_net), .CO(n36331));
    SB_CARRY add_4435_19 (.CI(n35954), .I0(n8535[16]), .I1(GND_net), .CO(n35955));
    SB_LUT4 add_4435_18_lut (.I0(GND_net), .I1(n8535[15]), .I2(GND_net), 
            .I3(n35953), .O(n8514[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_25_lut (.I0(GND_net), .I1(n8831[22]), .I2(GND_net), 
            .I3(n36329), .O(n8802[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_18 (.CI(n35953), .I0(n8535[15]), .I1(GND_net), .CO(n35954));
    SB_LUT4 add_4435_17_lut (.I0(GND_net), .I1(n8535[14]), .I2(GND_net), 
            .I3(n35952), .O(n8514[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_9 (.CI(n36598), .I0(n9146[6]), .I1(GND_net), .CO(n36599));
    SB_CARRY add_4451_25 (.CI(n36329), .I0(n8831[22]), .I1(GND_net), .CO(n36330));
    SB_CARRY add_4435_17 (.CI(n35952), .I0(n8535[14]), .I1(GND_net), .CO(n35953));
    SB_LUT4 add_4435_16_lut (.I0(GND_net), .I1(n8535[13]), .I2(GND_net), 
            .I3(n35951), .O(n8514[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_24_lut (.I0(GND_net), .I1(n8831[21]), .I2(GND_net), 
            .I3(n36328), .O(n8802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_16 (.CI(n35951), .I0(n8535[13]), .I1(GND_net), .CO(n35952));
    SB_CARRY add_3176_8 (.CI(n36958), .I0(n1802[22]), .I1(n1703), .CO(n36959));
    SB_LUT4 mult_14_add_1217_13_lut (.I0(GND_net), .I1(n1803[10]), .I2(GND_net), 
            .I3(n36875), .O(n1802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_15_lut (.I0(GND_net), .I1(n1798[12]), .I2(GND_net), 
            .I3(n36762), .O(n1797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_8_lut (.I0(GND_net), .I1(n9146[5]), .I2(n737_adj_3928), 
            .I3(n36597), .O(n9132[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_7_lut (.I0(GND_net), .I1(n1801[22]), .I2(n1699), 
            .I3(n36957), .O(n6821[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_8 (.CI(n36597), .I0(n9146[5]), .I1(n737_adj_3928), 
            .CO(n36598));
    SB_CARRY add_4451_24 (.CI(n36328), .I0(n8831[21]), .I1(GND_net), .CO(n36329));
    SB_LUT4 add_4451_23_lut (.I0(GND_net), .I1(n8831[20]), .I2(GND_net), 
            .I3(n36327), .O(n8802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_7_lut (.I0(GND_net), .I1(n9146[4]), .I2(n640_adj_3929), 
            .I3(n36596), .O(n9132[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_15 (.CI(n36762), .I0(n1798[12]), .I1(GND_net), 
            .CO(n36763));
    SB_CARRY add_4466_7 (.CI(n36596), .I0(n9146[4]), .I1(n640_adj_3929), 
            .CO(n36597));
    SB_LUT4 add_4466_6_lut (.I0(GND_net), .I1(n9146[3]), .I2(n543_adj_3930), 
            .I3(n36595), .O(n9132[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_23 (.CI(n36327), .I0(n8831[20]), .I1(GND_net), .CO(n36328));
    SB_LUT4 add_4435_15_lut (.I0(GND_net), .I1(n8535[12]), .I2(GND_net), 
            .I3(n35950), .O(n8514[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_22_lut (.I0(GND_net), .I1(n8831[19]), .I2(GND_net), 
            .I3(n36326), .O(n8802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_6 (.CI(n36595), .I0(n9146[3]), .I1(n543_adj_3930), 
            .CO(n36596));
    SB_CARRY add_4451_22 (.CI(n36326), .I0(n8831[19]), .I1(GND_net), .CO(n36327));
    SB_LUT4 add_4451_21_lut (.I0(GND_net), .I1(n8831[18]), .I2(GND_net), 
            .I3(n36325), .O(n8802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_7 (.CI(n36957), .I0(n1801[22]), .I1(n1699), .CO(n36958));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[19]), .I3(n34691), .O(n39_adj_3931)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n34691), .I0(GND_net), .I1(n76[19]), 
            .CO(n34692));
    SB_LUT4 add_4466_5_lut (.I0(GND_net), .I1(n9146[2]), .I2(n446_adj_3933), 
            .I3(n36594), .O(n9132[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_13 (.CI(n36875), .I0(n1803[10]), .I1(GND_net), 
            .CO(n36876));
    SB_CARRY add_4451_21 (.CI(n36325), .I0(n8831[18]), .I1(GND_net), .CO(n36326));
    SB_LUT4 mult_14_add_1212_14_lut (.I0(GND_net), .I1(n1798[11]), .I2(GND_net), 
            .I3(n36761), .O(n1797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_15 (.CI(n35950), .I0(n8535[12]), .I1(GND_net), .CO(n35951));
    SB_CARRY add_4466_5 (.CI(n36594), .I0(n9146[2]), .I1(n446_adj_3933), 
            .CO(n36595));
    SB_LUT4 add_4435_14_lut (.I0(GND_net), .I1(n8535[11]), .I2(GND_net), 
            .I3(n35949), .O(n8514[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_4_lut (.I0(GND_net), .I1(n9146[1]), .I2(n349_adj_3934), 
            .I3(n36593), .O(n9132[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_20_lut (.I0(GND_net), .I1(n8831[17]), .I2(GND_net), 
            .I3(n36324), .O(n8802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_14 (.CI(n36761), .I0(n1798[11]), .I1(GND_net), 
            .CO(n36762));
    SB_CARRY add_4466_4 (.CI(n36593), .I0(n9146[1]), .I1(n349_adj_3934), 
            .CO(n36594));
    SB_CARRY add_4451_20 (.CI(n36324), .I0(n8831[17]), .I1(GND_net), .CO(n36325));
    SB_LUT4 add_4451_19_lut (.I0(GND_net), .I1(n8831[16]), .I2(GND_net), 
            .I3(n36323), .O(n8802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_19 (.CI(n36323), .I0(n8831[16]), .I1(GND_net), .CO(n36324));
    SB_LUT4 add_4466_3_lut (.I0(GND_net), .I1(n9146[0]), .I2(n252_adj_3935), 
            .I3(n36592), .O(n9132[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_18_lut (.I0(GND_net), .I1(n8831[15]), .I2(GND_net), 
            .I3(n36322), .O(n8802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_14 (.CI(n35949), .I0(n8535[11]), .I1(GND_net), .CO(n35950));
    SB_LUT4 add_4435_13_lut (.I0(GND_net), .I1(n8535[10]), .I2(GND_net), 
            .I3(n35948), .O(n8514[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_18 (.CI(n36322), .I0(n8831[15]), .I1(GND_net), .CO(n36323));
    SB_CARRY add_4435_13 (.CI(n35948), .I0(n8535[10]), .I1(GND_net), .CO(n35949));
    SB_LUT4 state_23__I_0_add_2_26_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n79[23]), .I3(n34844), .O(\PID_CONTROLLER.err_31__N_3175 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[18]), .I3(n34690), .O(n37_adj_3937)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n34690), .I0(GND_net), .I1(n76[18]), 
            .CO(n34691));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n79[23]), .I3(n34843), .O(\PID_CONTROLLER.err_31__N_3175 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_17_lut (.I0(GND_net), .I1(n8831[14]), .I2(GND_net), 
            .I3(n36321), .O(n8802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[17]), .I3(n34689), .O(n35_adj_3939)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_25 (.CI(n34843), .I0(\motor_state[23] ), 
            .I1(n79[23]), .CO(n34844));
    SB_CARRY unary_minus_5_add_3_19 (.CI(n34689), .I0(GND_net), .I1(n76[17]), 
            .CO(n34690));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[16]), .I3(n34688), .O(n33_adj_3941)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(\motor_state[22] ), 
            .I2(n79[22]), .I3(n34842), .O(\PID_CONTROLLER.err_31__N_3175 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_12_lut (.I0(GND_net), .I1(n8535[9]), .I2(GND_net), 
            .I3(n35947), .O(n8514[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_6_lut (.I0(GND_net), .I1(n1800[22]), .I2(n1695), 
            .I3(n36956), .O(n6821[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_12_lut (.I0(GND_net), .I1(n1803[9]), .I2(GND_net), 
            .I3(n36874), .O(n1802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_12 (.CI(n35947), .I0(n8535[9]), .I1(GND_net), .CO(n35948));
    SB_LUT4 mult_14_add_1212_13_lut (.I0(GND_net), .I1(n1798[10]), .I2(GND_net), 
            .I3(n36760), .O(n1797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_3 (.CI(n36592), .I0(n9146[0]), .I1(n252_adj_3935), 
            .CO(n36593));
    SB_LUT4 add_4466_2_lut (.I0(GND_net), .I1(n62_adj_3944), .I2(n155_adj_3945), 
            .I3(GND_net), .O(n9132[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_13 (.CI(n36760), .I0(n1798[10]), .I1(GND_net), 
            .CO(n36761));
    SB_CARRY add_4466_2 (.CI(GND_net), .I0(n62_adj_3944), .I1(n155_adj_3945), 
            .CO(n36592));
    SB_CARRY add_4451_17 (.CI(n36321), .I0(n8831[14]), .I1(GND_net), .CO(n36322));
    SB_LUT4 add_4435_11_lut (.I0(GND_net), .I1(n8535[8]), .I2(GND_net), 
            .I3(n35946), .O(n8514[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n34842), .I0(\motor_state[22] ), 
            .I1(n79[22]), .CO(n34843));
    SB_LUT4 add_4451_16_lut (.I0(GND_net), .I1(n8831[13]), .I2(GND_net), 
            .I3(n36320), .O(n8802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(\motor_state[21] ), 
            .I2(n79[21]), .I3(n34841), .O(\PID_CONTROLLER.err_31__N_3175 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n34841), .I0(\motor_state[21] ), 
            .I1(n79[21]), .CO(n34842));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(\motor_state[20] ), 
            .I2(n79[20]), .I3(n34840), .O(\PID_CONTROLLER.err_31__N_3175 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n34840), .I0(\motor_state[20] ), 
            .I1(n79[20]), .CO(n34841));
    SB_LUT4 add_4465_14_lut (.I0(GND_net), .I1(n9132[11]), .I2(GND_net), 
            .I3(n36591), .O(n9117[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_16 (.CI(n36320), .I0(n8831[13]), .I1(GND_net), .CO(n36321));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n34688), .I0(GND_net), .I1(n76[16]), 
            .CO(n34689));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[15]), .I3(n34687), .O(n31_adj_3948)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4451_15_lut (.I0(GND_net), .I1(n8831[12]), .I2(GND_net), 
            .I3(n36319), .O(n8802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i331_2_lut (.I0(\Kd[5] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n492));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i97_2_lut (.I0(\Kd[1] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n143));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(\motor_state[19] ), 
            .I2(n79[19]), .I3(n34839), .O(\PID_CONTROLLER.err_31__N_3175 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n34687), .I0(GND_net), .I1(n76[15]), 
            .CO(n34688));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[14]), .I3(n34686), .O(n29_adj_3951)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n34839), .I0(\motor_state[19] ), 
            .I1(n79[19]), .CO(n34840));
    SB_LUT4 mult_12_i34_2_lut (.I0(\Kd[0] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i162_2_lut (.I0(\Kd[2] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n240));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i396_2_lut (.I0(\Kd[6] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n589_adj_3465));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4465_13_lut (.I0(GND_net), .I1(n9132[10]), .I2(GND_net), 
            .I3(n36590), .O(n9117[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_15 (.CI(n36319), .I0(n8831[12]), .I1(GND_net), .CO(n36320));
    SB_CARRY add_4435_11 (.CI(n35946), .I0(n8535[8]), .I1(GND_net), .CO(n35947));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(\motor_state[18] ), 
            .I2(n79[18]), .I3(n34838), .O(\PID_CONTROLLER.err_31__N_3175 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n34686), .I0(GND_net), .I1(n76[14]), 
            .CO(n34687));
    SB_CARRY state_23__I_0_add_2_20 (.CI(n34838), .I0(\motor_state[18] ), 
            .I1(n79[18]), .CO(n34839));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(\motor_state[17] ), 
            .I2(n79[17]), .I3(n34837), .O(\PID_CONTROLLER.err_31__N_3175 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_10_lut (.I0(GND_net), .I1(n8535[7]), .I2(GND_net), 
            .I3(n35945), .O(n8514[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1190__i1 (.Q(Kd_delay_counter[1]), .C(clk32MHz), 
           .D(n69[1]));   // verilog/motorControl.v(55[27:47])
    SB_CARRY mult_14_add_1217_12 (.CI(n36874), .I0(n1803[9]), .I1(GND_net), 
            .CO(n36875));
    SB_CARRY state_23__I_0_add_2_19 (.CI(n34837), .I0(\motor_state[17] ), 
            .I1(n79[17]), .CO(n34838));
    SB_LUT4 mult_14_add_1212_12_lut (.I0(GND_net), .I1(n1798[9]), .I2(GND_net), 
            .I3(n36759), .O(n1797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_13 (.CI(n36590), .I0(n9132[10]), .I1(GND_net), .CO(n36591));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[13]), .I3(n34685), .O(n27_adj_3955)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4465_12_lut (.I0(GND_net), .I1(n9132[9]), .I2(GND_net), 
            .I3(n36589), .O(n9117[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n34685), .I0(GND_net), .I1(n76[13]), 
            .CO(n34686));
    SB_CARRY mult_14_add_1212_12 (.CI(n36759), .I0(n1798[9]), .I1(GND_net), 
            .CO(n36760));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(\motor_state[16] ), 
            .I2(n79[16]), .I3(n34836), .O(\PID_CONTROLLER.err_31__N_3175 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_12 (.CI(n36589), .I0(n9132[9]), .I1(GND_net), .CO(n36590));
    SB_LUT4 add_4451_14_lut (.I0(GND_net), .I1(n8831[11]), .I2(GND_net), 
            .I3(n36318), .O(n8802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_11_lut (.I0(GND_net), .I1(n1803[8]), .I2(GND_net), 
            .I3(n36873), .O(n1802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_10 (.CI(n35945), .I0(n8535[7]), .I1(GND_net), .CO(n35946));
    SB_CARRY add_4451_14 (.CI(n36318), .I0(n8831[11]), .I1(GND_net), .CO(n36319));
    SB_LUT4 mult_14_add_1212_11_lut (.I0(GND_net), .I1(n1798[8]), .I2(GND_net), 
            .I3(n36758), .O(n1797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4465_11_lut (.I0(GND_net), .I1(n9132[8]), .I2(GND_net), 
            .I3(n36588), .O(n9117[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_9_lut (.I0(GND_net), .I1(n8535[6]), .I2(GND_net), 
            .I3(n35944), .O(n8514[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n34836), .I0(\motor_state[16] ), 
            .I1(n79[16]), .CO(n34837));
    SB_CARRY mult_14_add_1217_11 (.CI(n36873), .I0(n1803[8]), .I1(GND_net), 
            .CO(n36874));
    SB_CARRY mult_14_add_1212_11 (.CI(n36758), .I0(n1798[8]), .I1(GND_net), 
            .CO(n36759));
    SB_CARRY add_4465_11 (.CI(n36588), .I0(n9132[8]), .I1(GND_net), .CO(n36589));
    SB_LUT4 add_4451_13_lut (.I0(GND_net), .I1(n8831[10]), .I2(GND_net), 
            .I3(n36317), .O(n8802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_9 (.CI(n35944), .I0(n8535[6]), .I1(GND_net), .CO(n35945));
    SB_CARRY add_4451_13 (.CI(n36317), .I0(n8831[10]), .I1(GND_net), .CO(n36318));
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(\motor_state[15] ), 
            .I2(n79[15]), .I3(n34835), .O(\PID_CONTROLLER.err_31__N_3175 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_8_lut (.I0(GND_net), .I1(n8535[5]), .I2(n716_adj_3959), 
            .I3(n35943), .O(n8514[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n34835), .I0(\motor_state[15] ), 
            .I1(n79[15]), .CO(n34836));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[12]), .I3(n34684), .O(n25_adj_3960)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(\motor_state[14] ), 
            .I2(n79[14]), .I3(n34834), .O(\PID_CONTROLLER.err_31__N_3175 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n34684), .I0(GND_net), .I1(n76[12]), 
            .CO(n34685));
    SB_LUT4 add_4465_10_lut (.I0(GND_net), .I1(n9132[7]), .I2(GND_net), 
            .I3(n36587), .O(n9117[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_8 (.CI(n35943), .I0(n8535[5]), .I1(n716_adj_3959), 
            .CO(n35944));
    SB_LUT4 add_4451_12_lut (.I0(GND_net), .I1(n8831[9]), .I2(GND_net), 
            .I3(n36316), .O(n8802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n34834), .I0(\motor_state[14] ), 
            .I1(n79[14]), .CO(n34835));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(\motor_state[13] ), 
            .I2(n79[13]), .I3(n34833), .O(\PID_CONTROLLER.err_31__N_3175 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_12 (.CI(n36316), .I0(n8831[9]), .I1(GND_net), .CO(n36317));
    SB_LUT4 add_4451_11_lut (.I0(GND_net), .I1(n8831[8]), .I2(GND_net), 
            .I3(n36315), .O(n8802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n34833), .I0(\motor_state[13] ), 
            .I1(n79[13]), .CO(n34834));
    SB_CARRY add_4451_11 (.CI(n36315), .I0(n8831[8]), .I1(GND_net), .CO(n36316));
    SB_LUT4 add_4435_7_lut (.I0(GND_net), .I1(n8535[4]), .I2(n619_adj_3964), 
            .I3(n35942), .O(n8514[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[11]), .I3(n34683), .O(n23_adj_3965)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4435_7 (.CI(n35942), .I0(n8535[4]), .I1(n619_adj_3964), 
            .CO(n35943));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n34683), .I0(GND_net), .I1(n76[11]), 
            .CO(n34684));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(\motor_state[12] ), 
            .I2(n79[12]), .I3(n34832), .O(\PID_CONTROLLER.err_31__N_3175 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4435_6_lut (.I0(GND_net), .I1(n8535[3]), .I2(n522_adj_3968), 
            .I3(n35941), .O(n8514[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[10]), .I3(n34682), .O(n21_adj_3969)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n34832), .I0(\motor_state[12] ), 
            .I1(n79[12]), .CO(n34833));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(\motor_state[11] ), 
            .I2(n79[11]), .I3(n34831), .O(\PID_CONTROLLER.err_31__N_3175 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_6 (.CI(n35941), .I0(n8535[3]), .I1(n522_adj_3968), 
            .CO(n35942));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n34682), .I0(GND_net), .I1(n76[10]), 
            .CO(n34683));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n76[9]), .I3(n34681), .O(n19_adj_3972)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n34831), .I0(\motor_state[11] ), 
            .I1(n79[11]), .CO(n34832));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(\motor_state[10] ), 
            .I2(n79[10]), .I3(n34830), .O(\PID_CONTROLLER.err_31__N_3175 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_10 (.CI(n36587), .I0(n9132[7]), .I1(GND_net), .CO(n36588));
    SB_LUT4 mult_14_add_1217_10_lut (.I0(GND_net), .I1(n1803[7]), .I2(GND_net), 
            .I3(n36872), .O(n1802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_10_lut (.I0(GND_net), .I1(n8831[7]), .I2(GND_net), 
            .I3(n36314), .O(n8802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_10 (.CI(n36872), .I0(n1803[7]), .I1(GND_net), 
            .CO(n36873));
    SB_LUT4 add_4435_5_lut (.I0(GND_net), .I1(n8535[2]), .I2(n425_adj_3975), 
            .I3(n35940), .O(n8514[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_5 (.CI(n35940), .I0(n8535[2]), .I1(n425_adj_3975), 
            .CO(n35941));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n34830), .I0(\motor_state[10] ), 
            .I1(n79[10]), .CO(n34831));
    SB_CARRY add_4451_10 (.CI(n36314), .I0(n8831[7]), .I1(GND_net), .CO(n36315));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n34681), .I0(GND_net), .I1(n76[9]), 
            .CO(n34682));
    SB_LUT4 mult_14_add_1212_10_lut (.I0(GND_net), .I1(n1798[7]), .I2(GND_net), 
            .I3(n36757), .O(n1797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_9_lut (.I0(GND_net), .I1(n1803[6]), .I2(GND_net), 
            .I3(n36871), .O(n1802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4465_9_lut (.I0(GND_net), .I1(n9132[6]), .I2(GND_net), 
            .I3(n36586), .O(n9117[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(\motor_state[9] ), 
            .I2(n79[9]), .I3(n34829), .O(\PID_CONTROLLER.err_31__N_3175 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_9_lut (.I0(GND_net), .I1(n8831[6]), .I2(GND_net), 
            .I3(n36313), .O(n8802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n76[8]), .I3(n34680), .O(n17_adj_3977)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1212_10 (.CI(n36757), .I0(n1798[7]), .I1(GND_net), 
            .CO(n36758));
    SB_LUT4 add_4435_4_lut (.I0(GND_net), .I1(n8535[1]), .I2(n328_adj_3979), 
            .I3(n35939), .O(n8514[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n34680), .I0(GND_net), .I1(n76[8]), 
            .CO(n34681));
    SB_CARRY add_4465_9 (.CI(n36586), .I0(n9132[6]), .I1(GND_net), .CO(n36587));
    SB_CARRY mult_14_add_1217_9 (.CI(n36871), .I0(n1803[6]), .I1(GND_net), 
            .CO(n36872));
    SB_LUT4 mult_14_add_1212_9_lut (.I0(GND_net), .I1(n1798[6]), .I2(GND_net), 
            .I3(n36756), .O(n1797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4465_8_lut (.I0(GND_net), .I1(n9132[5]), .I2(n734_adj_3980), 
            .I3(n36585), .O(n9117[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_4 (.CI(n35939), .I0(n8535[1]), .I1(n328_adj_3979), 
            .CO(n35940));
    SB_CARRY add_4465_8 (.CI(n36585), .I0(n9132[5]), .I1(n734_adj_3980), 
            .CO(n36586));
    SB_LUT4 add_4465_7_lut (.I0(GND_net), .I1(n9132[4]), .I2(n637_adj_3981), 
            .I3(n36584), .O(n9117[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_9 (.CI(n36313), .I0(n8831[6]), .I1(GND_net), .CO(n36314));
    SB_LUT4 add_4435_3_lut (.I0(GND_net), .I1(n8535[0]), .I2(n231_adj_3982), 
            .I3(n35938), .O(n8514[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4435_3 (.CI(n35938), .I0(n8535[0]), .I1(n231_adj_3982), 
            .CO(n35939));
    SB_LUT4 add_4435_2_lut (.I0(GND_net), .I1(n41_adj_3983), .I2(n134_adj_3984), 
            .I3(GND_net), .O(n8514[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4435_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n34829), .I0(\motor_state[9] ), 
            .I1(n79[9]), .CO(n34830));
    SB_CARRY mult_14_add_1212_9 (.CI(n36756), .I0(n1798[6]), .I1(GND_net), 
            .CO(n36757));
    SB_LUT4 add_4451_8_lut (.I0(GND_net), .I1(n8831[5]), .I2(n692_adj_3985), 
            .I3(n36312), .O(n8802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_7 (.CI(n36584), .I0(n9132[4]), .I1(n637_adj_3981), 
            .CO(n36585));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(\motor_state[8] ), 
            .I2(n79[8]), .I3(n34828), .O(\PID_CONTROLLER.err_31__N_3175 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n76[7]), .I3(n34679), .O(n15_adj_3987)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4451_8 (.CI(n36312), .I0(n8831[5]), .I1(n692_adj_3985), 
            .CO(n36313));
    SB_CARRY add_4435_2 (.CI(GND_net), .I0(n41_adj_3983), .I1(n134_adj_3984), 
            .CO(n35938));
    SB_LUT4 add_4451_7_lut (.I0(GND_net), .I1(n8831[4]), .I2(n595_adj_3989), 
            .I3(n36311), .O(n8802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_21_lut (.I0(GND_net), .I1(n8514[18]), .I2(GND_net), 
            .I3(n35937), .O(n8492[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_6 (.CI(n36956), .I0(n1800[22]), .I1(n1695), .CO(n36957));
    SB_LUT4 add_3176_5_lut (.I0(GND_net), .I1(n1799[22]), .I2(n1691), 
            .I3(n36955), .O(n6821[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n34828), .I0(\motor_state[8] ), 
            .I1(n79[8]), .CO(n34829));
    SB_LUT4 add_4465_6_lut (.I0(GND_net), .I1(n9132[3]), .I2(n540_adj_3990), 
            .I3(n36583), .O(n9117[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_7 (.CI(n36311), .I0(n8831[4]), .I1(n595_adj_3989), 
            .CO(n36312));
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(\motor_state[7] ), 
            .I2(n79[7]), .I3(n34827), .O(\PID_CONTROLLER.err_31__N_3175 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n34679), .I0(GND_net), .I1(n76[7]), 
            .CO(n34680));
    SB_LUT4 add_4434_20_lut (.I0(GND_net), .I1(n8514[17]), .I2(GND_net), 
            .I3(n35936), .O(n8492[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_20 (.CI(n35936), .I0(n8514[17]), .I1(GND_net), .CO(n35937));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n76[6]), .I3(n34678), .O(n13_adj_3992)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1217_8_lut (.I0(GND_net), .I1(n1803[5]), .I2(n530), 
            .I3(n36870), .O(n1802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n34678), .I0(GND_net), .I1(n76[6]), 
            .CO(n34679));
    SB_LUT4 add_4451_6_lut (.I0(GND_net), .I1(n8831[3]), .I2(n498_adj_3994), 
            .I3(n36310), .O(n8802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_6 (.CI(n36310), .I0(n8831[3]), .I1(n498_adj_3994), 
            .CO(n36311));
    SB_LUT4 mult_14_add_1212_8_lut (.I0(GND_net), .I1(n1798[5]), .I2(n515), 
            .I3(n36755), .O(n1797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_6 (.CI(n36583), .I0(n9132[3]), .I1(n540_adj_3990), 
            .CO(n36584));
    SB_LUT4 add_4434_19_lut (.I0(GND_net), .I1(n8514[16]), .I2(GND_net), 
            .I3(n35935), .O(n8492[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_19 (.CI(n35935), .I0(n8514[16]), .I1(GND_net), .CO(n35936));
    SB_LUT4 add_4451_5_lut (.I0(GND_net), .I1(n8831[2]), .I2(n401_adj_3995), 
            .I3(n36309), .O(n8802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_18_lut (.I0(GND_net), .I1(n8514[15]), .I2(GND_net), 
            .I3(n35934), .O(n8492[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_18 (.CI(n35934), .I0(n8514[15]), .I1(GND_net), .CO(n35935));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n34827), .I0(\motor_state[7] ), 
            .I1(n79[7]), .CO(n34828));
    SB_CARRY add_4451_5 (.CI(n36309), .I0(n8831[2]), .I1(n401_adj_3995), 
            .CO(n36310));
    SB_LUT4 add_4465_5_lut (.I0(GND_net), .I1(n9132[2]), .I2(n443_adj_3996), 
            .I3(n36582), .O(n9117[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_17_lut (.I0(GND_net), .I1(n8514[14]), .I2(GND_net), 
            .I3(n35933), .O(n8492[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_17 (.CI(n35933), .I0(n8514[14]), .I1(GND_net), .CO(n35934));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(\motor_state[6] ), 
            .I2(n79[6]), .I3(n34826), .O(\PID_CONTROLLER.err_31__N_3175 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_16_lut (.I0(GND_net), .I1(n8514[13]), .I2(GND_net), 
            .I3(n35932), .O(n8492[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n76[5]), .I3(n34677), .O(n11_adj_3998)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4465_5 (.CI(n36582), .I0(n9132[2]), .I1(n443_adj_3996), 
            .CO(n36583));
    SB_LUT4 add_4451_4_lut (.I0(GND_net), .I1(n8831[1]), .I2(n304_adj_4000), 
            .I3(n36308), .O(n8802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_8 (.CI(n36870), .I0(n1803[5]), .I1(n530), 
            .CO(n36871));
    SB_CARRY mult_14_add_1212_8 (.CI(n36755), .I0(n1798[5]), .I1(n515), 
            .CO(n36756));
    SB_CARRY add_4434_16 (.CI(n35932), .I0(n8514[13]), .I1(GND_net), .CO(n35933));
    SB_LUT4 mult_14_add_1212_7_lut (.I0(GND_net), .I1(n1798[4]), .I2(n442), 
            .I3(n36754), .O(n1797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_7 (.CI(n36754), .I0(n1798[4]), .I1(n442), 
            .CO(n36755));
    SB_LUT4 add_4465_4_lut (.I0(GND_net), .I1(n9132[1]), .I2(n346_adj_4001), 
            .I3(n36581), .O(n9117[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_4 (.CI(n36581), .I0(n9132[1]), .I1(n346_adj_4001), 
            .CO(n36582));
    SB_LUT4 add_4434_15_lut (.I0(GND_net), .I1(n8514[12]), .I2(GND_net), 
            .I3(n35931), .O(n8492[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_6_lut (.I0(GND_net), .I1(n1798[3]), .I2(n369), 
            .I3(n36753), .O(n1797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4465_3_lut (.I0(GND_net), .I1(n9132[0]), .I2(n249_adj_4002), 
            .I3(n36580), .O(n9117[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_4 (.CI(n36308), .I0(n8831[1]), .I1(n304_adj_4000), 
            .CO(n36309));
    SB_CARRY add_4434_15 (.CI(n35931), .I0(n8514[12]), .I1(GND_net), .CO(n35932));
    SB_CARRY state_23__I_0_add_2_8 (.CI(n34826), .I0(\motor_state[6] ), 
            .I1(n79[6]), .CO(n34827));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(\motor_state[5] ), 
            .I2(n79[5]), .I3(n34825), .O(\PID_CONTROLLER.err_31__N_3175 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_14_lut (.I0(GND_net), .I1(n8514[11]), .I2(GND_net), 
            .I3(n35930), .O(n8492[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_14 (.CI(n35930), .I0(n8514[11]), .I1(GND_net), .CO(n35931));
    SB_CARRY state_23__I_0_add_2_7 (.CI(n34825), .I0(\motor_state[5] ), 
            .I1(n79[5]), .CO(n34826));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n34677), .I0(GND_net), .I1(n76[5]), 
            .CO(n34678));
    SB_LUT4 add_4434_13_lut (.I0(GND_net), .I1(n8514[10]), .I2(GND_net), 
            .I3(n35929), .O(n8492[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n76[4]), .I3(n34676), .O(n9_adj_4004)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(\motor_state[4] ), 
            .I2(n79[4]), .I3(n34824), .O(\PID_CONTROLLER.err_31__N_3175 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_3 (.CI(n36580), .I0(n9132[0]), .I1(n249_adj_4002), 
            .CO(n36581));
    SB_LUT4 add_4451_3_lut (.I0(GND_net), .I1(n8831[0]), .I2(n207_adj_4007), 
            .I3(n36307), .O(n8802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_13 (.CI(n35929), .I0(n8514[10]), .I1(GND_net), .CO(n35930));
    SB_CARRY add_4451_3 (.CI(n36307), .I0(n8831[0]), .I1(n207_adj_4007), 
            .CO(n36308));
    SB_LUT4 add_4451_2_lut (.I0(GND_net), .I1(n17_adj_4008), .I2(n110_adj_4009), 
            .I3(GND_net), .O(n8802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4465_2_lut (.I0(GND_net), .I1(n59_adj_4010), .I2(n152_adj_4011), 
            .I3(GND_net), .O(n9117[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4465_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_2 (.CI(GND_net), .I0(n17_adj_4008), .I1(n110_adj_4009), 
            .CO(n36307));
    SB_LUT4 add_4434_12_lut (.I0(GND_net), .I1(n8514[9]), .I2(GND_net), 
            .I3(n35928), .O(n8492[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_12 (.CI(n35928), .I0(n8514[9]), .I1(GND_net), .CO(n35929));
    SB_LUT4 add_4450_29_lut (.I0(GND_net), .I1(n8802[26]), .I2(GND_net), 
            .I3(n36306), .O(n8772[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_11_lut (.I0(GND_net), .I1(n8514[8]), .I2(GND_net), 
            .I3(n35927), .O(n8492[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_28_lut (.I0(GND_net), .I1(n8802[25]), .I2(GND_net), 
            .I3(n36305), .O(n8772[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4465_2 (.CI(GND_net), .I0(n59_adj_4010), .I1(n152_adj_4011), 
            .CO(n36580));
    SB_LUT4 add_4464_15_lut (.I0(GND_net), .I1(n9117[12]), .I2(GND_net), 
            .I3(n36579), .O(n9101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n34824), .I0(\motor_state[4] ), 
            .I1(n79[4]), .CO(n34825));
    SB_CARRY add_4434_11 (.CI(n35927), .I0(n8514[8]), .I1(GND_net), .CO(n35928));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(\motor_state[3] ), 
            .I2(n79[3]), .I3(n34823), .O(\PID_CONTROLLER.err_31__N_3175 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_28 (.CI(n36305), .I0(n8802[25]), .I1(GND_net), .CO(n36306));
    SB_CARRY add_3176_5 (.CI(n36955), .I0(n1799[22]), .I1(n1691), .CO(n36956));
    SB_LUT4 add_4450_27_lut (.I0(GND_net), .I1(n8802[24]), .I2(GND_net), 
            .I3(n36304), .O(n8772[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_10_lut (.I0(GND_net), .I1(n8514[7]), .I2(GND_net), 
            .I3(n35926), .O(n8492[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4464_14_lut (.I0(GND_net), .I1(n9117[11]), .I2(GND_net), 
            .I3(n36578), .O(n9101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n34676), .I0(GND_net), .I1(n76[4]), 
            .CO(n34677));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n76[3]), .I3(n34675), .O(n7_adj_4013)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4450_27 (.CI(n36304), .I0(n8802[24]), .I1(GND_net), .CO(n36305));
    SB_CARRY add_4434_10 (.CI(n35926), .I0(n8514[7]), .I1(GND_net), .CO(n35927));
    SB_CARRY state_23__I_0_add_2_5 (.CI(n34823), .I0(\motor_state[3] ), 
            .I1(n79[3]), .CO(n34824));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(\motor_state[2] ), 
            .I2(n79[2]), .I3(n34822), .O(\PID_CONTROLLER.err_31__N_3175 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_9_lut (.I0(GND_net), .I1(n8514[6]), .I2(GND_net), 
            .I3(n35925), .O(n8492[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_9 (.CI(n35925), .I0(n8514[6]), .I1(GND_net), .CO(n35926));
    SB_LUT4 add_4434_8_lut (.I0(GND_net), .I1(n8514[5]), .I2(n713_adj_4016), 
            .I3(n35924), .O(n8492[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_7_lut (.I0(GND_net), .I1(n1803[4]), .I2(n457_adj_4017), 
            .I3(n36869), .O(n1802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_6 (.CI(n36753), .I0(n1798[3]), .I1(n369), 
            .CO(n36754));
    SB_CARRY add_4464_14 (.CI(n36578), .I0(n9117[11]), .I1(GND_net), .CO(n36579));
    SB_LUT4 add_4450_26_lut (.I0(GND_net), .I1(n8802[23]), .I2(GND_net), 
            .I3(n36303), .O(n8772[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_26 (.CI(n36303), .I0(n8802[23]), .I1(GND_net), .CO(n36304));
    SB_LUT4 add_4464_13_lut (.I0(GND_net), .I1(n9117[10]), .I2(GND_net), 
            .I3(n36577), .O(n9101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_25_lut (.I0(GND_net), .I1(n8802[22]), .I2(GND_net), 
            .I3(n36302), .O(n8772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_5_lut (.I0(GND_net), .I1(n1798[2]), .I2(n296_adj_4018), 
            .I3(n36752), .O(n1797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4464_13 (.CI(n36577), .I0(n9117[10]), .I1(GND_net), .CO(n36578));
    SB_CARRY add_4450_25 (.CI(n36302), .I0(n8802[22]), .I1(GND_net), .CO(n36303));
    SB_LUT4 add_4464_12_lut (.I0(GND_net), .I1(n9117[9]), .I2(GND_net), 
            .I3(n36576), .O(n9101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4464_12 (.CI(n36576), .I0(n9117[9]), .I1(GND_net), .CO(n36577));
    SB_LUT4 add_4450_24_lut (.I0(GND_net), .I1(n8802[21]), .I2(GND_net), 
            .I3(n36301), .O(n8772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_4_lut (.I0(GND_net), .I1(n1798[22]), .I2(n1687), 
            .I3(n36954), .O(n6821[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_24 (.CI(n36301), .I0(n8802[21]), .I1(GND_net), .CO(n36302));
    SB_CARRY mult_14_add_1217_7 (.CI(n36869), .I0(n1803[4]), .I1(n457_adj_4017), 
            .CO(n36870));
    SB_CARRY mult_14_add_1212_5 (.CI(n36752), .I0(n1798[2]), .I1(n296_adj_4018), 
            .CO(n36753));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n34822), .I0(\motor_state[2] ), 
            .I1(n79[2]), .CO(n34823));
    SB_LUT4 add_4464_11_lut (.I0(GND_net), .I1(n9117[8]), .I2(GND_net), 
            .I3(n36575), .O(n9101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(\motor_state[1] ), 
            .I2(n79[1]), .I3(n34821), .O(\PID_CONTROLLER.err_31__N_3175 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_23_lut (.I0(GND_net), .I1(n8802[20]), .I2(GND_net), 
            .I3(n36300), .O(n8772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n34675), .I0(GND_net), .I1(n76[3]), 
            .CO(n34676));
    SB_CARRY add_4434_8 (.CI(n35924), .I0(n8514[5]), .I1(n713_adj_4016), 
            .CO(n35925));
    SB_CARRY add_4464_11 (.CI(n36575), .I0(n9117[8]), .I1(GND_net), .CO(n36576));
    SB_LUT4 mult_14_add_1212_4_lut (.I0(GND_net), .I1(n1798[1]), .I2(n223_adj_4020), 
            .I3(n36751), .O(n1797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_4 (.CI(n36954), .I0(n1798[22]), .I1(n1687), .CO(n36955));
    SB_LUT4 add_4464_10_lut (.I0(GND_net), .I1(n9117[7]), .I2(GND_net), 
            .I3(n36574), .O(n9101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n34821), .I0(\motor_state[1] ), 
            .I1(n79[1]), .CO(n34822));
    SB_CARRY add_4464_10 (.CI(n36574), .I0(n9117[7]), .I1(GND_net), .CO(n36575));
    SB_LUT4 mult_14_add_1217_6_lut (.I0(GND_net), .I1(n1803[3]), .I2(n384), 
            .I3(n36868), .O(n1802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_4 (.CI(n36751), .I0(n1798[1]), .I1(n223_adj_4020), 
            .CO(n36752));
    SB_LUT4 add_4464_9_lut (.I0(GND_net), .I1(n9117[6]), .I2(GND_net), 
            .I3(n36573), .O(n9101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n76[2]), .I3(n34674), .O(n5_adj_4021)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4464_9 (.CI(n36573), .I0(n9117[6]), .I1(GND_net), .CO(n36574));
    SB_LUT4 mult_14_add_1212_3_lut (.I0(GND_net), .I1(n1798[0]), .I2(n150_adj_4023), 
            .I3(n36750), .O(n1797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_3_lut (.I0(GND_net), .I1(n1797[22]), .I2(n1683), 
            .I3(n36953), .O(n6821[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_7_lut (.I0(GND_net), .I1(n8514[4]), .I2(n616_adj_4024), 
            .I3(n35923), .O(n8492[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_3 (.CI(n36953), .I0(n1797[22]), .I1(n1683), .CO(n36954));
    SB_CARRY add_4450_23 (.CI(n36300), .I0(n8802[20]), .I1(GND_net), .CO(n36301));
    SB_CARRY add_4434_7 (.CI(n35923), .I0(n8514[4]), .I1(n616_adj_4024), 
            .CO(n35924));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(\motor_state[0] ), 
            .I2(n79[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_31__N_3175 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4464_8_lut (.I0(GND_net), .I1(n9117[5]), .I2(n731_adj_4026), 
            .I3(n36572), .O(n9101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_6_lut (.I0(GND_net), .I1(n8514[3]), .I2(n519_adj_4027), 
            .I3(n35922), .O(n8492[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4464_8 (.CI(n36572), .I0(n9117[5]), .I1(n731_adj_4026), 
            .CO(n36573));
    SB_LUT4 add_4464_7_lut (.I0(GND_net), .I1(n9117[4]), .I2(n634_adj_4028), 
            .I3(n36571), .O(n9101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(\motor_state[0] ), 
            .I1(n79[0]), .CO(n34821));
    SB_LUT4 add_3176_2_lut (.I0(GND_net), .I1(n1796[22]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n6821[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n34674), .I0(GND_net), .I1(n76[2]), 
            .CO(n34675));
    SB_CARRY mult_14_add_1217_6 (.CI(n36868), .I0(n1803[3]), .I1(n384), 
            .CO(n36869));
    SB_LUT4 mult_14_add_1217_5_lut (.I0(GND_net), .I1(n1803[2]), .I2(n311_adj_4029), 
            .I3(n36867), .O(n1802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_3 (.CI(n36750), .I0(n1798[0]), .I1(n150_adj_4023), 
            .CO(n36751));
    SB_CARRY add_4464_7 (.CI(n36571), .I0(n9117[4]), .I1(n634_adj_4028), 
            .CO(n36572));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n76[1]), .I3(n34673), .O(n3_adj_4030)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4450_22_lut (.I0(GND_net), .I1(n8802[19]), .I2(GND_net), 
            .I3(n36299), .O(n8772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_22 (.CI(n36299), .I0(n8802[19]), .I1(GND_net), .CO(n36300));
    SB_LUT4 add_4464_6_lut (.I0(GND_net), .I1(n9117[3]), .I2(n537_adj_4032), 
            .I3(n36570), .O(n9101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_21_lut (.I0(GND_net), .I1(n8802[18]), .I2(GND_net), 
            .I3(n36298), .O(n8772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_2 (.CI(GND_net), .I0(n1796[22]), .I1(\PID_CONTROLLER.integral [9]), 
            .CO(n36953));
    SB_LUT4 add_4473_22_lut (.I0(GND_net), .I1(n9555[19]), .I2(GND_net), 
            .I3(n36952), .O(n9225[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_21 (.CI(n36298), .I0(n8802[18]), .I1(GND_net), .CO(n36299));
    SB_LUT4 add_4450_20_lut (.I0(GND_net), .I1(n8802[17]), .I2(GND_net), 
            .I3(n36297), .O(n8772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_6 (.CI(n35922), .I0(n8514[3]), .I1(n519_adj_4027), 
            .CO(n35923));
    SB_LUT4 mult_14_add_1212_2_lut (.I0(GND_net), .I1(n8_adj_4033), .I2(n77), 
            .I3(GND_net), .O(n1797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4464_6 (.CI(n36570), .I0(n9117[3]), .I1(n537_adj_4032), 
            .CO(n36571));
    SB_CARRY add_4450_20 (.CI(n36297), .I0(n8802[17]), .I1(GND_net), .CO(n36298));
    SB_LUT4 add_4450_19_lut (.I0(GND_net), .I1(n8802[16]), .I2(GND_net), 
            .I3(n36296), .O(n8772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_5_lut (.I0(GND_net), .I1(n8514[2]), .I2(n422_adj_4034), 
            .I3(n35921), .O(n8492[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4464_5_lut (.I0(GND_net), .I1(n9117[2]), .I2(n440_adj_4035), 
            .I3(n36569), .O(n9101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_19 (.CI(n36296), .I0(n8802[16]), .I1(GND_net), .CO(n36297));
    SB_LUT4 add_4450_18_lut (.I0(GND_net), .I1(n8802[15]), .I2(GND_net), 
            .I3(n36295), .O(n8772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_5 (.CI(n35921), .I0(n8514[2]), .I1(n422_adj_4034), 
            .CO(n35922));
    SB_CARRY mult_14_add_1217_5 (.CI(n36867), .I0(n1803[2]), .I1(n311_adj_4029), 
            .CO(n36868));
    SB_CARRY mult_14_add_1212_2 (.CI(GND_net), .I0(n8_adj_4033), .I1(n77), 
            .CO(n36750));
    SB_CARRY add_4464_5 (.CI(n36569), .I0(n9117[2]), .I1(n440_adj_4035), 
            .CO(n36570));
    SB_CARRY add_4450_18 (.CI(n36295), .I0(n8802[15]), .I1(GND_net), .CO(n36296));
    SB_LUT4 add_4450_17_lut (.I0(GND_net), .I1(n8802[14]), .I2(GND_net), 
            .I3(n36294), .O(n8772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_4_lut (.I0(GND_net), .I1(n8514[1]), .I2(n325_adj_4036), 
            .I3(n35920), .O(n8492[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_4 (.CI(n35920), .I0(n8514[1]), .I1(n325_adj_4036), 
            .CO(n35921));
    SB_LUT4 add_4464_4_lut (.I0(GND_net), .I1(n9117[1]), .I2(n343_adj_4037), 
            .I3(n36568), .O(n9101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4464_4 (.CI(n36568), .I0(n9117[1]), .I1(n343_adj_4037), 
            .CO(n36569));
    SB_CARRY add_4450_17 (.CI(n36294), .I0(n8802[14]), .I1(GND_net), .CO(n36295));
    SB_LUT4 add_4473_21_lut (.I0(GND_net), .I1(n9555[18]), .I2(GND_net), 
            .I3(n36951), .O(n9225[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_16_lut (.I0(GND_net), .I1(n8802[13]), .I2(GND_net), 
            .I3(n36293), .O(n8772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_3_lut (.I0(GND_net), .I1(n8514[0]), .I2(n228_adj_4038), 
            .I3(n35919), .O(n8492[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_24_lut (.I0(GND_net), .I1(n1797[21]), .I2(GND_net), 
            .I3(n36748), .O(n1796[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1190__i2 (.Q(Kd_delay_counter[2]), .C(clk32MHz), 
           .D(n69[2]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1190__i3 (.Q(Kd_delay_counter[3]), .C(clk32MHz), 
           .D(n69[3]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1190__i4 (.Q(Kd_delay_counter[4]), .C(clk32MHz), 
           .D(n69[4]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1190__i5 (.Q(Kd_delay_counter[5]), .C(clk32MHz), 
           .D(n69[5]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1190__i6 (.Q(Kd_delay_counter[6]), .C(clk32MHz), 
           .D(n69[6]));   // verilog/motorControl.v(55[27:47])
    SB_DFF pwm_count_1191__i1 (.Q(pwm_count[1]), .C(clk32MHz), .D(n70[1]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i2 (.Q(pwm_count[2]), .C(clk32MHz), .D(n70[2]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i3 (.Q(pwm_count[3]), .C(clk32MHz), .D(n70[3]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i4 (.Q(pwm_count[4]), .C(clk32MHz), .D(n70[4]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i5 (.Q(pwm_count[5]), .C(clk32MHz), .D(n70[5]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i6 (.Q(pwm_count[6]), .C(clk32MHz), .D(n70[6]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i7 (.Q(pwm_count[7]), .C(clk32MHz), .D(n70[7]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1191__i8 (.Q(pwm_count[8]), .C(clk32MHz), .D(n70[8]));   // verilog/motorControl.v(110[18:29])
    SB_DFFE \PID_CONTROLLER.integral_1192__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[1]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[2]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[3]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[4]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[5]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[6]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[7]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[8]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1192__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(n55_adj_3736), .D(n73[9]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 add_4464_3_lut (.I0(GND_net), .I1(n9117[0]), .I2(n246_adj_4039), 
            .I3(n36567), .O(n9101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_16 (.CI(n36293), .I0(n8802[13]), .I1(GND_net), .CO(n36294));
    SB_LUT4 add_4450_15_lut (.I0(GND_net), .I1(n8802[12]), .I2(GND_net), 
            .I3(n36292), .O(n8772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_3 (.CI(n35919), .I0(n8514[0]), .I1(n228_adj_4038), 
            .CO(n35920));
    SB_CARRY add_4464_3 (.CI(n36567), .I0(n9117[0]), .I1(n246_adj_4039), 
            .CO(n36568));
    SB_CARRY add_4450_15 (.CI(n36292), .I0(n8802[12]), .I1(GND_net), .CO(n36293));
    SB_LUT4 add_4450_14_lut (.I0(GND_net), .I1(n8802[11]), .I2(GND_net), 
            .I3(n36291), .O(n8772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4434_2_lut (.I0(GND_net), .I1(n38_adj_4040), .I2(n131_adj_4041), 
            .I3(GND_net), .O(n8492[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4434_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_21 (.CI(n36951), .I0(n9555[18]), .I1(GND_net), .CO(n36952));
    SB_LUT4 mult_14_add_1217_4_lut (.I0(GND_net), .I1(n1803[1]), .I2(n238_adj_4042), 
            .I3(n36866), .O(n1802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_24 (.CI(n36748), .I0(n1797[21]), .I1(GND_net), 
            .CO(n1683));
    SB_LUT4 add_4464_2_lut (.I0(GND_net), .I1(n56_adj_4043), .I2(n149_adj_4044), 
            .I3(GND_net), .O(n9101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4464_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_14 (.CI(n36291), .I0(n8802[11]), .I1(GND_net), .CO(n36292));
    SB_LUT4 add_4450_13_lut (.I0(GND_net), .I1(n8802[10]), .I2(GND_net), 
            .I3(n36290), .O(n8772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4434_2 (.CI(GND_net), .I0(n38_adj_4040), .I1(n131_adj_4041), 
            .CO(n35919));
    SB_CARRY add_4464_2 (.CI(GND_net), .I0(n56_adj_4043), .I1(n149_adj_4044), 
            .CO(n36567));
    SB_CARRY add_4450_13 (.CI(n36290), .I0(n8802[10]), .I1(GND_net), .CO(n36291));
    SB_LUT4 add_4450_12_lut (.I0(GND_net), .I1(n8802[9]), .I2(GND_net), 
            .I3(n36289), .O(n8772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_12 (.CI(n36289), .I0(n8802[9]), .I1(GND_net), .CO(n36290));
    SB_LUT4 mult_14_add_1211_23_lut (.I0(GND_net), .I1(n1797[20]), .I2(GND_net), 
            .I3(n36747), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_16_lut (.I0(GND_net), .I1(n9101[13]), .I2(GND_net), 
            .I3(n36566), .O(n9084[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_15_lut (.I0(GND_net), .I1(n9101[12]), .I2(GND_net), 
            .I3(n36565), .O(n9084[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4450_11_lut (.I0(GND_net), .I1(n8802[8]), .I2(GND_net), 
            .I3(n36288), .O(n8772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_11 (.CI(n36288), .I0(n8802[8]), .I1(GND_net), .CO(n36289));
    SB_LUT4 add_4450_10_lut (.I0(GND_net), .I1(n8802[7]), .I2(GND_net), 
            .I3(n36287), .O(n8772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_20_lut (.I0(GND_net), .I1(n9555[17]), .I2(GND_net), 
            .I3(n36950), .O(n9225[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_15 (.CI(n36565), .I0(n9101[12]), .I1(GND_net), .CO(n36566));
    SB_LUT4 add_4463_14_lut (.I0(GND_net), .I1(n9101[11]), .I2(GND_net), 
            .I3(n36564), .O(n9084[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_10 (.CI(n36287), .I0(n8802[7]), .I1(GND_net), .CO(n36288));
    SB_LUT4 add_4450_9_lut (.I0(GND_net), .I1(n8802[6]), .I2(GND_net), 
            .I3(n36286), .O(n8772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_4 (.CI(n36866), .I0(n1803[1]), .I1(n238_adj_4042), 
            .CO(n36867));
    SB_CARRY mult_14_add_1211_23 (.CI(n36747), .I0(n1797[20]), .I1(GND_net), 
            .CO(n36748));
    SB_CARRY add_4463_14 (.CI(n36564), .I0(n9101[11]), .I1(GND_net), .CO(n36565));
    SB_CARRY add_4450_9 (.CI(n36286), .I0(n8802[6]), .I1(GND_net), .CO(n36287));
    SB_LUT4 add_4450_8_lut (.I0(GND_net), .I1(n8802[5]), .I2(n689_adj_4045), 
            .I3(n36285), .O(n8772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_13_lut (.I0(GND_net), .I1(n9101[10]), .I2(GND_net), 
            .I3(n36563), .O(n9084[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_8 (.CI(n36285), .I0(n8802[5]), .I1(n689_adj_4045), 
            .CO(n36286));
    SB_LUT4 add_4450_7_lut (.I0(GND_net), .I1(n8802[4]), .I2(n592_adj_4046), 
            .I3(n36284), .O(n8772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_22_lut (.I0(GND_net), .I1(n1797[19]), .I2(GND_net), 
            .I3(n36746), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_13 (.CI(n36563), .I0(n9101[10]), .I1(GND_net), .CO(n36564));
    SB_CARRY add_4450_7 (.CI(n36284), .I0(n8802[4]), .I1(n592_adj_4046), 
            .CO(n36285));
    SB_LUT4 add_4450_6_lut (.I0(GND_net), .I1(n8802[3]), .I2(n495_adj_4047), 
            .I3(n36283), .O(n8772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_12_lut (.I0(GND_net), .I1(n9101[9]), .I2(GND_net), 
            .I3(n36562), .O(n9084[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_6 (.CI(n36283), .I0(n8802[3]), .I1(n495_adj_4047), 
            .CO(n36284));
    SB_LUT4 add_4450_5_lut (.I0(GND_net), .I1(n8802[2]), .I2(n398_adj_4048), 
            .I3(n36282), .O(n8772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_20 (.CI(n36950), .I0(n9555[17]), .I1(GND_net), .CO(n36951));
    SB_CARRY add_4450_5 (.CI(n36282), .I0(n8802[2]), .I1(n398_adj_4048), 
            .CO(n36283));
    SB_LUT4 mult_14_add_1217_3_lut (.I0(GND_net), .I1(n1803[0]), .I2(n165_adj_4049), 
            .I3(n36865), .O(n1802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n34673), .I0(GND_net), .I1(n76[1]), 
            .CO(n34674));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n76[0]), 
            .I3(VCC_net), .O(n75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_22 (.CI(n36746), .I0(n1797[19]), .I1(GND_net), 
            .CO(n36747));
    SB_LUT4 mult_14_add_1211_21_lut (.I0(GND_net), .I1(n1797[18]), .I2(GND_net), 
            .I3(n36745), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_12 (.CI(n36562), .I0(n9101[9]), .I1(GND_net), .CO(n36563));
    SB_CARRY mult_14_add_1217_3 (.CI(n36865), .I0(n1803[0]), .I1(n165_adj_4049), 
            .CO(n36866));
    SB_LUT4 add_4433_22_lut (.I0(GND_net), .I1(n8492[19]), .I2(GND_net), 
            .I3(n35918), .O(n8469[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_11_lut (.I0(GND_net), .I1(n9101[8]), .I2(GND_net), 
            .I3(n36561), .O(n9084[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_21_lut (.I0(GND_net), .I1(n8492[18]), .I2(GND_net), 
            .I3(n35917), .O(n8469[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_21 (.CI(n36745), .I0(n1797[18]), .I1(GND_net), 
            .CO(n36746));
    SB_CARRY add_4463_11 (.CI(n36561), .I0(n9101[8]), .I1(GND_net), .CO(n36562));
    SB_CARRY add_4433_21 (.CI(n35917), .I0(n8492[18]), .I1(GND_net), .CO(n35918));
    SB_LUT4 add_4463_10_lut (.I0(GND_net), .I1(n9101[7]), .I2(GND_net), 
            .I3(n36560), .O(n9084[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_20_lut (.I0(GND_net), .I1(n8492[17]), .I2(GND_net), 
            .I3(n35916), .O(n8469[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_2_lut (.I0(GND_net), .I1(n23_adj_4052), .I2(n92), 
            .I3(GND_net), .O(n1802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_20_lut (.I0(GND_net), .I1(n1797[17]), .I2(GND_net), 
            .I3(n36744), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_10 (.CI(n36560), .I0(n9101[7]), .I1(GND_net), .CO(n36561));
    SB_LUT4 add_4450_4_lut (.I0(GND_net), .I1(n8802[1]), .I2(n301_adj_4053), 
            .I3(n36281), .O(n8772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_20 (.CI(n35916), .I0(n8492[17]), .I1(GND_net), .CO(n35917));
    SB_LUT4 add_4473_19_lut (.I0(GND_net), .I1(n9555[16]), .I2(GND_net), 
            .I3(n36949), .O(n9225[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_9_lut (.I0(GND_net), .I1(n9101[6]), .I2(GND_net), 
            .I3(n36559), .O(n9084[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_19_lut (.I0(GND_net), .I1(n8492[16]), .I2(GND_net), 
            .I3(n35915), .O(n8469[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_20 (.CI(n36744), .I0(n1797[17]), .I1(GND_net), 
            .CO(n36745));
    SB_CARRY add_4463_9 (.CI(n36559), .I0(n9101[6]), .I1(GND_net), .CO(n36560));
    SB_CARRY add_4433_19 (.CI(n35915), .I0(n8492[16]), .I1(GND_net), .CO(n35916));
    SB_LUT4 add_4463_8_lut (.I0(GND_net), .I1(n9101[5]), .I2(n728_adj_4054), 
            .I3(n36558), .O(n9084[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_18_lut (.I0(GND_net), .I1(n8492[15]), .I2(GND_net), 
            .I3(n35914), .O(n8469[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_19 (.CI(n36949), .I0(n9555[16]), .I1(GND_net), .CO(n36950));
    SB_CARRY mult_14_add_1217_2 (.CI(GND_net), .I0(n23_adj_4052), .I1(n92), 
            .CO(n36865));
    SB_LUT4 mult_14_add_1211_19_lut (.I0(GND_net), .I1(n1797[16]), .I2(GND_net), 
            .I3(n36743), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_8 (.CI(n36558), .I0(n9101[5]), .I1(n728_adj_4054), 
            .CO(n36559));
    SB_CARRY add_4433_18 (.CI(n35914), .I0(n8492[15]), .I1(GND_net), .CO(n35915));
    SB_LUT4 add_4463_7_lut (.I0(GND_net), .I1(n9101[4]), .I2(n631_adj_4055), 
            .I3(n36557), .O(n9084[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_17_lut (.I0(GND_net), .I1(n8492[14]), .I2(GND_net), 
            .I3(n35913), .O(n8469[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_19 (.CI(n36743), .I0(n1797[16]), .I1(GND_net), 
            .CO(n36744));
    SB_CARRY add_4463_7 (.CI(n36557), .I0(n9101[4]), .I1(n631_adj_4055), 
            .CO(n36558));
    SB_CARRY add_4433_17 (.CI(n35913), .I0(n8492[14]), .I1(GND_net), .CO(n35914));
    SB_LUT4 add_4433_16_lut (.I0(GND_net), .I1(n8492[13]), .I2(GND_net), 
            .I3(n35912), .O(n8469[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_6_lut (.I0(GND_net), .I1(n9101[3]), .I2(n534_adj_4056), 
            .I3(n36556), .O(n9084[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_16 (.CI(n35912), .I0(n8492[13]), .I1(GND_net), .CO(n35913));
    SB_DFF \PID_CONTROLLER.err_prev__i1  (.Q(\PID_CONTROLLER.err_prev[0] ), 
           .C(clk32MHz), .D(n17967));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_add_1216_24_lut (.I0(GND_net), .I1(n1802[21]), .I2(GND_net), 
            .I3(n36863), .O(n1801[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_18_lut (.I0(GND_net), .I1(n1797[15]), .I2(GND_net), 
            .I3(n36742), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_6 (.CI(n36556), .I0(n9101[3]), .I1(n534_adj_4056), 
            .CO(n36557));
    SB_LUT4 add_4433_15_lut (.I0(GND_net), .I1(n8492[12]), .I2(GND_net), 
            .I3(n35911), .O(n8469[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n76[0]), 
            .CO(n34673));
    SB_LUT4 add_4463_5_lut (.I0(GND_net), .I1(n9101[2]), .I2(n437_adj_4057), 
            .I3(n36555), .O(n9084[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_15 (.CI(n35911), .I0(n8492[12]), .I1(GND_net), .CO(n35912));
    SB_LUT4 add_4433_14_lut (.I0(GND_net), .I1(n8492[11]), .I2(GND_net), 
            .I3(n35910), .O(n8469[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_18 (.CI(n36742), .I0(n1797[15]), .I1(GND_net), 
            .CO(n36743));
    SB_CARRY add_4463_5 (.CI(n36555), .I0(n9101[2]), .I1(n437_adj_4057), 
            .CO(n36556));
    SB_CARRY add_4433_14 (.CI(n35910), .I0(n8492[11]), .I1(GND_net), .CO(n35911));
    SB_LUT4 add_4463_4_lut (.I0(GND_net), .I1(n9101[1]), .I2(n340_adj_4058), 
            .I3(n36554), .O(n9084[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_13_lut (.I0(GND_net), .I1(n8492[10]), .I2(GND_net), 
            .I3(n35909), .O(n8469[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_18_lut (.I0(GND_net), .I1(n9555[15]), .I2(GND_net), 
            .I3(n36948), .O(n9225[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_24 (.CI(n36863), .I0(n1802[21]), .I1(GND_net), 
            .CO(n1703));
    SB_LUT4 mult_14_add_1211_17_lut (.I0(GND_net), .I1(n1797[14]), .I2(GND_net), 
            .I3(n36741), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_4 (.CI(n36554), .I0(n9101[1]), .I1(n340_adj_4058), 
            .CO(n36555));
    SB_CARRY add_4450_4 (.CI(n36281), .I0(n8802[1]), .I1(n301_adj_4053), 
            .CO(n36282));
    SB_LUT4 add_4450_3_lut (.I0(GND_net), .I1(n8802[0]), .I2(n204_adj_4059), 
            .I3(n36280), .O(n8772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_13 (.CI(n35909), .I0(n8492[10]), .I1(GND_net), .CO(n35910));
    SB_LUT4 add_4433_12_lut (.I0(GND_net), .I1(n8492[9]), .I2(GND_net), 
            .I3(n35908), .O(n8469[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_3 (.CI(n36280), .I0(n8802[0]), .I1(n204_adj_4059), 
            .CO(n36281));
    SB_CARRY add_4433_12 (.CI(n35908), .I0(n8492[9]), .I1(GND_net), .CO(n35909));
    SB_LUT4 add_4450_2_lut (.I0(GND_net), .I1(n14_adj_4060), .I2(n107_adj_4061), 
            .I3(GND_net), .O(n8772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4450_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_23_lut (.I0(GND_net), .I1(n1802[20]), .I2(GND_net), 
            .I3(n36862), .O(n1801[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_17 (.CI(n36741), .I0(n1797[14]), .I1(GND_net), 
            .CO(n36742));
    SB_LUT4 add_4433_11_lut (.I0(GND_net), .I1(n8492[8]), .I2(GND_net), 
            .I3(n35907), .O(n8469[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_3_lut (.I0(GND_net), .I1(n9101[0]), .I2(n243_adj_4062), 
            .I3(n36553), .O(n9084[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4450_2 (.CI(GND_net), .I0(n14_adj_4060), .I1(n107_adj_4061), 
            .CO(n36280));
    SB_LUT4 add_4449_30_lut (.I0(GND_net), .I1(n8772[27]), .I2(GND_net), 
            .I3(n36279), .O(n8741[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_11 (.CI(n35907), .I0(n8492[8]), .I1(GND_net), .CO(n35908));
    SB_LUT4 add_4433_10_lut (.I0(GND_net), .I1(n8492[7]), .I2(GND_net), 
            .I3(n35906), .O(n8469[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_16_lut (.I0(GND_net), .I1(n1797[13]), .I2(GND_net), 
            .I3(n36740), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4463_3 (.CI(n36553), .I0(n9101[0]), .I1(n243_adj_4062), 
            .CO(n36554));
    SB_LUT4 add_4449_29_lut (.I0(GND_net), .I1(n8772[26]), .I2(GND_net), 
            .I3(n36278), .O(n8741[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_29 (.CI(n36278), .I0(n8772[26]), .I1(GND_net), .CO(n36279));
    SB_CARRY add_4433_10 (.CI(n35906), .I0(n8492[7]), .I1(GND_net), .CO(n35907));
    SB_LUT4 add_4433_9_lut (.I0(GND_net), .I1(n8492[6]), .I2(GND_net), 
            .I3(n35905), .O(n8469[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4463_2_lut (.I0(GND_net), .I1(n53_adj_4063), .I2(n146_adj_4064), 
            .I3(GND_net), .O(n9084[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4463_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_28_lut (.I0(GND_net), .I1(n8772[25]), .I2(GND_net), 
            .I3(n36277), .O(n8741[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_28 (.CI(n36277), .I0(n8772[25]), .I1(GND_net), .CO(n36278));
    SB_CARRY add_4433_9 (.CI(n35905), .I0(n8492[6]), .I1(GND_net), .CO(n35906));
    SB_LUT4 add_4433_8_lut (.I0(GND_net), .I1(n8492[5]), .I2(n710_adj_4065), 
            .I3(n35904), .O(n8469[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_8 (.CI(n35904), .I0(n8492[5]), .I1(n710_adj_4065), 
            .CO(n35905));
    SB_CARRY mult_14_add_1216_23 (.CI(n36862), .I0(n1802[20]), .I1(GND_net), 
            .CO(n36863));
    SB_CARRY add_4463_2 (.CI(GND_net), .I0(n53_adj_4063), .I1(n146_adj_4064), 
            .CO(n36553));
    SB_CARRY mult_14_add_1211_16 (.CI(n36740), .I0(n1797[13]), .I1(GND_net), 
            .CO(n36741));
    SB_LUT4 add_4449_27_lut (.I0(GND_net), .I1(n8772[24]), .I2(GND_net), 
            .I3(n36276), .O(n8741[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_17_lut (.I0(GND_net), .I1(n9084[14]), .I2(GND_net), 
            .I3(n36552), .O(n9066[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_16_lut (.I0(GND_net), .I1(n9084[13]), .I2(GND_net), 
            .I3(n36551), .O(n9066[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4433_7_lut (.I0(GND_net), .I1(n8492[4]), .I2(n613_adj_4066), 
            .I3(n35903), .O(n8469[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_27 (.CI(n36276), .I0(n8772[24]), .I1(GND_net), .CO(n36277));
    SB_LUT4 add_4449_26_lut (.I0(GND_net), .I1(n8772[23]), .I2(GND_net), 
            .I3(n36275), .O(n8741[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_7 (.CI(n35903), .I0(n8492[4]), .I1(n613_adj_4066), 
            .CO(n35904));
    SB_LUT4 add_4433_6_lut (.I0(GND_net), .I1(n8492[3]), .I2(n516_adj_4067), 
            .I3(n35902), .O(n8469[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_16 (.CI(n36551), .I0(n9084[13]), .I1(GND_net), .CO(n36552));
    SB_CARRY add_4449_26 (.CI(n36275), .I0(n8772[23]), .I1(GND_net), .CO(n36276));
    SB_LUT4 add_4449_25_lut (.I0(GND_net), .I1(n8772[22]), .I2(GND_net), 
            .I3(n36274), .O(n8741[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4433_6 (.CI(n35902), .I0(n8492[3]), .I1(n516_adj_4067), 
            .CO(n35903));
    SB_LUT4 add_4433_5_lut (.I0(GND_net), .I1(n8492[2]), .I2(n419_adj_4068), 
            .I3(n35901), .O(n8469[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_25 (.CI(n36274), .I0(n8772[22]), .I1(GND_net), .CO(n36275));
    SB_CARRY add_4433_5 (.CI(n35901), .I0(n8492[2]), .I1(n419_adj_4068), 
            .CO(n35902));
    SB_LUT4 i39803_3_lut (.I0(n48426), .I1(pwm_23__N_3310[7]), .I2(n15), 
            .I3(GND_net), .O(n47706));   // verilog/motorControl.v(44[31:51])
    defparam i39803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_17_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(n57[31]), 
            .I3(n34672), .O(pwm_23__N_3310[24])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n57[31]), 
            .I3(n34671), .O(pwm_23__N_3310[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_18 (.CI(n36948), .I0(n9555[15]), .I1(GND_net), .CO(n36949));
    SB_LUT4 add_4433_4_lut (.I0(GND_net), .I1(n8492[1]), .I2(n322_adj_4070), 
            .I3(n35900), .O(n8469[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_22_lut (.I0(GND_net), .I1(n1802[19]), .I2(GND_net), 
            .I3(n36861), .O(n1801[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_15_lut (.I0(GND_net), .I1(n1797[12]), .I2(GND_net), 
            .I3(n36739), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_15_lut (.I0(GND_net), .I1(n9084[12]), .I2(GND_net), 
            .I3(n36550), .O(n9066[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_24_lut (.I0(GND_net), .I1(n8772[21]), .I2(GND_net), 
            .I3(n36273), .O(n8741[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_24 (.CI(n36273), .I0(n8772[21]), .I1(GND_net), .CO(n36274));
    SB_CARRY add_4433_4 (.CI(n35900), .I0(n8492[1]), .I1(n322_adj_4070), 
            .CO(n35901));
    SB_LUT4 add_4433_3_lut (.I0(GND_net), .I1(n8492[0]), .I2(n225_adj_4071), 
            .I3(n35899), .O(n8469[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_15 (.CI(n36739), .I0(n1797[12]), .I1(GND_net), 
            .CO(n36740));
    SB_CARRY add_4462_15 (.CI(n36550), .I0(n9084[12]), .I1(GND_net), .CO(n36551));
    SB_LUT4 add_4449_23_lut (.I0(GND_net), .I1(n8772[20]), .I2(GND_net), 
            .I3(n36272), .O(n8741[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_23 (.CI(n36272), .I0(n8772[20]), .I1(GND_net), .CO(n36273));
    SB_CARRY add_4433_3 (.CI(n35899), .I0(n8492[0]), .I1(n225_adj_4071), 
            .CO(n35900));
    SB_LUT4 add_4433_2_lut (.I0(GND_net), .I1(n35_adj_4072), .I2(n128_adj_4073), 
            .I3(GND_net), .O(n8469[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4433_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_22_lut (.I0(GND_net), .I1(n8772[19]), .I2(GND_net), 
            .I3(n36271), .O(n8741[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_22 (.CI(n36861), .I0(n1802[19]), .I1(GND_net), 
            .CO(n36862));
    SB_CARRY unary_minus_17_add_3_25 (.CI(n34671), .I0(GND_net), .I1(n57[31]), 
            .CO(n34672));
    SB_LUT4 add_4462_14_lut (.I0(GND_net), .I1(n9084[11]), .I2(GND_net), 
            .I3(n36549), .O(n9066[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_22 (.CI(n36271), .I0(n8772[19]), .I1(GND_net), .CO(n36272));
    SB_CARRY add_4433_2 (.CI(GND_net), .I0(n35_adj_4072), .I1(n128_adj_4073), 
            .CO(n35899));
    SB_LUT4 add_4473_17_lut (.I0(GND_net), .I1(n9555[14]), .I2(GND_net), 
            .I3(n36947), .O(n9225[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n57[22]), 
            .I3(n34670), .O(pwm_23__N_3310[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_14_lut (.I0(GND_net), .I1(n1797[11]), .I2(GND_net), 
            .I3(n36738), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_23_lut (.I0(GND_net), .I1(n8469[20]), .I2(GND_net), 
            .I3(n35898), .O(n8445[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_21_lut (.I0(GND_net), .I1(n8772[18]), .I2(GND_net), 
            .I3(n36270), .O(n8741[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_22_lut (.I0(GND_net), .I1(n8469[19]), .I2(GND_net), 
            .I3(n35897), .O(n8445[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_17 (.CI(n36947), .I0(n9555[14]), .I1(GND_net), .CO(n36948));
    SB_CARRY add_4462_14 (.CI(n36549), .I0(n9084[11]), .I1(GND_net), .CO(n36550));
    SB_LUT4 mult_14_add_1216_21_lut (.I0(GND_net), .I1(n1802[18]), .I2(GND_net), 
            .I3(n36860), .O(n1801[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_22 (.CI(n35897), .I0(n8469[19]), .I1(GND_net), .CO(n35898));
    SB_LUT4 add_4473_16_lut (.I0(GND_net), .I1(n9555[13]), .I2(GND_net), 
            .I3(n36946), .O(n9225[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_24 (.CI(n34670), .I0(GND_net), .I1(n57[22]), 
            .CO(n34671));
    SB_CARRY add_4473_16 (.CI(n36946), .I0(n9555[13]), .I1(GND_net), .CO(n36947));
    SB_LUT4 unary_minus_17_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n57[21]), 
            .I3(n34669), .O(pwm_23__N_3310[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_21 (.CI(n36860), .I0(n1802[18]), .I1(GND_net), 
            .CO(n36861));
    SB_LUT4 mult_14_add_1216_20_lut (.I0(GND_net), .I1(n1802[17]), .I2(GND_net), 
            .I3(n36859), .O(n1801[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_21 (.CI(n36270), .I0(n8772[18]), .I1(GND_net), .CO(n36271));
    SB_CARRY unary_minus_17_add_3_23 (.CI(n34669), .I0(GND_net), .I1(n57[21]), 
            .CO(n34670));
    SB_CARRY mult_14_add_1211_14 (.CI(n36738), .I0(n1797[11]), .I1(GND_net), 
            .CO(n36739));
    SB_LUT4 add_4432_21_lut (.I0(GND_net), .I1(n8469[18]), .I2(GND_net), 
            .I3(n35896), .O(n8445[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n57[20]), 
            .I3(n34668), .O(pwm_23__N_3310[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_13_lut (.I0(GND_net), .I1(n9084[10]), .I2(GND_net), 
            .I3(n36548), .O(n9066[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_20_lut (.I0(GND_net), .I1(n8772[17]), .I2(GND_net), 
            .I3(n36269), .O(n8741[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_21 (.CI(n35896), .I0(n8469[18]), .I1(GND_net), .CO(n35897));
    SB_LUT4 add_4432_20_lut (.I0(GND_net), .I1(n8469[17]), .I2(GND_net), 
            .I3(n35895), .O(n8445[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_20 (.CI(n36269), .I0(n8772[17]), .I1(GND_net), .CO(n36270));
    SB_CARRY unary_minus_17_add_3_22 (.CI(n34668), .I0(GND_net), .I1(n57[20]), 
            .CO(n34669));
    SB_CARRY add_4432_20 (.CI(n35895), .I0(n8469[17]), .I1(GND_net), .CO(n35896));
    SB_LUT4 unary_minus_17_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n57[19]), 
            .I3(n34667), .O(pwm_23__N_3310[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_19_lut (.I0(GND_net), .I1(n8469[16]), .I2(GND_net), 
            .I3(n35894), .O(n8445[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_21 (.CI(n34667), .I0(GND_net), .I1(n57[19]), 
            .CO(n34668));
    SB_CARRY add_4462_13 (.CI(n36548), .I0(n9084[10]), .I1(GND_net), .CO(n36549));
    SB_LUT4 add_4449_19_lut (.I0(GND_net), .I1(n8772[16]), .I2(GND_net), 
            .I3(n36268), .O(n8741[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_19 (.CI(n35894), .I0(n8469[16]), .I1(GND_net), .CO(n35895));
    SB_CARRY add_4449_19 (.CI(n36268), .I0(n8772[16]), .I1(GND_net), .CO(n36269));
    SB_CARRY mult_14_add_1216_20 (.CI(n36859), .I0(n1802[17]), .I1(GND_net), 
            .CO(n36860));
    SB_LUT4 add_4462_12_lut (.I0(GND_net), .I1(n9084[9]), .I2(GND_net), 
            .I3(n36547), .O(n9066[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_18_lut (.I0(GND_net), .I1(n8469[15]), .I2(GND_net), 
            .I3(n35893), .O(n8445[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_18_lut (.I0(GND_net), .I1(n8772[15]), .I2(GND_net), 
            .I3(n36267), .O(n8741[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4473_15_lut (.I0(GND_net), .I1(n9555[12]), .I2(GND_net), 
            .I3(n36945), .O(n9225[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_18 (.CI(n35893), .I0(n8469[15]), .I1(GND_net), .CO(n35894));
    SB_LUT4 add_4432_17_lut (.I0(GND_net), .I1(n8469[14]), .I2(GND_net), 
            .I3(n35892), .O(n8445[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4473_15 (.CI(n36945), .I0(n9555[12]), .I1(GND_net), .CO(n36946));
    SB_LUT4 unary_minus_17_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n57[18]), 
            .I3(n34666), .O(pwm_23__N_3310[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_19_lut (.I0(GND_net), .I1(n1802[16]), .I2(GND_net), 
            .I3(n36858), .O(n1801[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_20 (.CI(n34666), .I0(GND_net), .I1(n57[18]), 
            .CO(n34667));
    SB_LUT4 mult_14_add_1211_13_lut (.I0(GND_net), .I1(n1797[10]), .I2(GND_net), 
            .I3(n36737), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_17 (.CI(n35892), .I0(n8469[14]), .I1(GND_net), .CO(n35893));
    SB_LUT4 add_4473_14_lut (.I0(GND_net), .I1(n9555[11]), .I2(GND_net), 
            .I3(n36944), .O(n9225[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_12 (.CI(n36547), .I0(n9084[9]), .I1(GND_net), .CO(n36548));
    SB_CARRY mult_14_add_1216_19 (.CI(n36858), .I0(n1802[16]), .I1(GND_net), 
            .CO(n36859));
    SB_CARRY mult_14_add_1211_13 (.CI(n36737), .I0(n1797[10]), .I1(GND_net), 
            .CO(n36738));
    SB_LUT4 add_4432_16_lut (.I0(GND_net), .I1(n8469[13]), .I2(GND_net), 
            .I3(n35891), .O(n8445[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_11_lut (.I0(GND_net), .I1(n9084[8]), .I2(GND_net), 
            .I3(n36546), .O(n9066[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_18_lut (.I0(GND_net), .I1(n1802[15]), .I2(GND_net), 
            .I3(n36857), .O(n1801[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4462_11 (.CI(n36546), .I0(n9084[8]), .I1(GND_net), .CO(n36547));
    SB_LUT4 mult_14_add_1211_12_lut (.I0(GND_net), .I1(n1797[9]), .I2(GND_net), 
            .I3(n36736), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4462_10_lut (.I0(GND_net), .I1(n9084[7]), .I2(GND_net), 
            .I3(n36545), .O(n9066[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_18 (.CI(n36267), .I0(n8772[15]), .I1(GND_net), .CO(n36268));
    SB_CARRY add_4462_10 (.CI(n36545), .I0(n9084[7]), .I1(GND_net), .CO(n36546));
    SB_LUT4 add_4462_9_lut (.I0(GND_net), .I1(n9084[6]), .I2(GND_net), 
            .I3(n36544), .O(n9066[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4462_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4432_16 (.CI(n35891), .I0(n8469[13]), .I1(GND_net), .CO(n35892));
    SB_LUT4 add_4449_17_lut (.I0(GND_net), .I1(n8772[14]), .I2(GND_net), 
            .I3(n36266), .O(n8741[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_15_lut (.I0(GND_net), .I1(n8469[12]), .I2(GND_net), 
            .I3(n35890), .O(n8445[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_17 (.CI(n36266), .I0(n8772[14]), .I1(GND_net), .CO(n36267));
    SB_CARRY add_4432_15 (.CI(n35890), .I0(n8469[12]), .I1(GND_net), .CO(n35891));
    SB_LUT4 add_4449_16_lut (.I0(GND_net), .I1(n8772[13]), .I2(GND_net), 
            .I3(n36265), .O(n8741[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4432_14_lut (.I0(GND_net), .I1(n8469[11]), .I2(GND_net), 
            .I3(n35889), .O(n8445[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4432_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_18 (.CI(n36857), .I0(n1802[15]), .I1(GND_net), 
            .CO(n36858));
    SB_CARRY add_4473_14 (.CI(n36944), .I0(n9555[11]), .I1(GND_net), .CO(n36945));
    SB_CARRY add_4449_16 (.CI(n36265), .I0(n8772[13]), .I1(GND_net), .CO(n36266));
    SB_LUT4 mult_14_i291_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[3]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i207_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_3507));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i272_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n404));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(n878), .I3(n17_adj_3860), 
            .O(GATES_5__N_3138[0]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2044;
    SB_LUT4 i5_4_lut_adj_848 (.I0(Kd_delay_counter[5]), .I1(Kd_delay_counter[3]), 
            .I2(Kd_delay_counter[6]), .I3(Kd_delay_counter[4]), .O(n12_adj_4079));   // verilog/motorControl.v(56[10:29])
    defparam i5_4_lut_adj_848.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_849 (.I0(Kd_delay_counter[1]), .I1(n12_adj_4079), 
            .I2(Kd_delay_counter[2]), .I3(Kd_delay_counter[0]), .O(n43362));   // verilog/motorControl.v(56[10:29])
    defparam i6_4_lut_adj_849.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i227_2_lut (.I0(\Kd[3] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i461_2_lut (.I0(\Kd[7] ), .I1(n58[2]), .I2(GND_net), 
            .I3(GND_net), .O(n686));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i292_2_lut (.I0(\Kd[4] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n434));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i6_3_lut_3_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n67[3]), 
            .I2(n67[2]), .I3(GND_net), .O(n6_adj_3715));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i39216_3_lut_4_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n67[3]), 
            .I2(n67[2]), .I3(\PID_CONTROLLER.result [2]), .O(n47118));   // verilog/motorControl.v(47[21:37])
    defparam i39216_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_12_i357_2_lut (.I0(\Kd[5] ), .I1(n58[15]), .I2(GND_net), 
            .I3(GND_net), .O(n531));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i337_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n501));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n598));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[18]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[19]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[20]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[21]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[22]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i87_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n128_adj_4073));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4072));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i152_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n225_adj_4071));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_850 (.I0(pwm_23__N_3307), .I1(n1_adj_3675), .I2(PWMLimit[4]), 
            .I3(n387), .O(n18625));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_850.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_851 (.I0(pwm_23__N_3307), .I1(n1_adj_3674), .I2(PWMLimit[6]), 
            .I3(n387), .O(n18627));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_851.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i217_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n322_adj_4070));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i32_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[31]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_852 (.I0(pwm_23__N_3307), .I1(n1), .I2(PWMLimit[10]), 
            .I3(n387), .O(n18631));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_852.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i282_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n419_adj_4068));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n516_adj_4067));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n613_adj_4066));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i477_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n710_adj_4065));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i99_2_lut (.I0(\Kd[1] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n146_adj_4064));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i36_2_lut (.I0(\Kd[0] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4063));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_853 (.I0(pwm_23__N_3307), .I1(n23155), .I2(PWMLimit[13]), 
            .I3(n387), .O(n18634));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_853.LUT_INIT = 16'ha088;
    SB_LUT4 mult_12_i164_2_lut (.I0(\Kd[2] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n243_adj_4062));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i73_2_lut (.I0(\Kd[1] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4061));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i10_2_lut (.I0(\Kd[0] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4060));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i138_2_lut (.I0(\Kd[2] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n204_adj_4059));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i229_2_lut (.I0(\Kd[3] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n340_adj_4058));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_854 (.I0(pwm_23__N_3307), .I1(n23686), .I2(PWMLimit[17]), 
            .I3(n387), .O(n18638));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_854.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_855 (.I0(pwm_23__N_3307), .I1(n23926), .I2(PWMLimit[19]), 
            .I3(n387), .O(n18640));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_855.LUT_INIT = 16'ha088;
    SB_LUT4 mult_12_i294_2_lut (.I0(\Kd[4] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n437_adj_4057));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_856 (.I0(\PID_CONTROLLER.result [29]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(pwm_23__N_3310[24]), .I3(\PID_CONTROLLER.result [25]), .O(n43808));   // verilog/motorControl.v(44[31:51])
    defparam i2_4_lut_adj_856.LUT_INIT = 16'h7ffe;
    SB_LUT4 i3_4_lut_adj_857 (.I0(\PID_CONTROLLER.result [27]), .I1(n43808), 
            .I2(pwm_23__N_3310[24]), .I3(\PID_CONTROLLER.result [24]), .O(n8_adj_4080));   // verilog/motorControl.v(44[31:51])
    defparam i3_4_lut_adj_857.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_4_lut (.I0(\PID_CONTROLLER.result [28]), .I1(n8_adj_4080), 
            .I2(\PID_CONTROLLER.result [30]), .I3(pwm_23__N_3310[24]), .O(n43813));   // verilog/motorControl.v(44[31:51])
    defparam i4_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 mult_12_i359_2_lut (.I0(\Kd[5] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n534_adj_4056));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_833_i15_2_lut (.I0(\PID_CONTROLLER.result [7]), .I1(pwm_23__N_3310[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_833_i11_2_lut (.I0(\PID_CONTROLLER.result [5]), .I1(pwm_23__N_3310[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4081));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i424_2_lut (.I0(\Kd[6] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n631_adj_4055));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_833_i4_3_lut (.I0(n46520), .I1(pwm_23__N_3310[1]), 
            .I2(\PID_CONTROLLER.result [1]), .I3(GND_net), .O(n4_adj_4082));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40522_3_lut (.I0(n4_adj_4082), .I1(pwm_23__N_3310[5]), .I2(n11_adj_4081), 
            .I3(GND_net), .O(n48425));   // verilog/motorControl.v(44[31:51])
    defparam i40522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40523_3_lut (.I0(n48425), .I1(\pwm_23__N_3310[6] ), .I2(n13_adj_11), 
            .I3(GND_net), .O(n48426));   // verilog/motorControl.v(44[31:51])
    defparam i40523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40058_4_lut (.I0(n13_adj_11), .I1(n11_adj_4081), .I2(n9_adj_12), 
            .I3(n47225), .O(n47961));
    defparam i40058_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 pwm_23__I_833_i8_3_lut (.I0(n6_adj_4085), .I1(\pwm_23__N_3310[4] ), 
            .I2(n9_adj_12), .I3(GND_net), .O(n8));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i489_2_lut (.I0(\Kd[7] ), .I1(n58[16]), .I2(GND_net), 
            .I3(GND_net), .O(n728_adj_4054));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i203_2_lut (.I0(\Kd[3] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n301_adj_4053));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4052));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[0]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4049));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i268_2_lut (.I0(\Kd[4] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n398_adj_4048));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i333_2_lut (.I0(\Kd[5] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n495_adj_4047));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i398_2_lut (.I0(\Kd[6] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n592_adj_4046));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i463_2_lut (.I0(\Kd[7] ), .I1(n58[3]), .I2(GND_net), 
            .I3(GND_net), .O(n689_adj_4045));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39259_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(PWMLimit[2]), .O(n47161));   // verilog/motorControl.v(45[12:27])
    defparam i39259_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_12_i101_2_lut (.I0(\Kd[1] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n149_adj_4044));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i38_2_lut (.I0(\Kd[0] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4043));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4042));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_4041));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4040));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i166_2_lut (.I0(\Kd[2] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n246_adj_4039));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i154_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n228_adj_4038));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i231_2_lut (.I0(\Kd[3] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n343_adj_4037));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i219_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n325_adj_4036));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i296_2_lut (.I0(\Kd[4] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n440_adj_4035));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i284_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n422_adj_4034));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4033));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i361_2_lut (.I0(\Kd[5] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n537_adj_4032));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[1]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4029));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i426_2_lut (.I0(\Kd[6] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n634_adj_4028));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n519_adj_4027));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i491_2_lut (.I0(\Kd[7] ), .I1(n58[17]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4026));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[0]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n616_adj_4024));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4023));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[2]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4020));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[1]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4018));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4017));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i479_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n713_adj_4016));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[2]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i150_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n222));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[3]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[3]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i103_2_lut (.I0(\Kd[1] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n152_adj_4011));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i40_2_lut (.I0(\Kd[0] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59_adj_4010));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i75_2_lut (.I0(\Kd[1] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4009));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i12_2_lut (.I0(\Kd[0] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4008));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28766_4_lut_4_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n34094), .I3(n9577[0]), .O(n4_adj_3646));   // verilog/motorControl.v(43[17:23])
    defparam i28766_4_lut_4_lut_4_lut.LUT_INIT = 16'hfa80;
    SB_LUT4 mult_12_i140_2_lut (.I0(\Kd[2] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n207_adj_4007));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[4]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[4]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[5]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i168_2_lut (.I0(\Kd[2] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n249_adj_4002));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i233_2_lut (.I0(\Kd[3] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n346_adj_4001));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i205_2_lut (.I0(\Kd[3] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n304_adj_4000));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[5]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[6]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i298_2_lut (.I0(\Kd[4] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n443_adj_3996));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i270_2_lut (.I0(\Kd[4] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n401_adj_3995));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28710_4_lut_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n34094), .I3(n9577[0]), .O(n4_adj_3644));   // verilog/motorControl.v(43[17:23])
    defparam i28710_4_lut_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_12_i335_2_lut (.I0(\Kd[5] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n498_adj_3994));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[6]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[7]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i363_2_lut (.I0(\Kd[5] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n540_adj_3990));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i400_2_lut (.I0(\Kd[6] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n595_adj_3989));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[7]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[8]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i465_2_lut (.I0(\Kd[7] ), .I1(n58[4]), .I2(GND_net), 
            .I3(GND_net), .O(n692_adj_3985));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i91_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n134_adj_3984));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3983));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i156_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n231_adj_3982));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i428_2_lut (.I0(\Kd[6] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n637_adj_3981));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i493_2_lut (.I0(\Kd[7] ), .I1(n58[18]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_3980));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i221_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n328_adj_3979));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[8]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[9]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i286_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n425_adj_3975));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[10]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[9]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[11]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[10]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n522_adj_3968));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[12]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[11]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n619_adj_3964));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[13]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[14]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[12]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i481_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n716_adj_3959));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[15]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[16]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[13]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[17]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[18]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[14]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[19]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[15]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[20]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[21]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i105_2_lut (.I0(\Kd[1] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n155_adj_3945));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i42_2_lut (.I0(\Kd[0] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_3944));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[22]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[16]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39322_3_lut_4_lut (.I0(\PID_CONTROLLER.result [3]), .I1(pwm_23__N_3310[3]), 
            .I2(pwm_23__N_3310[2]), .I3(\PID_CONTROLLER.result [2]), .O(n47225));   // verilog/motorControl.v(44[31:51])
    defparam i39322_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 pwm_23__I_833_i6_3_lut_3_lut (.I0(\PID_CONTROLLER.result [3]), 
            .I1(pwm_23__N_3310[3]), .I2(pwm_23__N_3310[2]), .I3(GND_net), 
            .O(n6_adj_4085));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_833_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[17]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[18]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[23]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i170_2_lut (.I0(\Kd[2] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n252_adj_3935));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i235_2_lut (.I0(\Kd[3] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n349_adj_3934));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i300_2_lut (.I0(\Kd[4] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n446_adj_3933));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[19]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i365_2_lut (.I0(\Kd[5] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n543_adj_3930));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i430_2_lut (.I0(\Kd[6] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n640_adj_3929));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i495_2_lut (.I0(\Kd[7] ), .I1(n58[19]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_3928));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n137_adj_3927));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3926));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i77_2_lut (.I0(\Kd[1] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_3925));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i14_2_lut (.I0(\Kd[0] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_3924));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i158_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n234_adj_3923));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i223_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_3922));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i142_2_lut (.I0(\Kd[2] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n210_adj_3921));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i288_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n428_adj_3920));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i207_2_lut (.I0(\Kd[3] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n307_adj_3919));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i272_2_lut (.I0(\Kd[4] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n404_adj_3918));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i337_2_lut (.I0(\Kd[5] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n501_adj_3917));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n525_adj_3916));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i402_2_lut (.I0(\Kd[6] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n598_adj_3915));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n622_adj_3914));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i467_2_lut (.I0(\Kd[7] ), .I1(n58[5]), .I2(GND_net), 
            .I3(GND_net), .O(n695_adj_3913));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i483_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n719_adj_3912));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i107_2_lut (.I0(\Kd[1] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n158_adj_3911));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i44_2_lut (.I0(\Kd[0] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n65_adj_3910));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i172_2_lut (.I0(\Kd[2] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n255_adj_3909));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n64[0]));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n282[0]));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[20]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i237_2_lut (.I0(\Kd[3] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n352_adj_3904));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i302_2_lut (.I0(\Kd[4] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n449_adj_3903));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_4_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4086));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i367_2_lut (.I0(\Kd[5] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n546_adj_3902));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i432_2_lut (.I0(\Kd[6] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n643_adj_3901));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i497_2_lut (.I0(\Kd[7] ), .I1(n58[20]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_3900));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i109_2_lut (.I0(\Kd[1] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n161_adj_3899));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i46_2_lut (.I0(\Kd[0] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_3898));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\Kd[3] ), .I1(n58[25]), .I2(n4_adj_3668), 
            .I3(n9584[1]), .O(n9618[2]));   // verilog/motorControl.v(43[26:45])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_12_i174_2_lut (.I0(\Kd[2] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n258_adj_3897));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_3896));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3895));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i239_2_lut (.I0(\Kd[3] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n355_adj_3894));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3893));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[21]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3889));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i304_2_lut (.I0(\Kd[4] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n452_adj_3887));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3886));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i369_2_lut (.I0(\Kd[5] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n549_adj_3884));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24_4_lut (.I0(GATES_5__N_3398[4]), .I1(\GATES_5__N_3398[5] ), 
            .I2(n17_adj_3860), .I3(n878), .O(GATES_5__N_3138[5]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i24_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i2_4_lut_adj_858 (.I0(hall1), .I1(\GATES_5__N_3398[5] ), .I2(hall2), 
            .I3(hall3), .O(GATES_5__N_3398[4]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_4_lut_adj_858.LUT_INIT = 16'h1050;
    SB_LUT4 GATES_5__I_0_i5_4_lut (.I0(n878), .I1(GATES_5__N_3398[4]), .I2(n17_adj_3860), 
            .I3(\GATES_5__N_3398[5] ), .O(GATES_5__N_3138[4]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i5_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i3_4_lut_adj_859 (.I0(pwm_count[8]), .I1(n865), .I2(n868), 
            .I3(n16), .O(n19_adj_4088));
    defparam i3_4_lut_adj_859.LUT_INIT = 16'h0223;
    SB_LUT4 i36418_3_lut (.I0(n866), .I1(n44276), .I2(n853), .I3(GND_net), 
            .O(n44318));
    defparam i36418_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i36414_4_lut (.I0(n862), .I1(n864), .I2(n859), .I3(n861), 
            .O(n44314));
    defparam i36414_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36416_4_lut (.I0(n857), .I1(n856), .I2(n867), .I3(n863), 
            .O(n44316));
    defparam i36416_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_860 (.I0(n44318), .I1(n19_adj_4088), .I2(n855), 
            .I3(n860), .O(n29_adj_4089));
    defparam i13_4_lut_adj_860.LUT_INIT = 16'h0004;
    SB_LUT4 i2_4_lut_adj_861 (.I0(n29_adj_4089), .I1(hall3), .I2(n44316), 
            .I3(n44314), .O(n6_adj_4090));
    defparam i2_4_lut_adj_861.LUT_INIT = 16'h333b;
    SB_LUT4 GATES_5__I_0_i4_4_lut (.I0(n5), .I1(GATES_5__N_3398[3]), .I2(n17_adj_3860), 
            .I3(n6_adj_4090), .O(GATES_5__N_3138[3]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i4_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 i37_3_lut_3_lut (.I0(\PID_CONTROLLER.result [9]), .I1(pwm_23__N_3310[9]), 
            .I2(n18), .I3(GND_net), .O(n29));   // verilog/motorControl.v(44[31:51])
    defparam i37_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i2_3_lut_adj_862 (.I0(hall2), .I1(\GATES_5__N_3398[5] ), .I2(hall3), 
            .I3(GND_net), .O(GATES_5__N_3398[3]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_3_lut_adj_862.LUT_INIT = 16'h0202;
    SB_LUT4 GATES_5__I_0_i3_4_lut (.I0(n46595), .I1(hall2), .I2(n17_adj_3860), 
            .I3(hall3), .O(GATES_5__N_3138[2]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i3_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mult_12_i434_2_lut (.I0(\Kd[6] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n646_adj_3879));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[22]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i95_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n140_adj_3875));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3874));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i499_2_lut (.I0(\Kd[7] ), .I1(n58[21]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_3873));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i160_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n237_adj_3872));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[23]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38950_2_lut_4_lut (.I0(hall2), .I1(\GATES_5__N_3398[5] ), .I2(hall3), 
            .I3(n878), .O(n46595));   // verilog/motorControl.v(86[14] 109[8])
    defparam i38950_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mult_10_i225_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n334_adj_3867));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i1_1_lut (.I0(\PID_CONTROLLER.err[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[0]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i290_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n431_adj_3864));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3863));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i79_2_lut (.I0(\Kd[1] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_3862));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i16_2_lut (.I0(\Kd[0] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3861));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3859));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i2_1_lut (.I0(\PID_CONTROLLER.err[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[1]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3851));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n528_adj_3849));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i3_1_lut (.I0(\PID_CONTROLLER.err[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[2]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_adj_3847));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i144_2_lut (.I0(\Kd[2] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n213_adj_3846));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3845));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i4_1_lut (.I0(\PID_CONTROLLER.err[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[3]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i485_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n722_adj_3842));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i5_1_lut (.I0(\PID_CONTROLLER.err[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[4]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i209_2_lut (.I0(\Kd[3] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n310_adj_3840));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i111_2_lut (.I0(\Kd[1] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n164_adj_3839));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i48_2_lut (.I0(\Kd[0] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71_adj_3838));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i274_2_lut (.I0(\Kd[4] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n407_adj_3837));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i339_2_lut (.I0(\Kd[5] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n504_adj_3836));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i176_2_lut (.I0(\Kd[2] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n261_adj_3835));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i6_1_lut (.I0(\PID_CONTROLLER.err[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[5]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_3833));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i404_2_lut (.I0(\Kd[6] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n601_adj_3831));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i241_2_lut (.I0(\Kd[3] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n358_adj_3830));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i7_1_lut (.I0(\PID_CONTROLLER.err[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[6]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i8_1_lut (.I0(\PID_CONTROLLER.err[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[7]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i306_2_lut (.I0(\Kd[4] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n455_adj_3827));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i9_1_lut (.I0(\PID_CONTROLLER.err[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[8]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i469_2_lut (.I0(\Kd[7] ), .I1(n58[6]), .I2(GND_net), 
            .I3(GND_net), .O(n698_adj_3825));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i371_2_lut (.I0(\Kd[5] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n552_adj_3824));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i97_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n143_adj_3823));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3822));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i162_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n240_adj_3821));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i436_2_lut (.I0(\Kd[6] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n649_adj_3820));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3819));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i227_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n337_adj_3816));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i292_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n434_adj_3815));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n531_adj_3814));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n628_adj_3813));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i501_2_lut (.I0(\Kd[7] ), .I1(n58[22]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_3812));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i487_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n725_adj_3811));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i113_2_lut (.I0(\Kd[1] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n167_adj_3810));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i50_2_lut (.I0(\Kd[0] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_3809));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i99_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n146_adj_3808));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3807));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i164_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n243_adj_3806));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i229_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n340));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i294_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n437_adj_3804));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i178_2_lut (.I0(\Kd[2] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n264_adj_3803));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n534));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n631));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i489_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n728));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i243_2_lut (.I0(\Kd[3] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n361_adj_3799));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i308_2_lut (.I0(\Kd[4] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n458_adj_3792));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i101_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n149_adj_3788));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3787));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i166_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n246_adj_3786));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i373_2_lut (.I0(\Kd[5] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n555_adj_3785));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i231_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n343));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n440));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i81_2_lut (.I0(\Kd[1] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_3782));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i18_2_lut (.I0(\Kd[0] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_3781));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i10_1_lut (.I0(\PID_CONTROLLER.err[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[9]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n537_adj_3779));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i11_1_lut (.I0(\PID_CONTROLLER.err[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[10]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i146_2_lut (.I0(\Kd[2] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n216_adj_3777));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i426_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n634));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i438_2_lut (.I0(\Kd[6] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n652_adj_3776));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i491_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i211_2_lut (.I0(\Kd[3] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n313_adj_3773));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i12_1_lut (.I0(\PID_CONTROLLER.err[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[11]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29007_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(n58[25]), 
            .I3(GND_net), .O(n9584[0]));   // verilog/motorControl.v(43[26:45])
    defparam i29007_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i28975_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(\Kd[2] ), 
            .I3(GND_net), .O(n34352));   // verilog/motorControl.v(43[26:45])
    defparam i28975_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(n373), .I1(n4_adj_3668), .I2(n34352), 
            .I3(n58[25]), .O(n7_adj_3670));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6966;
    SB_LUT4 i39183_2_lut_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(n67[21]), 
            .I2(\PID_CONTROLLER.result [9]), .I3(n67[9]), .O(n47085));
    defparam i39183_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i39193_2_lut_4_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n67[16]), 
            .I2(\PID_CONTROLLER.result [7]), .I3(n67[7]), .O(n47095));
    defparam i39193_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i29031_3_lut_4_lut (.I0(n9618[2]), .I1(\Kd[4] ), .I2(n58[25]), 
            .I3(n6_adj_4093), .O(n8_adj_3671));   // verilog/motorControl.v(43[26:45])
    defparam i29031_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 mult_12_i276_2_lut (.I0(\Kd[4] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n410_adj_3771));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i503_2_lut (.I0(\Kd[7] ), .I1(n58[23]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_3770));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i341_2_lut (.I0(\Kd[5] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n507_adj_3769));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i215_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n319));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i13_1_lut (.I0(\PID_CONTROLLER.err[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[12]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i115_2_lut (.I0(\Kd[1] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n170_adj_3767));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i406_2_lut (.I0(\Kd[6] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n604_adj_3766));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i471_2_lut (.I0(\Kd[7] ), .I1(n58[7]), .I2(GND_net), 
            .I3(GND_net), .O(n701_adj_3764));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i180_2_lut (.I0(\Kd[2] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n267));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kd[5] ), .I1(n58[25]), .I2(\Kd[4] ), 
            .I3(n6_adj_4093), .O(n8_adj_3672));   // verilog/motorControl.v(43[26:45])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hb748;
    SB_LUT4 i29023_3_lut_4_lut (.I0(n9584[1]), .I1(\Kd[3] ), .I2(n58[25]), 
            .I3(n4_adj_3668), .O(n6_adj_4093));   // verilog/motorControl.v(43[26:45])
    defparam i29023_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 sub_11_inv_0_i14_1_lut (.I0(\PID_CONTROLLER.err[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[13]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i245_2_lut (.I0(\Kd[3] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n364_adj_3762));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29002_2_lut_3_lut (.I0(\Kd[0] ), .I1(n58[25]), .I2(\Kd[1] ), 
            .I3(GND_net), .O(n34377));   // verilog/motorControl.v(43[26:45])
    defparam i29002_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mult_12_i310_2_lut (.I0(\Kd[4] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n461));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i15_1_lut (.I0(\PID_CONTROLLER.err[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[14]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i103_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n152_adj_3759));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i40_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i375_2_lut (.I0(\Kd[5] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n558));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_863 (.I0(n9618[2]), .I1(\Kd[4] ), .I2(n58[25]), 
            .I3(n6_adj_4093), .O(n9584[3]));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut_adj_863.LUT_INIT = 16'h956a;
    SB_LUT4 mult_10_i168_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n249));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i233_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n346));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n443_adj_3755));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i440_2_lut (.I0(\Kd[6] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n655_adj_3754));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i16_1_lut (.I0(\PID_CONTROLLER.err[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[15]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n540));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i2_2_lut (.I0(\Kd[0] ), .I1(n58[0]), .I2(GND_net), 
            .I3(GND_net), .O(n191[0]));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i505_2_lut (.I0(\Kd[7] ), .I1(n58[24]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_3752));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i428_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n637));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i493_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_3748));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3747));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3746));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i17_1_lut (.I0(\PID_CONTROLLER.err[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[16]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i18_1_lut (.I0(\PID_CONTROLLER.err[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[17]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3743));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i105_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n155_adj_3741));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i170_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n252));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i235_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n349));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i19_1_lut (.I0(\PID_CONTROLLER.err[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[18]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n446));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut (.I0(n19_adj_3972), .I1(n25_adj_3960), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4094));   // verilog/motorControl.v(40[38:63])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n33_adj_3941), .I1(n43_adj_3890), .I2(n27_adj_3955), 
            .I3(n35_adj_3939), .O(n24_adj_4095));   // verilog/motorControl.v(40[38:63])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n41_adj_3905), .I1(n45_adj_3877), .I2(n31_adj_3948), 
            .I3(n23_adj_3965), .O(n22_adj_4096));   // verilog/motorControl.v(40[38:63])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n29_adj_3951), .I1(n24_adj_4095), .I2(n18_adj_4094), 
            .I3(n37_adj_3937), .O(n26_adj_4097));   // verilog/motorControl.v(40[38:63])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_864 (.I0(n21_adj_3969), .I1(n26_adj_4097), .I2(n22_adj_4096), 
            .I3(n39_adj_3931), .O(n43573));   // verilog/motorControl.v(40[38:63])
    defparam i13_4_lut_adj_864.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_4_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(IntegralLimit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4098));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(IntegralLimit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4099));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(IntegralLimit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4100));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40142_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4100), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4099), .O(n48045));
    defparam i40142_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i40140_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[10]), 
            .I2(IntegralLimit[11]), .I3(n48045), .O(n48043));
    defparam i40140_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i39389_4_lut (.I0(n11_adj_3998), .I1(n9_adj_4004), .I2(n7_adj_4013), 
            .I3(n5_adj_4021), .O(n47292));
    defparam i39389_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_4_i13_rep_571_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n50913));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i13_rep_571_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40146_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n50913), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4098), .O(n48049));
    defparam i40146_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i40134_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48049), .O(n48037));
    defparam i40134_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i39403_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47306));
    defparam i39403_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_4_i35_rep_559_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n50901));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i35_rep_559_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4101));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28775_3_lut_4_lut (.I0(n9577[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_3646), .O(n6_adj_3612));   // verilog/motorControl.v(43[17:23])
    defparam i28775_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 LessThan_4_i30_4_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[16]), .O(n30_adj_4102));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_4_i5_2_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(IntegralLimit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4103));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40150_4_lut (.I0(n9_adj_4099), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n5_adj_4103), .I3(IntegralLimit[3]), .O(n48053));
    defparam i40150_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i28698_2_lut_3_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[1] ), .I3(GND_net), .O(n34094));   // verilog/motorControl.v(43[17:23])
    defparam i28698_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i40148_4_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n11_adj_4098), 
            .I2(IntegralLimit[6]), .I3(n48053), .O(n48051));
    defparam i40148_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i39421_4_lut (.I0(n17_adj_4100), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n48051), .I3(IntegralLimit[7]), .O(n47324));
    defparam i39421_4_lut.LUT_INIT = 16'haeab;
    SB_LUT4 i40444_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[9]), 
            .I2(IntegralLimit[10]), .I3(n47324), .O(n48347));
    defparam i40444_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i40912_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[11]), 
            .I2(IntegralLimit[12]), .I3(n48347), .O(n48815));
    defparam i40912_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i40136_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48815), .O(n48039));
    defparam i40136_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_865 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n9577[1]), .I3(n4_adj_3644), .O(n9612[2]));   // verilog/motorControl.v(43[17:23])
    defparam i1_2_lut_3_lut_4_lut_adj_865.LUT_INIT = 16'h8778;
    SB_LUT4 i40703_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48039), .O(n48606));
    defparam i40703_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i41019_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[17]), 
            .I2(IntegralLimit[18]), .I3(n48606), .O(n48922));
    defparam i41019_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i41137_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[19]), 
            .I2(IntegralLimit[20]), .I3(n48922), .O(n49040));
    defparam i41137_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_4_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4104));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39465_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(IntegralLimit[9]), .O(n47368));
    defparam i39465_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 LessThan_4_i24_4_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[21]), .O(n24_adj_4105));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i40544_3_lut (.I0(n6_adj_4104), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48447));   // verilog/motorControl.v(40[10:34])
    defparam i40544_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39395_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[12]), 
            .I2(IntegralLimit[21]), .I3(n48043), .O(n47298));
    defparam i39395_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_4_i45_rep_524_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n50866));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i45_rep_524_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i40560_3_lut (.I0(n24_adj_4105), .I1(n8_adj_4086), .I2(n47368), 
            .I3(GND_net), .O(n48463));   // verilog/motorControl.v(40[10:34])
    defparam i40560_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39777_4_lut (.I0(n48447), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[11]), .O(n47680));   // verilog/motorControl.v(40[10:34])
    defparam i39777_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_6_i4_4_lut (.I0(n75[0]), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3_adj_4030), .I3(\PID_CONTROLLER.integral [0]), .O(n4_adj_4106));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i40536_3_lut (.I0(n4_adj_4106), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n11_adj_3998), .I3(GND_net), .O(n48439));   // verilog/motorControl.v(40[38:63])
    defparam i40536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40537_3_lut (.I0(n48439), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n13_adj_3992), .I3(GND_net), .O(n48440));   // verilog/motorControl.v(40[38:63])
    defparam i40537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i8_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n17_adj_3977), .I3(GND_net), .O(n8_adj_4107));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39383_2_lut (.I0(n17_adj_3977), .I1(n9_adj_4004), .I2(GND_net), 
            .I3(GND_net), .O(n47286));
    defparam i39383_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_6_i6_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n7_adj_4013), .I3(GND_net), .O(n6_adj_4108));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i16_3_lut (.I0(n8_adj_4107), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n43573), .I3(GND_net), .O(n16_adj_4109));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39385_4_lut (.I0(n17_adj_3977), .I1(n15_adj_3987), .I2(n13_adj_3992), 
            .I3(n47292), .O(n47288));
    defparam i39385_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i40687_4_lut (.I0(n16_adj_4109), .I1(n6_adj_4108), .I2(n43573), 
            .I3(n47286), .O(n48590));   // verilog/motorControl.v(40[38:63])
    defparam i40687_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39787_3_lut (.I0(n48440), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n15_adj_3987), .I3(GND_net), .O(n47690));   // verilog/motorControl.v(40[38:63])
    defparam i39787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40988_4_lut (.I0(n47690), .I1(n48590), .I2(n43573), .I3(n47288), 
            .O(n48891));   // verilog/motorControl.v(40[38:63])
    defparam i40988_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_4_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(IntegralLimit[1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), .O(n4_adj_4110));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i40540_3_lut (.I0(n4_adj_4110), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48443));   // verilog/motorControl.v(40[10:34])
    defparam i40540_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39406_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48037), .O(n47309));
    defparam i39406_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i40942_4_lut (.I0(n30_adj_4102), .I1(n10_adj_4101), .I2(n50901), 
            .I3(n47306), .O(n48845));   // verilog/motorControl.v(40[10:34])
    defparam i40942_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39779_4_lut (.I0(n48443), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[14]), .O(n47682));   // verilog/motorControl.v(40[10:34])
    defparam i39779_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i41103_4_lut (.I0(n47682), .I1(n48845), .I2(n50901), .I3(n47309), 
            .O(n49006));   // verilog/motorControl.v(40[10:34])
    defparam i41103_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i41104_3_lut (.I0(n49006), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n49007));   // verilog/motorControl.v(40[10:34])
    defparam i41104_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40122_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(n49040), .O(n48025));
    defparam i40122_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i40829_4_lut (.I0(n47680), .I1(n48463), .I2(n50866), .I3(n47298), 
            .O(n48732));   // verilog/motorControl.v(40[10:34])
    defparam i40829_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39785_4_lut (.I0(n49007), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[19]), .O(n47688));   // verilog/motorControl.v(40[10:34])
    defparam i39785_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i40989_3_lut (.I0(n48891), .I1(n75[23]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48892));   // verilog/motorControl.v(40[38:63])
    defparam i40989_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40986_3_lut (.I0(n47688), .I1(n48732), .I2(n48025), .I3(GND_net), 
            .O(n48889));   // verilog/motorControl.v(40[10:34])
    defparam i40986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_866 (.I0(n48889), .I1(n48892), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[23]), .O(n55_adj_3736));   // verilog/motorControl.v(40[10:63])
    defparam i8_4_lut_adj_866.LUT_INIT = 16'h80c8;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n543));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_3735));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i430_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n640));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i495_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[4] ), 
            .I1(\PID_CONTROLLER.result [8]), .I2(deadband[8]), .I3(GND_net), 
            .O(n8_adj_3542));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 i39345_2_lut_4_lut (.I0(deadband[21]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(deadband[9]), .I3(\PID_CONTROLLER.result [9]), .O(n47248));
    defparam i39345_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i16_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result [21]), .I2(deadband[21]), .I3(GND_net), 
            .O(n16_adj_3540));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i16_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i18_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[10] ), 
            .I1(\PID_CONTROLLER.result [11]), .I2(deadband[11]), .I3(GND_net), 
            .O(n18_adj_3539));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i18_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [2]), 
            .I1(\PID_CONTROLLER.result [3]), .I2(deadband[3]), .I3(GND_net), 
            .O(n6_adj_3538));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [5]), 
            .I1(\PID_CONTROLLER.result[6] ), .I2(deadband[6]), .I3(GND_net), 
            .O(n10_adj_3563));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 i39357_2_lut_4_lut (.I0(deadband[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(deadband[7]), .I3(\PID_CONTROLLER.result [7]), .O(n47260));
    defparam i39357_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i12_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [7]), 
            .I1(\PID_CONTROLLER.result [16]), .I2(deadband[16]), .I3(GND_net), 
            .O(n12_adj_3531));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i12_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_20_i8_3_lut_3_lut (.I0(\PID_CONTROLLER.result[4] ), .I1(\PID_CONTROLLER.result [8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_3512));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39219_2_lut_4_lut (.I0(PWMLimit[21]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(PWMLimit[9]), .I3(\PID_CONTROLLER.result [9]), .O(n47121));
    defparam i39219_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_20_i16_3_lut_3_lut (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result [21]), .I2(PWMLimit[21]), .I3(GND_net), 
            .O(n16_adj_3510));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_11_inv_0_i20_1_lut (.I0(\PID_CONTROLLER.err[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[19]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i83_2_lut (.I0(\Kd[1] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_3725));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i20_2_lut (.I0(\Kd[0] ), .I1(n58[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3724));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i148_2_lut (.I0(\Kd[2] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n219_adj_3718));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i107_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n158));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i44_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n65));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i172_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n255));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i213_2_lut (.I0(\Kd[3] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n316_adj_3714));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i237_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n352));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n449_adj_3713));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i278_2_lut (.I0(\Kd[4] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n413_adj_3712));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i343_2_lut (.I0(\Kd[5] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n510_adj_3710));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n546));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i21_1_lut (.I0(\PID_CONTROLLER.err[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[20]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i408_2_lut (.I0(\Kd[6] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n607_adj_3708));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i432_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n643));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i497_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i10_3_lut_3_lut (.I0(\PID_CONTROLLER.result [5]), 
            .I1(\PID_CONTROLLER.result[6] ), .I2(PWMLimit[6]), .I3(GND_net), 
            .O(n10_adj_3514));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i473_2_lut (.I0(\Kd[7] ), .I1(n58[8]), .I2(GND_net), 
            .I3(GND_net), .O(n704_adj_3704));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i22_1_lut (.I0(\PID_CONTROLLER.err[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[21]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29088_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n34487));   // verilog/motorControl.v(43[17:23])
    defparam i29088_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i28759_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(GND_net), .O(n9577[0]));   // verilog/motorControl.v(43[17:23])
    defparam i28759_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 sub_11_inv_0_i23_1_lut (.I0(\PID_CONTROLLER.err[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[22]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i109_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i46_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n68));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i174_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n258));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39236_2_lut_4_lut (.I0(PWMLimit[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(PWMLimit[7]), .I3(\PID_CONTROLLER.result [7]), .O(n47138));
    defparam i39236_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_20_i12_3_lut_3_lut (.I0(\PID_CONTROLLER.result [7]), 
            .I1(\PID_CONTROLLER.result [16]), .I2(PWMLimit[16]), .I3(GND_net), 
            .O(n12));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_867 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n9577[1]), .I3(n4_adj_3646), .O(n9577[2]));   // verilog/motorControl.v(43[17:23])
    defparam i1_2_lut_3_lut_4_lut_adj_867.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i239_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n355));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i239_2_lut.LUT_INIT = 16'h8888;
    
endmodule
