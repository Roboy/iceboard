// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue May 19 17:48:20 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    
    wire n45509;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(354[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(362[15:20])
    
    wire pwm_setpoint_23__N_183, n209, n211, n61602, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, 
        n260, n261, n262, n263, n264, n265, n266, n267, n268, 
        n269, n270, n296, n330, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n1856, n1854, n356, n62598, n62595, n379, n62592, n20251, 
        n418, n419, n420, n421, n422, n423, n424, n425, n426, 
        n427, n428, n429, n430, n431, n432, n433, n434, n435, 
        n436, n437, n438, n439, n440, n441, n62715;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n62745;
    wire [7:0]commutation_state_7__N_184;
    
    wire commutation_state_7__N_192, n27253, n27252, n40, n30905, 
        GHA_N_331, GLA_N_348, GHB_N_353, GLB_N_362, GHC_N_367, GLC_N_376, 
        dti_N_380, n27251, n27247, n27246, RX_N_2, n1852, n1850, 
        n1848, n1846, n62739, n1844, n1842, n1840;
    wire [31:0]motor_state_23__N_67;
    wire [23:0]displacement_23__N_43;
    
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, 
        n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
        n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
        n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
        read_N_385, n1365, n28, n22, n19, n17, n16, n15, n13, 
        n11, n9, n8, n7, n6, n5, n4, n24, n61887, n62472, 
        n62466, n62463, n1788, n1889, n1891, n1893, n1895, n1897, 
        n1899, n1901, n1903, n1905;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n27245;
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [5:0]color_bit_N_478;
    
    wire n5040, n5039, n5038, n5037, n5036, n5035, n5034, n5032, 
        n5031, n5030, n5029, n5028, n10, n5027, n5026, n5025, 
        n5024, n5023, n27243, n62733, n45561, n27242, n27241, 
        n27240, n27237, n27236, n62020, n19_adj_5685, n17_adj_5686, 
        n16_adj_5687, n15_adj_5688, n13_adj_5689, n11_adj_5690, n2916, 
        n45560, n45508, n61003, n3, n4_adj_5691, n5_adj_5692, n6_adj_5693, 
        n7_adj_5694, n8_adj_5695, n9_adj_5696, n10_adj_5697, n11_adj_5698, 
        n12, n13_adj_5699, n14, n15_adj_5700, n16_adj_5701, n17_adj_5702, 
        n18, n19_adj_5703, n20, n21, n22_adj_5704, n23, n24_adj_5705, 
        n25, n45559, n2, n45558, n14_adj_5706, n15_adj_5707, n16_adj_5708, 
        n17_adj_5709, n18_adj_5710, n19_adj_5711, n20_adj_5712, n21_adj_5713, 
        n22_adj_5714, n23_adj_5715, n24_adj_5716, n25_adj_5717, n27234, 
        n27233, n27232, n27231, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n45557;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n2925, n3543, n5022, n62637, 
        n20312, n27230, n45493, n27228, n27227, n2978, n45507, 
        n45556, n62727, n7_adj_5718, n26384, n52283, n52282, n52281, 
        n52280, n52157, n52279, n52278, n52277, n52276, n52275, 
        n52274, n52273, n52272, n52271, n52270, n52269, n52268, 
        n52267, n52266, n52265, n52264, n52263, n52262, n52261, 
        n52260, n52259, n52258, n52257, n52256, n52161, n52255, 
        n52254, n52253, n52252, n52251, n52250, n26347, n52249, 
        n52248, n52218, n52247, n52246, n52245, n52244, n52243, 
        n52242, n52241, n52224, n52240, n52239, n52238, n52237, 
        n52236, n52235, n52234, n52233, n26327, n52232, n52231, 
        n52230, n52229, n52228, n52227, n52226, n26319, n52156, 
        n26317, n52221, n52222, n52223, n52225, n52160, n52220, 
        n52162, n52163, n52164, n52165, n52166, n52167, n52168, 
        n52169, n26302, n52170, n26300, n52171, n52172, n52173, 
        n52174, n52175, n26294, n52176, n26292, n52177, n52178, 
        n52179, n52180, n52181, n52182, n52183, n26284, n26283, 
        n52184, n26281, n52185, n52186, n52187, n26277, n26276, 
        n26275, n52188, n52189, n52190, n52191, n52192, n52193, 
        n52194, n52195, n52196, n52197, n52198, n52199, n52200, 
        n52201, n52202, n52203, n52204, n52205, n52206, n52207, 
        n52352, n52208, n52209, n52210, n52211, n52212, n26215, 
        n52213, n26213, n52214, n26207, n52216, n51937, n12_adj_5719, 
        n8_adj_5720, n1130, n45555, n45554, n45492, n45506, n45553, 
        n52154, n45552, n45551, n45550, n45505, n45549, n45548, 
        n45504, n45503, n45502, n45547, n45546, n45491, n45545, 
        n45544, n45490, n45501, n45543, n1513, n45542, n45541, 
        n45540, n45489, n45539, n45538, n6_adj_5721, n45537, n45536, 
        n45535, n45534, n2076, n62721, n22887, n37855, n37991, 
        n45533, n37902, n37969, n37857, n62589, n62586, n27226, 
        n27224, n27223, n27222, n4858, n4855, n4847, n7_adj_5722, 
        n6_adj_5723, Kp_23__N_969, n15_adj_5724, n27218, n6_adj_5725, 
        Kp_23__N_675, Kp_23__N_645, n4_adj_5726, n62709, n27213, n22878, 
        n27203, n27200, \FRAME_MATCHER.i_31__N_2485 , Kp_23__N_1724, 
        n15_adj_5727, n15_adj_5728, n27192, n52215, n27148, n27144, 
        n27136, n27133, n27130, n27129, n27128, n27127, n27126, 
        n27124, n27123, n27122, n27121, n27120, n27119, n27118, 
        n27117, n27116, n27115, n27114, n27113, n27112, n27111, 
        n27110, n27109, n27108, n27105, n27104, n27101, n27100, 
        n27099, n27097, n27096, n27095, n27094, n27093, n27092, 
        n27091, n27090, n27089, n27088, n27087, n27086, n27085, 
        n27084, n27083, n27082, n27081, n27080, n27079, n27078, 
        n27062, n27061, n27057, n27056, n27055, n27054, n27053, 
        n27052, n27051, n27050, n27049, n27048, n27047, n27046, 
        n27045, n27044, n27043, n27042, n27041, n27040, n27039, 
        n27038, n27028, n27023, n27022, n27021, n27020, n27019, 
        n27018, n27017, n27016, n27015, n27014, n27010, n27009, 
        n62, n26986, n26985, n26982, n26979, n26978, n26977, n26976, 
        n26975, n26972, n26969, n26968, n26960, n26957, n26956, 
        n26953, n26946, n26944, n26943, n26934, n26932, n26930, 
        n26929, n26925, n26924, n26923, n26922, n26920, n26916, 
        n26915, n51553, n51555, n51557, n51559, n51561, n10_adj_5729, 
        n51563, n51565, n9_adj_5730, n8_adj_5731, n7_adj_5732, n6_adj_5733, 
        n5_adj_5734, n4_adj_5735, n40_adj_5736, n28111, n28105, n32, 
        n24_adj_5737, n19_adj_5738, n17_adj_5739, n16_adj_5740, n15_adj_5741, 
        n13_adj_5742, n11_adj_5743, n9_adj_5744, n8_adj_5745, n7_adj_5746, 
        n6_adj_5747, n5_adj_5748, n4_adj_5749, n28096, n28095, n28093, 
        n4_adj_5750, n3_adj_5751, n28052, n28046, n28044, n27987, 
        n27986, n27985, n27981, n27979, n27978, n27970, n27968, 
        n27962, n27960, n27945, n27935, n52831, n6_adj_5752, n6_adj_5753, 
        n5_adj_5754, n26691, n52309, n53350, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n143, n151, n152, n155, n181, n203, n204, n214, n220;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3691 ;
    
    wire n375, n56666, n56663, n10_adj_5755, n27772, n15_adj_5756, 
        n11_adj_5757, n54562, n52878, n27757, n45532;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, position_31__N_3803, n5021, n5020, n5019, n5018, 
        n5017, n5016, n5015, n5014, n5013, n5012, n5010, n61601;
    wire [1:0]a_new_adj_5900;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5759, position_31__N_3803_adj_5760, n38310, n61189, 
        n26, n25_adj_5761, n24_adj_5762, n23_adj_5763, n4_adj_5764, 
        n3_adj_5765;
    wire [7:0]data_adj_5912;   // verilog/eeprom.v(23[12:16])
    wire [7:0]state_7__N_3892;
    
    wire n24_adj_5766, n62568, n62703, n5057, n5056, n5055, n5054, 
        n5053, n5052, n2_adj_5767, n62079, n27662, n5051, clk_out;
    wire [15:0]data_adj_5920;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_5922;   // verilog/tli4970.v(29[13:18])
    
    wire n27659, n27656, n27653, n27650, n27647, n27644, n27637, 
        n45531, n22771, n45799, n10_adj_5778, n5050, n5049, n5048, 
        n5047, n5046, n5045, n5044, n5043, n5042, n5041, state_7__N_4293, 
        n22915, n45798, n26787, n26786, n22_adj_5779, n21_adj_5780, 
        n27614, n27613, n27612, n27611, n27609, n27608, n27607, 
        n27606, n27605, n27604, n27603, n27602, n27601, n27600, 
        n27599, n27598, n27597, n26782, n6543, n27595, n27594, 
        r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n27593, n27590, n4_adj_5781, n27584, n27583, n27579;
    wire [24:0]o_Rx_DV_N_3464;
    
    wire n62565, n27572, n20_adj_5782, n19_adj_5783, n18_adj_5784, 
        n17_adj_5785, n16_adj_5786, n51551;
    wire [2:0]r_SM_Main_adj_5933;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5934;   // verilog/uart_tx.v(33[16:29])
    
    wire n45797, n45796, n25295, n25293, n45795, n27551, n27549, 
        n27543, n15_adj_5797, n14_adj_5798, n13_adj_5799, n12_adj_5800, 
        n11_adj_5801, n51567, n27524, n27523, n27522, n45530;
    wire [7:0]state_adj_5946;   // verilog/i2c_controller.v(33[12:17])
    
    wire n27521, n52310;
    wire [7:0]counter_adj_5947;   // verilog/i2c_controller.v(36[12:19])
    
    wire enable_slow_N_4187, n27520, n27519, n27518, n10_adj_5803, 
        n9_adj_5804, n8_adj_5805, n7_adj_5806, n27517, n6_adj_5807, 
        n5_adj_5808, n27516, n27515, n27514, n27513, n27512;
    wire [7:0]state_7__N_4084;
    
    wire n27511, n27510, n27509, n27508, n5_adj_5809, n27507, n27506, 
        n27505, n27504, n27503, n22880, n6352, n27502, n27501, 
        n27500, n27499, n27498;
    wire [7:0]state_7__N_4100;
    
    wire n45794, n27497, n27496, n27495, n27486, n27485, n27484, 
        n45793, n27483, n27482, n26769, n27470, n27469, n27468, 
        n27467, n27466, n27465, n45792, n45791, n45790, n45789, 
        n26768, n27464, n27463, n27462, n45788, n52303, n27461, 
        n27460, n27459, n25264, n52311, n52842, n22568, n26655, 
        n27458, n27457, n27456, n27455, n27454, n27453, n27452, 
        n51577, n23_adj_5810, n6_adj_5811, n11_adj_5812, n11_adj_5813, 
        n51579, n27439, n38306, n45787, n45786, n45785, n45784, 
        n35696, n68, n35706, n35720, n35727, n45783, n45782, n27433, 
        n78, n82, n52217, n45781, n22907, n45780, n41, n45779, 
        n45778, n45777, n45776, n45775, n45500, n45774, n25356, 
        n45773, n4_adj_5814, n45772, n45771, n59836, n45770, n45769, 
        n45768, n45767, n45766, n22875, n45765, n62688, n45764, 
        n10_adj_5815, n23688, n22896, n56196, n9_adj_5816, n45763, 
        n45762, n13_adj_5817, n25346, n62532, n56672, n23958, n23945, 
        n45761, n59809, n38302, n59807, n32_adj_5818, n27430, n45760, 
        n25081, n4_adj_5819, n6_adj_5820, n8_adj_5821, n9_adj_5822, 
        n11_adj_5823, n13_adj_5824, n14_adj_5825, n15_adj_5826, n4_adj_5827, 
        n6_adj_5828, n8_adj_5829, n9_adj_5830, n48, n49, n50, n51, 
        n52, n53, n54, n55, n45759, n45758, n25039, n45529, 
        n45528, n9582, n20140, n45757, n25021, n25014, n25013, 
        n52158, n52312, n45756, n60471, n52313, n52848, n26705, 
        n52318, n52317, n52316, n52315, n52314, n52304, n52219, 
        n60461, n61603, n60455, n62685, n52301, n52300, n52299, 
        n52298, n52297, n26402, n52296, n45755, n25768, n25766, 
        n25761, n52432, n52434, n25750, n52430, n52412, n25739, 
        n25734, n25713, n25709, n25707, n25705, n25699, n26176, 
        n24962, n26400, n52307, n52302, n52308, n26399, n45488, 
        n52295, n12_adj_5831, n52294, n52293, n52292, n52291, n52290, 
        n52306, n52289, n26391, n26390, n24938, n52053, n45754, 
        n45527, n490, n45526, n45525, n472, n399, n52305, n417, 
        n45753, n45524, n45752, n51575, n45751, n45750, n344_adj_5832, 
        n45499, n27391, n45498, n253_adj_5833, n45749, n271, n326, 
        n45523, n62430, n62427, n62418, n62415, n62403, n14_adj_5834, 
        n180, n45748, n198, n10_adj_5835, n125, n27387, n27379, 
        n27375, n27370, n27365, n38354, n35, n53_adj_5836, n107, 
        n52155, n51669, n27331, n27327, n22918, n22893, n45497, 
        n45522, n46065, n46064, n52288, n46063, n45747, n45746, 
        n23824, n45496, n45521, n45495, n46062, n45745, n45744, 
        n46061, n23338, n46060, n46059, n27321, n27317, n27312, 
        n23375, n45520, n26749, n26746, n52427, n26743, n26740, 
        n26737, n27259, n27257, n27256, n27255, n52159, n45743, 
        n45519, n45494, n45518, n22774, n45742, n45741, n26731, 
        n52287, n45487, n52286, n45517, n14_adj_5837, n13_adj_5838, 
        n52285, n26734, n52284, n45516, n45515, n45514, n45486, 
        n23594, n48661, n54861, n45513, n23531, n33996, n45512, 
        n60412, n52513, n5_adj_5839, n45511, n23427, n4_adj_5840, 
        n3_adj_5841, n45510, n55054, n22870, n56825, n22594, n47529, 
        n22765, n47509, n47989, n545, n47452, n6_adj_5842, n9_adj_5843, 
        n4_adj_5844, n47380, n61591, n10_adj_5845, n4_adj_5846, n60212, 
        n16_adj_5847, n62667, n60167, n60154, n60152, n4_adj_5848, 
        n62658, n60110, n56674, n56673, n60092, n60080, n56668, 
        n56667, n50845, n24_adj_5849, n56665, n17_adj_5850, n25_adj_5851, 
        n53300, n53298, n50941, n56463, n56664, n56475, n59386, 
        n59385, n55846, n54039, n54035, n55830, n52928, n52496, 
        n52584, n52564, n59364, n55814, n52741, n55011, n54720, 
        n51153, n55798, n52939, n52922, n53140, n53137, n52979, 
        n55782, n59353, n15_adj_5852, n29, n14_adj_5853, n53069, 
        n53055, n53035, n27, n23_adj_5854, n59349, n54886, n54882, 
        n55766, n54842, n59342, n59339, n55750, n59325, n55734, 
        n59312, n59311, n59310, n59309, n59308, n62103, n62102, 
        n59307, n59306, n56302, n62086, n62080, n53122, n53113, 
        n53098, n53092, n52362, n56826, n62021, n53161, n59565, 
        n53125, n59279, n62835, n52409, n61981, n52424, n62829, 
        n61935, n62823, n61699, n52435, n54312, n56306, n62817, 
        n61980, n61874, n51549, n59538, n62811, n51585, n62805, 
        n9_adj_5855, n62799, n62793, n8_adj_5856, n52641, n52925, 
        n51655, n51659, n51663, n51667, n51673, n51677, n51681, 
        n62787, n61784, n61783, n62401, n59198, n59196, n62781, 
        n59192, n52455, n51817, n62775, n6_adj_5857, n61604, n61592, 
        n62640, n62769, n52656, n24_adj_5858, n55156, n20_adj_5859, 
        n51973, n62763, n15_adj_5860, n14_adj_5861, n62757, n56589, 
        n56588, n62751, n62840, n6_adj_5862;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 i24349_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i24349_2_lut.LUT_INIT = 16'h8888;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_188 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_183));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_190 (.Q(dti), .C(clk16MHz), .E(n24938), .D(dti_N_380));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 add_156_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n45522), .O(n1269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[0]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4100[3])) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_43[0]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5702));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_156_18 (.CI(n45522), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n45523));
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .GND_net(GND_net), 
            .state({state}), .VCC_net(VCC_net), .n20312(n20312), .bit_ctr({Open_0, 
            Open_1, Open_2, bit_ctr[1:0]}), .n7(n7_adj_5718), .\neopxl_color[9] (neopxl_color[9]), 
            .\neopxl_color[8] (neopxl_color[8]), .\color_bit_N_478[1] (color_bit_N_478[1]), 
            .n27543(n27543), .n51153(n51153), .n25081(n25081), .\bit_ctr[3] (bit_ctr[3]), 
            .\bit_ctr[4] (bit_ctr[4]), .NEOPXL_c(NEOPXL_c), .\neopxl_color[16] (neopxl_color[16]), 
            .\neopxl_color[17] (neopxl_color[17]), .\neopxl_color[18] (neopxl_color[18]), 
            .\neopxl_color[19] (neopxl_color[19]), .\neopxl_color[22] (neopxl_color[22]), 
            .\neopxl_color[23] (neopxl_color[23]), .\neopxl_color[20] (neopxl_color[20]), 
            .\neopxl_color[21] (neopxl_color[21]), .LED_c(LED_c), .n38354(n38354), 
            .n47529(n47529), .n56665(n56665), .n56663(n56663), .n62592(n62592), 
            .n62640(n62640), .\neopxl_color[10] (neopxl_color[10]), .\neopxl_color[11] (neopxl_color[11]), 
            .n62472(n62472), .n47509(n47509)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 i13537_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n55830), 
            .I3(n27), .O(n27243));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13537_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5696));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13845_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n25734), .I3(GND_net), .O(n27551));   // verilog/coms.v(130[12] 305[6])
    defparam i13845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[19] [7]), .I1(n10_adj_5755), .I2(n25734), 
            .I3(n52362), .O(n51549));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1780 (.I0(\data_in_frame[19] [4]), .I1(n53298), 
            .I2(n25734), .I3(rx_data[4]), .O(n51567));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1780.LUT_INIT = 16'h3a0a;
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5701));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n55156));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i13399_3_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n25739), .I3(GND_net), .O(n27105));   // verilog/coms.v(130[12] 305[6])
    defparam i13399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5695));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13873_3_lut (.I0(n53350), .I1(r_Bit_Index[0]), .I2(n25264), 
            .I3(GND_net), .O(n27579));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13873_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5700));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1068_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3464[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5830));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1068_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n51973));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut.LUT_INIT = 16'hd054;
    SB_LUT4 i1_2_lut (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), .I1(Ki[1]), 
            .I2(GND_net), .I3(GND_net), .O(n107));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5694));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1068_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3464[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3464[0]), .O(n4_adj_5827));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1068_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mux_252_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_67[6]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_1068_i8_3_lut (.I0(n6_adj_5828), .I1(o_Rx_DV_N_3464[4]), 
            .I2(n9_adj_5830), .I3(GND_net), .O(n8_adj_5829));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1068_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5693));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i44773_3_lut (.I0(state_7__N_4084[0]), .I1(n37902), .I2(enable_slow_N_4187), 
            .I3(GND_net), .O(n59385));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i44773_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_5946[0]), .I1(n59385), .I2(n6352), 
            .I3(n6_adj_5721), .O(n8_adj_5856));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i13866_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[0]), 
            .I2(counter_adj_5947[0]), .I3(n22875), .O(n27572));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13866_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i20329_3_lut (.I0(n214), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(n33996));
    defparam i20329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24258_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i24258_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1781 (.I0(n33996), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_5836));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5692));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13247_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n52427), .I3(GND_net), .O(n26953));   // verilog/coms.v(130[12] 305[6])
    defparam i13247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47080_4_lut (.I0(n8_adj_5829), .I1(n4_adj_5827), .I2(n9_adj_5830), 
            .I3(n59538), .O(n61980));   // verilog/uart_rx.v(119[17:57])
    defparam i47080_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47081_3_lut (.I0(n61980), .I1(o_Rx_DV_N_3464[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n61981));   // verilog/uart_rx.v(119[17:57])
    defparam i47081_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13877_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n55782), 
            .I3(n27), .O(n27583));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13877_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13878_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[0]), .I2(n11_adj_5757), 
            .I3(state_7__N_4293), .O(n27584));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13878_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_252_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_67[7]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i46974_3_lut (.I0(n61981), .I1(o_Rx_DV_N_3464[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n61874));   // verilog/uart_rx.v(119[17:57])
    defparam i46974_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n25013), 
            .D(n1284), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n25013), 
            .D(n1283), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i46890_3_lut (.I0(n61874), .I1(o_Rx_DV_N_3464[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4855));   // verilog/uart_rx.v(119[17:57])
    defparam i46890_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n25013), 
            .D(n1282), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n25013), 
            .D(n1281), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n25013), 
            .D(n1280), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i1_2_lut_adj_1782 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[2]), .I2(GND_net), .I3(GND_net), .O(n180));
    defparam i1_2_lut_adj_1782.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n25013), 
            .D(n1279), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n25013), 
            .D(n1278), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n25013), 
            .D(n1277), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n25013), 
            .D(n1276), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i1_2_lut_adj_1783 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[3]), .I2(GND_net), .I3(GND_net), .O(n253_adj_5833));
    defparam i1_2_lut_adj_1783.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n25013), 
            .D(n1275), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i13546_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[2]), 
            .I2(counter_adj_5947[0]), .I3(n22918), .O(n27252));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13546_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47724 (.I0(byte_transmit_counter[3]), 
            .I1(n61003), .I2(n59386), .I3(byte_transmit_counter[4]), .O(n62667));
    defparam byte_transmit_counter_3__bdd_4_lut_47724.LUT_INIT = 16'he4aa;
    SB_LUT4 n62667_bdd_4_lut (.I0(n62667), .I1(n41), .I2(n52053), .I3(byte_transmit_counter[4]), 
            .O(tx_data[2]));
    defparam n62667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n25013), 
            .D(n1274), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n25013), 
            .D(n1273), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i1_2_lut_adj_1784 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[4]), .I2(GND_net), .I3(GND_net), .O(n326));
    defparam i1_2_lut_adj_1784.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1785 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[5]), .I2(GND_net), .I3(GND_net), .O(n399));
    defparam i1_2_lut_adj_1785.LUT_INIT = 16'h8888;
    SB_LUT4 i13539_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n55798), 
            .I3(n27), .O(n27245));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13539_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i591_2_lut (.I0(n1365), .I1(n37857), .I2(GND_net), .I3(GND_net), 
            .O(n2925));   // verilog/TinyFPGA_B.v(386[18] 388[12])
    defparam i591_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_252_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_67[8]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_252_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_67[9]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1786 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[6]), .I2(GND_net), .I3(GND_net), .O(n472));
    defparam i1_2_lut_adj_1786.LUT_INIT = 16'h8888;
    SB_LUT4 i22037_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[10]));
    defparam i22037_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_67[10]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_252_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_67[11]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i44958_4_lut (.I0(data_ready), .I1(n6543), .I2(n24_adj_5849), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n59339));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i44958_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i45303_2_lut (.I0(n24_adj_5849), .I1(n6543), .I2(GND_net), 
            .I3(GND_net), .O(n59342));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i45303_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13540_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n55750), 
            .I3(n27), .O(n27246));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13540_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49_4_lut (.I0(n59342), .I1(n59339), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5723), .O(n50845));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 add_237_5_lut (.I0(current[3]), .I1(duty[6]), .I2(n62401), 
            .I3(n45488), .O(n267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_237_13_lut (.I0(current[11]), .I1(duty[14]), .I2(n62401), 
            .I3(n45496), .O(n259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_1787 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[7]), .I2(GND_net), .I3(GND_net), .O(n545));
    defparam i1_2_lut_adj_1787.LUT_INIT = 16'h8888;
    SB_LUT4 i13884_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n52435), 
            .I3(GND_net), .O(n27590));   // verilog/coms.v(130[12] 305[6])
    defparam i13884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_156_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n45521), .O(n1270)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_17 (.CI(n45521), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n45522));
    SB_LUT4 add_156_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n45520), .O(n1271)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5691));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13541_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n55766), 
            .I3(n27), .O(n27247));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13541_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n25013), 
            .D(n1272), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n25013), 
            .D(n1271), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_156_16 (.CI(n45520), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n45521));
    SB_LUT4 LessThan_1068_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3464[3]), 
            .I2(o_Rx_DV_N_3464[2]), .I3(GND_net), .O(n6_adj_5828));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1068_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n25013), 
            .D(n1270), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[23]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[22]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[21]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 add_156_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n45519), .O(n1272)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_13 (.CI(n45496), .I0(duty[14]), .I1(n62401), .CO(n45497));
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_CARRY add_156_15 (.CI(n45519), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n45520));
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 add_237_12_lut (.I0(current[10]), .I1(duty[13]), .I2(n62401), 
            .I3(n45495), .O(n260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_12_lut.LUT_INIT = 16'hA3AC;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_CARRY add_237_5 (.CI(n45488), .I0(duty[6]), .I1(n62401), .CO(n45489));
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n25013), 
            .D(n1269), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 add_156_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n45518), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_14 (.CI(n45518), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n45519));
    SB_CARRY add_237_12 (.CI(n45495), .I0(duty[13]), .I1(n62401), .CO(n45496));
    SB_LUT4 add_156_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n45517), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_13 (.CI(n45517), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n45518));
    SB_LUT4 add_156_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n45516), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_12 (.CI(n45516), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n45517));
    SB_LUT4 add_237_11_lut (.I0(current[9]), .I1(duty[12]), .I2(n62401), 
            .I3(n45494), .O(n261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_11_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i20034_3_lut (.I0(n220), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691 [11]));
    defparam i20034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_252_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_67[12]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_237_4_lut (.I0(current[2]), .I1(duty[5]), .I2(n62401), 
            .I3(n45487), .O(n268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_156_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n45515), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_11 (.CI(n45515), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n45516));
    SB_LUT4 add_156_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n45514), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_11 (.CI(n45494), .I0(duty[12]), .I1(n62401), .CO(n45495));
    SB_CARRY add_156_10 (.CI(n45514), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n45515));
    SB_LUT4 add_156_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n45513), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_9 (.CI(n45513), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n45514));
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n25013), 
            .D(n1268), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 n62715_bdd_4_lut (.I0(n62715), .I1(duty[2]), .I2(n268), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n62715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i44638_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3464[3]), 
            .I2(o_Rx_DV_N_3464[2]), .I3(r_Clock_Count[2]), .O(n59538));   // verilog/uart_rx.v(119[17:57])
    defparam i44638_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_adj_1788 (.I0(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I1(Ki[0]), .I2(GND_net), .I3(GND_net), .O(n35));
    defparam i1_2_lut_adj_1788.LUT_INIT = 16'h8888;
    SB_LUT4 add_156_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n45512), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_4 (.CI(n45487), .I0(duty[5]), .I1(n62401), .CO(n45488));
    SB_LUT4 add_237_10_lut (.I0(current[8]), .I1(duty[11]), .I2(n62401), 
            .I3(n45493), .O(n262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_10_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_156_8 (.CI(n45512), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n45513));
    SB_LUT4 LessThan_17_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5688));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5689));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5685));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5686));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5732));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_156_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n45511), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n25013), 
            .D(n1267), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 LessThan_17_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5730));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5690));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_156_19 (.CI(n45523), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n45524));
    SB_LUT4 LessThan_17_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5734));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45210_4_lut (.I0(n11_adj_5690), .I1(n9_adj_5730), .I2(n7_adj_5732), 
            .I3(n5_adj_5734), .O(n60110));
    defparam i45210_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_156_7 (.CI(n45511), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n45512));
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5731), .I1(current_limit[9]), 
            .I2(n19_adj_5685), .I3(GND_net), .O(n16_adj_5687));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5735));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n25013), 
            .D(n1266), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i46701_3_lut (.I0(n4_adj_5735), .I1(current_limit[5]), .I2(n11_adj_5690), 
            .I3(GND_net), .O(n61601));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i46701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46702_3_lut (.I0(n61601), .I1(current_limit[6]), .I2(n13_adj_5689), 
            .I3(GND_net), .O(n61602));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i46702_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n25013), 
            .D(n1265), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 add_156_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n45510), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45192_4_lut (.I0(n17_adj_5686), .I1(n15_adj_5688), .I2(n13_adj_5689), 
            .I3(n60110), .O(n60092));
    defparam i45192_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46987_4_lut (.I0(n16_adj_5687), .I1(n6_adj_5733), .I2(n19_adj_5685), 
            .I3(n60080), .O(n61887));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i46987_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45561_3_lut (.I0(n61602), .I1(current_limit[7]), .I2(n15_adj_5688), 
            .I3(GND_net), .O(n60461));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i45561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47179_4_lut (.I0(n60461), .I1(n61887), .I2(n19_adj_5685), 
            .I3(n60092), .O(n62079));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i47179_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47180_3_lut (.I0(n62079), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n62080));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i47180_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5835));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(dti_counter[7]), .I1(dti_counter[4]), .I2(dti_counter[5]), 
            .I3(dti_counter[6]), .O(n14_adj_5834));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5834), .I2(n10_adj_5835), 
            .I3(dti_counter[3]), .O(n20251));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5846));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'h7bde;
    SB_LUT4 i47119_3_lut (.I0(n62080), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i47119_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47419_2_lut (.I0(n20251), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_380));
    defparam i47419_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 LessThan_1071_i9_2_lut (.I0(r_Clock_Count_adj_5934[4]), .I1(o_Rx_DV_N_3464[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5822));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1071_i13_2_lut (.I0(r_Clock_Count_adj_5934[6]), .I1(o_Rx_DV_N_3464[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5824));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1071_i11_2_lut (.I0(r_Clock_Count_adj_5934[5]), .I1(o_Rx_DV_N_3464[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5823));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n54882));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n54886));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n54886), .I3(n54882), .O(n296));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1061_1_lut (.I0(n296), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n4847));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1061_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n25013), 
            .D(n1264), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_CARRY add_237_10 (.CI(n45493), .I0(duty[11]), .I1(n62401), .CO(n45494));
    SB_CARRY add_156_6 (.CI(n45510), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n45511));
    SB_LUT4 add_156_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n45509), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_5 (.CI(n45509), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n45510));
    SB_LUT4 add_156_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n45508), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_4 (.CI(n45508), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n45509));
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n25013), 
            .D(n1263), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_183), 
            .I3(n45561), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_237_9_lut (.I0(current[7]), .I1(duty[10]), .I2(n62401), 
            .I3(n45492), .O(n263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n4847), .I1(GND_net), .I2(pwm_setpoint_23__N_183), 
            .I3(n45560), .O(n5012)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n45560), .I0(GND_net), .I1(pwm_setpoint_23__N_183), 
            .CO(n45561));
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(n4847), .I1(GND_net), .I2(n3), 
            .I3(n45559), .O(n5013)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_24 (.CI(n45559), .I0(GND_net), .I1(n3), 
            .CO(n45560));
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(n4847), .I1(GND_net), .I2(n4_adj_5691), 
            .I3(n45558), .O(n5014)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n45558), .I0(GND_net), .I1(n4_adj_5691), 
            .CO(n45559));
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [2]), 
            .O(n52243));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(n4847), .I1(GND_net), .I2(n5_adj_5692), 
            .I3(n45557), .O(n5015)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [3]), 
            .O(n52242));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1793.LUT_INIT = 16'h2300;
    SB_LUT4 i13931_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n52432), .I3(GND_net), .O(n27637));   // verilog/coms.v(130[12] 305[6])
    defparam i13931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1794 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [4]), 
            .O(n52241));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1794.LUT_INIT = 16'h2300;
    SB_LUT4 i13269_3_lut_4_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26975));   // verilog/coms.v(130[12] 305[6])
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n45557), .I0(GND_net), .I1(n5_adj_5692), 
            .CO(n45558));
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(n4847), .I1(GND_net), .I2(n6_adj_5693), 
            .I3(n45556), .O(n5016)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_21 (.CI(n45556), .I0(GND_net), .I1(n6_adj_5693), 
            .CO(n45557));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1795 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [5]), 
            .O(n52240));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1795.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1796 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [6]), 
            .O(n52239));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1796.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1797 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [7]), 
            .O(n52223));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1797.LUT_INIT = 16'h2300;
    SB_LUT4 i13262_3_lut_4_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26968));   // verilog/coms.v(130[12] 305[6])
    defparam i13262_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(control_mode[3]), .I1(control_mode[6]), 
            .I2(control_mode[2]), .I3(control_mode[4]), .O(n56196));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n56196), .I1(control_mode[7]), .I2(control_mode[5]), 
            .I3(GND_net), .O(n22887));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1799 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [0]), 
            .O(n52238));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1799.LUT_INIT = 16'h2300;
    SB_LUT4 n62637_bdd_4_lut (.I0(n62637), .I1(neopxl_color[6]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[0]), .O(n62640));
    defparam n62637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1800 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [1]), 
            .O(n52237));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1800.LUT_INIT = 16'h2300;
    SB_LUT4 i13250_3_lut_4_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26956));   // verilog/coms.v(130[12] 305[6])
    defparam i13250_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1801 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [2]), 
            .O(n52236));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1801.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1802 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [3]), 
            .O(n52235));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1802.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_adj_1803 (.I0(control_mode[0]), .I1(n22887), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5724));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_1803.LUT_INIT = 16'hfdfd;
    SB_LUT4 i13240_3_lut_4_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26946));   // verilog/coms.v(130[12] 305[6])
    defparam i13240_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_252_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_67[18]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(n4847), .I1(GND_net), .I2(n7_adj_5694), 
            .I3(n45555), .O(n5017)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_237_3_lut (.I0(current[1]), .I1(duty[4]), .I2(n62401), 
            .I3(n45486), .O(n269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_156_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n45507), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13238_3_lut_4_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26944));   // verilog/coms.v(130[12] 305[6])
    defparam i13238_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13_4_lut_adj_1804 (.I0(\data_in_frame[19] [3]), .I1(n53298), 
            .I2(n25734), .I3(rx_data[3]), .O(n51575));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1804.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1805 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [4]), 
            .O(n52234));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1805.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_21_add_3_20 (.CI(n45555), .I0(GND_net), .I1(n7_adj_5694), 
            .CO(n45556));
    SB_LUT4 i13_4_lut_adj_1806 (.I0(\data_in_frame[19] [2]), .I1(n53298), 
            .I2(n25734), .I3(rx_data[2]), .O(n51577));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1806.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13372_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n20140), .I3(GND_net), .O(n27078));   // verilog/coms.v(130[12] 305[6])
    defparam i13372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13237_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5933[1]), 
            .I2(r_SM_Main_adj_5933[2]), .I3(n6_adj_5842), .O(n26943));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13237_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i13373_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n20140), .I3(GND_net), .O(n27079));   // verilog/coms.v(130[12] 305[6])
    defparam i13373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13395_3_lut (.I0(\data_in_frame[16] [0]), .I1(rx_data[0]), 
            .I2(n25739), .I3(GND_net), .O(n27101));   // verilog/coms.v(130[12] 305[6])
    defparam i13395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1807 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [5]), 
            .O(n52233));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1807.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(n4847), .I1(GND_net), .I2(n8_adj_5695), 
            .I3(n45554), .O(n5018)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'h8228;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1808 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [6]), 
            .O(n52232));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1808.LUT_INIT = 16'h2300;
    SB_LUT4 i13938_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n52432), .I3(GND_net), .O(n27644));   // verilog/coms.v(130[12] 305[6])
    defparam i13938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_252_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i1_3_lut (.I0(encoder0_position_scaled[0]), .I1(motor_state_23__N_67[0]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i1_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n45554), .I0(GND_net), .I1(n8_adj_5695), 
            .CO(n45555));
    SB_LUT4 i13941_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n52432), .I3(GND_net), .O(n27647));   // verilog/coms.v(130[12] 305[6])
    defparam i13941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(n4847), .I1(GND_net), .I2(n9_adj_5696), 
            .I3(n45553), .O(n5019)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13944_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n52432), .I3(GND_net), .O(n27650));   // verilog/coms.v(130[12] 305[6])
    defparam i13944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[16] [7]), 
            .O(n52231));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [0]), 
            .O(n26327));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1811 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [1]), 
            .O(n52230));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1811.LUT_INIT = 16'h2300;
    SB_LUT4 mux_250_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_67[1]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13224_3_lut_4_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26930));   // verilog/coms.v(130[12] 305[6])
    defparam i13224_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY unary_minus_21_add_3_18 (.CI(n45553), .I0(GND_net), .I1(n9_adj_5696), 
            .CO(n45554));
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(n4847), .I1(GND_net), .I2(n10_adj_5697), 
            .I3(n45552), .O(n5020)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13947_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n52432), .I3(GND_net), .O(n27653));   // verilog/coms.v(130[12] 305[6])
    defparam i13947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_252_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_67[2]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13950_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n52432), .I3(GND_net), .O(n27656));   // verilog/coms.v(130[12] 305[6])
    defparam i13950_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n45552), .I0(GND_net), .I1(n10_adj_5697), 
            .CO(n45553));
    SB_LUT4 i13374_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n20140), .I3(GND_net), .O(n27080));   // verilog/coms.v(130[12] 305[6])
    defparam i13374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13223_3_lut_4_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26929));   // verilog/coms.v(130[12] 305[6])
    defparam i13223_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13219_3_lut_4_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26925));   // verilog/coms.v(130[12] 305[6])
    defparam i13219_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1812 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [2]), 
            .O(n52229));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1812.LUT_INIT = 16'h2300;
    SB_LUT4 i13218_3_lut_4_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26924));   // verilog/coms.v(130[12] 305[6])
    defparam i13218_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n25013), 
            .D(n1262), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i13375_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n20140), .I3(GND_net), .O(n27081));   // verilog/coms.v(130[12] 305[6])
    defparam i13375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13376_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n20140), .I3(GND_net), .O(n27082));   // verilog/coms.v(130[12] 305[6])
    defparam i13376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [3]), 
            .O(n52228));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 i13214_3_lut_4_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26920));   // verilog/coms.v(130[12] 305[6])
    defparam i13214_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(n4847), .I1(GND_net), .I2(n11_adj_5698), 
            .I3(n45551), .O(n5021)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1090_25_lut (.I0(GND_net), .I1(n5010), .I2(n5034), .I3(n45799), 
            .O(n418)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13377_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n20140), .I3(GND_net), .O(n27083));   // verilog/coms.v(130[12] 305[6])
    defparam i13377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13378_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n20140), .I3(GND_net), .O(n27084));   // verilog/coms.v(130[12] 305[6])
    defparam i13378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13379_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n20140), .I3(GND_net), .O(n27085));   // verilog/coms.v(130[12] 305[6])
    defparam i13379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1071_i15_2_lut (.I0(r_Clock_Count_adj_5934[7]), .I1(o_Rx_DV_N_3464[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5826));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i21460_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n20140), .I3(GND_net), .O(n27086));
    defparam i21460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21462_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n20140), .I3(GND_net), .O(n27087));
    defparam i21462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13382_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n20140), .I3(GND_net), .O(n27088));   // verilog/coms.v(130[12] 305[6])
    defparam i13382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13210_3_lut_4_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26916));   // verilog/coms.v(130[12] 305[6])
    defparam i13210_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13383_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n20140), .I3(GND_net), .O(n27089));   // verilog/coms.v(130[12] 305[6])
    defparam i13383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13384_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n20140), .I3(GND_net), .O(n27090));   // verilog/coms.v(130[12] 305[6])
    defparam i13384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1090_24_lut (.I0(GND_net), .I1(n5010), .I2(n5035), .I3(n45798), 
            .O(n419)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n25013), 
            .D(n1261), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_CARRY unary_minus_21_add_3_16 (.CI(n45551), .I0(GND_net), .I1(n11_adj_5698), 
            .CO(n45552));
    SB_LUT4 i13953_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n52432), .I3(GND_net), .O(n27659));   // verilog/coms.v(130[12] 305[6])
    defparam i13953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_252_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_67[3]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13209_3_lut_4_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26915));   // verilog/coms.v(130[12] 305[6])
    defparam i13209_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13956_3_lut (.I0(\data_in_frame[20] [7]), .I1(rx_data[7]), 
            .I2(n52432), .I3(GND_net), .O(n27662));   // verilog/coms.v(130[12] 305[6])
    defparam i13956_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [4]), 
            .O(n52227));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [5]), 
            .O(n52226));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1816 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [6]), 
            .O(n52225));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1816.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1817 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [7]), 
            .O(n52155));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1817.LUT_INIT = 16'h2300;
    SB_LUT4 mux_250_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_67[4]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1818 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [0]), 
            .O(n26319));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1818.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1819 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [1]), 
            .O(n52220));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1819.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1820 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [2]), 
            .O(n26317));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1820.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_1071_i4_4_lut (.I0(r_Clock_Count_adj_5934[0]), .I1(o_Rx_DV_N_3464[1]), 
            .I2(r_Clock_Count_adj_5934[1]), .I3(o_Rx_DV_N_3464[0]), .O(n4_adj_5819));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_156_3 (.CI(n45507), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n45508));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [3]), 
            .O(n52221));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 mux_250_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_67[5]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [4]), 
            .O(n52222));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h2300;
    SB_LUT4 i13385_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n20140), .I3(GND_net), .O(n27091));   // verilog/coms.v(130[12] 305[6])
    defparam i13385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24553_2_lut_2_lut (.I0(duty[14]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5043));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24553_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13386_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n20140), .I3(GND_net), .O(n27092));   // verilog/coms.v(130[12] 305[6])
    defparam i13386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13387_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n20140), .I3(GND_net), .O(n27093));   // verilog/coms.v(130[12] 305[6])
    defparam i13387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13388_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n20140), .I3(GND_net), .O(n27094));   // verilog/coms.v(130[12] 305[6])
    defparam i13388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13389_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n20140), .I3(GND_net), .O(n27095));   // verilog/coms.v(130[12] 305[6])
    defparam i13389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [5]), 
            .O(n52224));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h2300;
    SB_LUT4 i46883_3_lut (.I0(n4_adj_5819), .I1(o_Rx_DV_N_3464[5]), .I2(n11_adj_5823), 
            .I3(GND_net), .O(n61783));   // verilog/uart_tx.v(117[17:57])
    defparam i46883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [6]), 
            .O(n52159));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [7]), 
            .O(n52219));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h2300;
    SB_CARRY add_1090_24 (.CI(n45798), .I0(n5010), .I1(n5035), .CO(n45799));
    SB_LUT4 add_1090_23_lut (.I0(GND_net), .I1(n5010), .I2(n5036), .I3(n45797), 
            .O(n420)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [0]), 
            .O(n52161));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [1]), 
            .O(n52162));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h2300;
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n25013), 
            .D(n1260), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [2]), 
            .O(n52163));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(n4847), .I1(GND_net), .I2(n12), 
            .I3(n45550), .O(n5022)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n45550), .I0(GND_net), .I1(n12), 
            .CO(n45551));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(n4847), .I1(GND_net), .I2(n13_adj_5699), 
            .I3(n45549), .O(n5023)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [3]), 
            .O(n52164));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [4]), 
            .O(n52165));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_21_add_3_14 (.CI(n45549), .I0(GND_net), .I1(n13_adj_5699), 
            .CO(n45550));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(n4847), .I1(GND_net), .I2(n14), 
            .I3(n45548), .O(n5024)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13843_3_lut_4_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27549));   // verilog/coms.v(130[12] 305[6])
    defparam i13843_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_1090_23 (.CI(n45797), .I0(n5010), .I1(n5036), .CO(n45798));
    SB_LUT4 i46884_3_lut (.I0(n61783), .I1(o_Rx_DV_N_3464[6]), .I2(n13_adj_5824), 
            .I3(GND_net), .O(n61784));   // verilog/uart_tx.v(117[17:57])
    defparam i46884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45512_4_lut (.I0(n13_adj_5824), .I1(n11_adj_5823), .I2(n9_adj_5822), 
            .I3(n59565), .O(n60412));
    defparam i45512_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_1090_22_lut (.I0(GND_net), .I1(n5012), .I2(n5037), .I3(n45796), 
            .O(n421)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [5]), 
            .O(n52166));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 i13837_4_lut_4_lut (.I0(n25081), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n27543));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13837_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i21013_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n20140), .I3(GND_net), .O(n27096));
    defparam i21013_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1090_22 (.CI(n45796), .I0(n5012), .I1(n5037), .CO(n45797));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_43[23]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_43[22]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 i20987_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n20140), .I3(GND_net), .O(n27097));
    defparam i20987_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_43[21]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_43[20]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_43[19]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 add_1090_21_lut (.I0(GND_net), .I1(n5013), .I2(n5038), .I3(n45795), 
            .O(n422)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_1071_i8_3_lut (.I0(n6_adj_5820), .I1(o_Rx_DV_N_3464[4]), 
            .I2(n9_adj_5822), .I3(GND_net), .O(n8_adj_5821));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_43[18]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_43[17]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_43[16]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_43[15]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_43[14]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_43[13]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_43[12]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_43[11]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_43[10]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_43[9]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_43[8]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_43[7]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_43[6]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_43[5]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_43[4]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_43[3]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [6]), 
            .O(n52167));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h2300;
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_43[2]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_43[1]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n25013), 
            .D(n1259), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 i13393_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n20140), .I3(GND_net), .O(n27099));   // verilog/coms.v(130[12] 305[6])
    defparam i13393_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[1]));   // verilog/TinyFPGA_B.v(320[10] 327[6])
    SB_LUT4 i46589_3_lut (.I0(n61784), .I1(o_Rx_DV_N_3464[7]), .I2(n15_adj_5826), 
            .I3(GND_net), .O(n14_adj_5825));   // verilog/uart_tx.v(117[17:57])
    defparam i46589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20896_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n20140), .I3(GND_net), .O(n27100));
    defparam i20896_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n25013), 
            .D(n1258), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n50845));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 i46289_4_lut (.I0(n14_adj_5825), .I1(n8_adj_5821), .I2(n15_adj_5826), 
            .I3(n60412), .O(n61189));   // verilog/uart_tx.v(117[17:57])
    defparam i46289_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[19] [7]), 
            .O(n52168));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h2300;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n51973));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_1090_21 (.CI(n45795), .I0(n5013), .I1(n5038), .CO(n45796));
    SB_CARRY unary_minus_21_add_3_13 (.CI(n45548), .I0(GND_net), .I1(n14), 
            .CO(n45549));
    SB_LUT4 add_1090_20_lut (.I0(GND_net), .I1(n5014), .I2(n5039), .I3(n45794), 
            .O(n423)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_20 (.CI(n45794), .I0(n5014), .I1(n5039), .CO(n45795));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(n4847), .I1(GND_net), .I2(n15_adj_5700), 
            .I3(n45547), .O(n5025)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1090_19_lut (.I0(GND_net), .I1(n5015), .I2(n5040), .I3(n45793), 
            .O(n424)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_19 (.CI(n45793), .I0(n5015), .I1(n5040), .CO(n45794));
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n25013), 
            .D(n1257), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 add_1090_18_lut (.I0(GND_net), .I1(n5016), .I2(n5041), .I3(n45792), 
            .O(n425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n45547), .I0(GND_net), .I1(n15_adj_5700), 
            .CO(n45548));
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(bit_ctr[3]), .I2(n38354), 
            .I3(bit_ctr[4]), .O(n4_adj_5814));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hd555;
    SB_DFF read_202 (.Q(state_7__N_3892[0]), .C(clk16MHz), .D(n55156));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n25013), 
            .D(n1256), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_237_9 (.CI(n45492), .I0(duty[10]), .I1(n62401), .CO(n45493));
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n25013), 
            .D(n1255), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n25013), 
            .D(n1254), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i24554_2_lut_2_lut (.I0(duty[13]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5044));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24554_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY add_1090_18 (.CI(n45792), .I0(n5016), .I1(n5041), .CO(n45793));
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(n4847), .I1(GND_net), .I2(n16_adj_5701), 
            .I3(n45546), .O(n5026)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'h8228;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF dti_counter_1928__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [0]), 
            .O(n52169));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h2300;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i46290_3_lut (.I0(n61189), .I1(o_Rx_DV_N_3464[8]), .I2(r_Clock_Count_adj_5934[8]), 
            .I3(GND_net), .O(n4858));   // verilog/uart_tx.v(117[17:57])
    defparam i46290_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n45546), .I0(GND_net), .I1(n16_adj_5701), 
            .CO(n45547));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [1]), 
            .O(n26302));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_LUT4 add_1090_17_lut (.I0(GND_net), .I1(n5017), .I2(n5042), .I3(n45791), 
            .O(n426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_17 (.CI(n45791), .I0(n5017), .I1(n5042), .CO(n45792));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47669 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n62595));
    defparam byte_transmit_counter_0__bdd_4_lut_47669.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main_adj_5933[0]), .I1(o_Rx_DV_N_3464[24]), 
            .I2(n27), .I3(GND_net), .O(n14_adj_5861));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 n62595_bdd_4_lut (.I0(n62595), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n62598));
    defparam n62595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1836 (.I0(n29), .I1(o_Rx_DV_N_3464[12]), .I2(n23_adj_5854), 
            .I3(n4858), .O(n15_adj_5860));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut_adj_1836.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5860), .I1(r_SM_Main_adj_5933[2]), .I2(n14_adj_5861), 
            .I3(r_SM_Main_adj_5933[1]), .O(n62840));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(n4847), .I1(GND_net), .I2(n17_adj_5702), 
            .I3(n45545), .O(n5027)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n45545), .I0(GND_net), .I1(n17_adj_5702), 
            .CO(n45546));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1837 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [2]), 
            .O(n52170));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1837.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1838 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [3]), 
            .O(n26300));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1838.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1839 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [4]), 
            .O(n52171));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1839.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [5]), 
            .O(n52172));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n51937));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_1090_16_lut (.I0(GND_net), .I1(n5018), .I2(n5043), .I3(n45790), 
            .O(n427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_16 (.CI(n45790), .I0(n5018), .I1(n5043), .CO(n45791));
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5850));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_LUT4 add_1090_15_lut (.I0(GND_net), .I1(n5019), .I2(n5044), .I3(n45789), 
            .O(n428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_15 (.CI(n45789), .I0(n5019), .I1(n5044), .CO(n45790));
    SB_LUT4 add_1090_14_lut (.I0(GND_net), .I1(n5020), .I2(n5045), .I3(n45788), 
            .O(n429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_14 (.CI(n45788), .I0(n5020), .I1(n5045), .CO(n45789));
    SB_LUT4 n62589_bdd_4_lut (.I0(n62589), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(color_bit_N_478[1]), .O(n62592));
    defparam n62589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_1090_13_lut (.I0(GND_net), .I1(n5021), .I2(n5046), .I3(n45787), 
            .O(n430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_13 (.CI(n45787), .I0(n5021), .I1(n5046), .CO(n45788));
    SB_LUT4 add_1090_12_lut (.I0(GND_net), .I1(n5022), .I2(n5047), .I3(n45786), 
            .O(n431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(n4847), .I1(GND_net), .I2(n18), 
            .I3(n45544), .O(n5028)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [6]), 
            .O(n52173));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n45544), .I0(GND_net), .I1(n18), 
            .CO(n45545));
    SB_LUT4 add_156_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(n4847), .I1(GND_net), .I2(n19_adj_5703), 
            .I3(n45543), .O(n5029)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1090_12 (.CI(n45786), .I0(n5022), .I1(n5047), .CO(n45787));
    SB_LUT4 add_1090_11_lut (.I0(GND_net), .I1(n5023), .I2(n5048), .I3(n45785), 
            .O(n432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_11 (.CI(n45785), .I0(n5023), .I1(n5048), .CO(n45786));
    SB_LUT4 i13733_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n25734), .I3(GND_net), .O(n27439));   // verilog/coms.v(130[12] 305[6])
    defparam i13733_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n45543), .I0(GND_net), .I1(n19_adj_5703), 
            .CO(n45544));
    SB_LUT4 add_1090_10_lut (.I0(GND_net), .I1(n5024), .I2(n5049), .I3(n45784), 
            .O(n433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_10 (.CI(n45784), .I0(n5024), .I1(n5049), .CO(n45785));
    SB_LUT4 add_1090_9_lut (.I0(GND_net), .I1(n5025), .I2(n5050), .I3(n45783), 
            .O(n434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_9 (.CI(n45783), .I0(n5025), .I1(n5050), .CO(n45784));
    SB_LUT4 add_1090_8_lut (.I0(GND_net), .I1(n5026), .I2(n5051), .I3(n45782), 
            .O(n435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47640 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[12] [2]), .I2(\data_out_frame[13] [2]), 
            .I3(byte_transmit_counter[2]), .O(n62565));
    defparam byte_transmit_counter_0__bdd_4_lut_47640.LUT_INIT = 16'he4aa;
    SB_LUT4 n62565_bdd_4_lut (.I0(n62565), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[2]), 
            .O(n62568));
    defparam n62565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_1090_8 (.CI(n45782), .I0(n5026), .I1(n5051), .CO(n45783));
    SB_LUT4 i13_4_lut_adj_1842 (.I0(\data_in_frame[19] [0]), .I1(n53298), 
            .I2(n25734), .I3(rx_data[0]), .O(n51579));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1842.LUT_INIT = 16'h3a0a;
    SB_LUT4 add_1090_7_lut (.I0(GND_net), .I1(n5027), .I2(n5052), .I3(n45781), 
            .O(n436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(n4847), .I1(GND_net), .I2(n20), 
            .I3(n45542), .O(n5030)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13545_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[1]), 
            .I2(counter_adj_5947[0]), .I3(n22875), .O(n27251));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13545_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY add_237_3 (.CI(n45486), .I0(duty[4]), .I1(n62401), .CO(n45487));
    SB_LUT4 i644_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2978));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i644_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13727_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n52435), 
            .I3(GND_net), .O(n27433));   // verilog/coms.v(130[12] 305[6])
    defparam i13727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13724_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n54720), .I3(GND_net), .O(n27430));   // verilog/coms.v(130[12] 305[6])
    defparam i13724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [7]), 
            .O(n52174));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 i13685_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n54720), .I3(GND_net), .O(n27391));   // verilog/coms.v(130[12] 305[6])
    defparam i13685_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [0]), 
            .O(n52175));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_LUT4 i13681_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n52435), 
            .I3(GND_net), .O(n27387));   // verilog/coms.v(130[12] 305[6])
    defparam i13681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_2_lut (.I0(IntegralLimit[11]), .I1(n143), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5810));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24555_2_lut_2_lut (.I0(duty[12]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5045));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24555_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13673_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n52435), 
            .I3(GND_net), .O(n27379));   // verilog/coms.v(130[12] 305[6])
    defparam i13673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1845 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [1]), 
            .O(n26294));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1845.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [2]), 
            .O(n52176));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [3]), 
            .O(n26292));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [4]), 
            .O(n52177));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 i13669_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n52435), 
            .I3(GND_net), .O(n27375));   // verilog/coms.v(130[12] 305[6])
    defparam i13669_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [5]), 
            .O(n52178));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_CARRY add_1090_7 (.CI(n45781), .I0(n5027), .I1(n5052), .CO(n45782));
    SB_LUT4 add_1090_6_lut (.I0(GND_net), .I1(n5028), .I2(n5053), .I3(n45780), 
            .O(n437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13664_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n52435), 
            .I3(GND_net), .O(n27370));   // verilog/coms.v(130[12] 305[6])
    defparam i13664_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13659_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n52435), 
            .I3(GND_net), .O(n27365));   // verilog/coms.v(130[12] 305[6])
    defparam i13659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[3] [7]), .I1(n25709), .I2(n25766), 
            .I3(rx_data[7]), .O(n51655));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_CARRY add_1090_6 (.CI(n45780), .I0(n5028), .I1(n5053), .CO(n45781));
    SB_LUT4 add_1090_5_lut (.I0(GND_net), .I1(n5029), .I2(n5054), .I3(n45779), 
            .O(n438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1090_5 (.CI(n45779), .I0(n5029), .I1(n5054), .CO(n45780));
    SB_LUT4 add_1090_4_lut (.I0(GND_net), .I1(n5030), .I2(n5055), .I3(n45778), 
            .O(n439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n25013), 
            .D(n1285), .R(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_DFFESR GHC_197 (.Q(GHC), .C(clk16MHz), .E(n24962), .D(GHC_N_367), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i24556_2_lut_2_lut (.I0(duty[11]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5046));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24556_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESR GHB_195 (.Q(GHB), .C(clk16MHz), .E(n24962), .D(GHB_N_353), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_193 (.Q(GHA), .C(clk16MHz), .E(n24962), .D(GHA_N_331), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5862), .D(commutation_state_7__N_184[0]), .S(commutation_state_7__N_192));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_194 (.Q(INLA_c_0), .C(clk16MHz), .E(n24962), .D(GLA_N_348), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLB_196 (.Q(INLB_c_0), .C(clk16MHz), .E(n24962), .D(GLB_N_362), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1850 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [6]), 
            .O(n52179));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1850.LUT_INIT = 16'h2300;
    SB_DFFESR GLC_198 (.Q(INLC_c_0), .C(clk16MHz), .E(n24962), .D(GLC_N_376), 
            .R(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dti_counter_1928__i1 (.Q(dti_counter[1]), .C(clk16MHz), .D(n54));   // verilog/TinyFPGA_B.v(174[23:37])
    GND i1 (.Y(GND_net));
    SB_DFF reset_203 (.Q(reset), .C(clk16MHz), .D(n50941));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    SB_CARRY add_1090_4 (.CI(n45778), .I0(n5030), .I1(n5055), .CO(n45779));
    SB_DFF dti_counter_1928__i2 (.Q(dti_counter[2]), .C(clk16MHz), .D(n53));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1928__i3 (.Q(dti_counter[3]), .C(clk16MHz), .D(n52));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1928__i4 (.Q(dti_counter[4]), .C(clk16MHz), .D(n51));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1928__i5 (.Q(dti_counter[5]), .C(clk16MHz), .D(n50));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1928__i6 (.Q(dti_counter[6]), .C(clk16MHz), .D(n49));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1928__i7 (.Q(dti_counter[7]), .C(clk16MHz), .D(n48));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5699));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_1851 (.I0(\data_in_frame[3] [4]), .I1(n25709), 
            .I2(n25766), .I3(rx_data[4]), .O(n51659));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1851.LUT_INIT = 16'h3a0a;
    SB_CARRY unary_minus_21_add_3_7 (.CI(n45542), .I0(GND_net), .I1(n20), 
            .CO(n45543));
    SB_LUT4 add_1090_3_lut (.I0(GND_net), .I1(n5031), .I2(n5056), .I3(n45777), 
            .O(n440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1852 (.I0(\data_in_frame[3] [3]), .I1(n25709), 
            .I2(n25766), .I3(rx_data[3]), .O(n51663));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1852.LUT_INIT = 16'h3a0a;
    SB_CARRY add_1090_3 (.CI(n45777), .I0(n5031), .I1(n5056), .CO(n45778));
    SB_LUT4 i12_4_lut_adj_1853 (.I0(\data_in_frame[3] [2]), .I1(n25709), 
            .I2(n25766), .I3(rx_data[2]), .O(n51667));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1853.LUT_INIT = 16'h3a0a;
    SB_LUT4 add_1090_2_lut (.I0(GND_net), .I1(n5032), .I2(n5057), .I3(GND_net), 
            .O(n441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1090_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(n4847), .I1(GND_net), .I2(n21), 
            .I3(n45541), .O(n5031)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_156_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n45507));
    SB_CARRY add_1090_2 (.CI(GND_net), .I0(n5032), .I1(n5057), .CO(n45777));
    SB_LUT4 i24720_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n38306), .I2(GND_net), 
            .I3(GND_net), .O(n38310));
    defparam i24720_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_237_8_lut (.I0(current[6]), .I1(duty[9]), .I2(n62401), 
            .I3(n45491), .O(n264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_237_23_lut (.I0(current[15]), .I1(duty[23]), .I2(n62401), 
            .I3(n45506), .O(n249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_23_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n45541), .I0(GND_net), .I1(n21), 
            .CO(n45542));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(n296), .I1(GND_net), .I2(n22_adj_5704), 
            .I3(n45540), .O(n5032)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n45540), .I0(GND_net), .I1(n22_adj_5704), 
            .CO(n45541));
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(n379), .I1(GND_net), .I2(n23), 
            .I3(n45539), .O(n4_adj_5844)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_4_lut_adj_1854 (.I0(\data_in_frame[3] [1]), .I1(n25709), 
            .I2(n25766), .I3(rx_data[1]), .O(n51669));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1854.LUT_INIT = 16'h3a0a;
    SB_CARRY unary_minus_21_add_3_4 (.CI(n45539), .I0(GND_net), .I1(n23), 
            .CO(n45540));
    SB_LUT4 add_237_22_lut (.I0(current[15]), .I1(duty[23]), .I2(n62401), 
            .I3(n45505), .O(n250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_22_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [7]), 
            .O(n52180));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5705), 
            .I3(n45538), .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n45776), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [0]), 
            .O(n52181));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n45538), .I0(GND_net), .I1(n24_adj_5705), 
            .CO(n45539));
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n45775), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n4_adj_5844), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n59192)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n45538));
    SB_CARRY add_237_22 (.CI(n45505), .I0(duty[23]), .I1(n62401), .CO(n45506));
    SB_CARRY unary_minus_19_add_3_14 (.CI(n45775), .I0(GND_net), .I1(n2), 
            .CO(n45776));
    SB_LUT4 add_156_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n45537), .O(n1254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_156_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n45536), .O(n1255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [1]), 
            .O(n52182));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h2300;
    SB_CARRY add_156_32 (.CI(n45536), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n45537));
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5706), 
            .I3(n45774), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_13 (.CI(n45774), .I0(GND_net), .I1(n14_adj_5706), 
            .CO(n45775));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [2]), 
            .O(n52183));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 add_156_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n45535), .O(n1256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_237_21_lut (.I0(current[15]), .I1(duty[22]), .I2(n62401), 
            .I3(n45504), .O(n251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_21_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_237_8 (.CI(n45491), .I0(duty[9]), .I1(n62401), .CO(n45492));
    SB_CARRY add_237_21 (.CI(n45504), .I0(duty[22]), .I1(n62401), .CO(n45505));
    SB_CARRY add_156_31 (.CI(n45535), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n45536));
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5707), 
            .I3(n45773), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_12 (.CI(n45773), .I0(GND_net), .I1(n15_adj_5707), 
            .CO(n45774));
    SB_LUT4 add_237_20_lut (.I0(current[15]), .I1(duty[21]), .I2(n62401), 
            .I3(n45503), .O(n252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_20_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_156_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n45534), .O(n1257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_30 (.CI(n45534), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n45535));
    SB_LUT4 add_156_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n45533), .O(n1258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_237_2_lut (.I0(GND_net), .I1(duty[3]), .I2(n211), .I3(GND_net), 
            .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_20 (.CI(n45503), .I0(duty[21]), .I1(n62401), .CO(n45504));
    SB_LUT4 add_237_7_lut (.I0(current[5]), .I1(duty[8]), .I2(n62401), 
            .I3(n45490), .O(n265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i21453_3_lut (.I0(n25761), .I1(rx_data[7]), .I2(\data_in_frame[5] [7]), 
            .I3(GND_net), .O(n27757));   // verilog/coms.v(94[13:20])
    defparam i21453_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5708), 
            .I3(n45772), .O(n337)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_11 (.CI(n45772), .I0(GND_net), .I1(n16_adj_5708), 
            .CO(n45773));
    SB_LUT4 i13625_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n25766), 
            .I3(GND_net), .O(n27331));   // verilog/coms.v(130[12] 305[6])
    defparam i13625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_237_19_lut (.I0(current[15]), .I1(duty[20]), .I2(n62401), 
            .I3(n45502), .O(n253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_19_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_156_29 (.CI(n45533), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n45534));
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5709), 
            .I3(n45771), .O(n338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_156_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n45532), .O(n1259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_19 (.CI(n45502), .I0(duty[20]), .I1(n62401), .CO(n45503));
    SB_LUT4 add_237_18_lut (.I0(current[15]), .I1(duty[19]), .I2(n62401), 
            .I3(n45501), .O(n254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_18_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13043_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n25761), 
            .I3(GND_net), .O(n26749));   // verilog/coms.v(130[12] 305[6])
    defparam i13043_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_156_28 (.CI(n45532), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n45533));
    SB_CARRY add_237_18 (.CI(n45501), .I0(duty[19]), .I1(n62401), .CO(n45502));
    SB_CARRY unary_minus_19_add_3_10 (.CI(n45771), .I0(GND_net), .I1(n17_adj_5709), 
            .CO(n45772));
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5710), 
            .I3(n45770), .O(n339)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_9 (.CI(n45770), .I0(GND_net), .I1(n18_adj_5710), 
            .CO(n45771));
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5711), 
            .I3(n45769), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13040_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n25761), 
            .I3(GND_net), .O(n26746));   // verilog/coms.v(130[12] 305[6])
    defparam i13040_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_19_add_3_8 (.CI(n45769), .I0(GND_net), .I1(n19_adj_5711), 
            .CO(n45770));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1859 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [3]), 
            .O(n26284));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1859.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5712), 
            .I3(n45768), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_7 (.CI(n45768), .I0(GND_net), .I1(n20_adj_5712), 
            .CO(n45769));
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5713), 
            .I3(n45767), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_156_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n45531), .O(n1260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_27 (.CI(n45531), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n45532));
    SB_CARRY unary_minus_19_add_3_6 (.CI(n45767), .I0(GND_net), .I1(n21_adj_5713), 
            .CO(n45768));
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5714), 
            .I3(n45766), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_5 (.CI(n45766), .I0(GND_net), .I1(n22_adj_5714), 
            .CO(n45767));
    SB_LUT4 add_156_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n45530), .O(n1261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5715), 
            .I3(n45765), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_4 (.CI(n45765), .I0(GND_net), .I1(n23_adj_5715), 
            .CO(n45766));
    SB_CARRY add_156_26 (.CI(n45530), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n45531));
    SB_LUT4 add_156_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n45529), .O(n1262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5716), 
            .I3(n45764), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_3 (.CI(n45764), .I0(GND_net), .I1(n24_adj_5716), 
            .CO(n45765));
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n25_adj_5717), 
            .I3(VCC_net), .O(n59198)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5717), 
            .CO(n45764));
    SB_CARRY add_156_25 (.CI(n45529), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n45530));
    SB_LUT4 add_237_17_lut (.I0(current[15]), .I1(duty[18]), .I2(n62401), 
            .I3(n45500), .O(n255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_17_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5767), .I3(n45763), .O(displacement_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5765), .I3(n45762), .O(displacement_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_156_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n45528), .O(n1263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n45762), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5765), .CO(n45763));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5764), .I3(n45761), .O(displacement_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_17 (.CI(n45500), .I0(duty[18]), .I1(n62401), .CO(n45501));
    SB_CARRY add_156_24 (.CI(n45528), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n45529));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n45761), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5764), .CO(n45762));
    SB_LUT4 add_237_16_lut (.I0(current[15]), .I1(duty[17]), .I2(n62401), 
            .I3(n45499), .O(n256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_16_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_237_7 (.CI(n45490), .I0(duty[8]), .I1(n62401), .CO(n45491));
    SB_LUT4 add_156_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n45527), .O(n1264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5808), .I3(n45760), .O(displacement_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n45760), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5808), .CO(n45761));
    SB_CARRY add_156_23 (.CI(n45527), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n45528));
    SB_CARRY add_237_16 (.CI(n45499), .I0(duty[17]), .I1(n62401), .CO(n45500));
    SB_CARRY add_237_2 (.CI(GND_net), .I0(duty[3]), .I1(n211), .CO(n45486));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5807), .I3(n45759), .O(displacement_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n45759), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5807), .CO(n45760));
    SB_LUT4 add_156_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n45526), .O(n1265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_156_22 (.CI(n45526), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n45527));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5806), .I3(n45758), .O(displacement_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_237_6_lut (.I0(current[4]), .I1(duty[7]), .I2(n62401), 
            .I3(n45489), .O(n266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_237_15_lut (.I0(current[15]), .I1(duty[16]), .I2(n62401), 
            .I3(n45498), .O(n257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i12_4_lut_adj_1860 (.I0(\data_in_frame[2] [4]), .I1(n25713), 
            .I2(n25768), .I3(rx_data[4]), .O(n51673));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1860.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n45758), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5806), .CO(n45759));
    SB_LUT4 i44933_4_lut (.I0(n3543), .I1(\FRAME_MATCHER.i [1]), .I2(n82), 
            .I3(n35696), .O(n59325));   // verilog/coms.v(94[13:20])
    defparam i44933_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5805), .I3(n45757), .O(displacement_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22089_4_lut (.I0(n59325), .I1(n78), .I2(rx_data[3]), .I3(\data_in_frame[2] [3]), 
            .O(n35720));   // verilog/coms.v(94[13:20])
    defparam i22089_4_lut.LUT_INIT = 16'hfac0;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n45757), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5805), .CO(n45758));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5804), .I3(n45756), .O(displacement_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22090_3_lut (.I0(n35720), .I1(\data_in_frame[2] [3]), .I2(reset), 
            .I3(GND_net), .O(n27317));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1861 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [4]), 
            .O(n26283));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1861.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1862 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [5]), 
            .O(n52184));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1862.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1863 (.I0(\data_in_frame[2] [1]), .I1(n25713), 
            .I2(n25768), .I3(rx_data[1]), .O(n51677));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1863.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n45756), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5804), .CO(n45757));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5803), .I3(n45755), .O(displacement_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1864 (.I0(\FRAME_MATCHER.i [0]), .I1(n10), .I2(GND_net), 
            .I3(GND_net), .O(n82));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1864.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [6]), 
            .O(n26281));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [7]), 
            .O(n52185));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1867 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [0]), 
            .O(n52186));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1867.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [1]), 
            .O(n52187));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n45755), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5803), .CO(n45756));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5801), .I3(n45754), .O(displacement_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n45754), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5801), .CO(n45755));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [2]), 
            .O(n26277));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5800), .I3(n45753), .O(displacement_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n45753), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5800), .CO(n45754));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [3]), 
            .O(n26276));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut (.I0(n9582), .I1(n419), .I2(current[15]), 
            .I3(duty[23]), .O(n62835));
    defparam n9582_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [4]), 
            .O(n26275));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 n62835_bdd_4_lut (.I0(n62835), .I1(duty[22]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam n62835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5799), .I3(n45752), .O(displacement_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n45752), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5799), .CO(n45753));
    SB_LUT4 i2_3_lut (.I0(n35727), .I1(n38302), .I2(\FRAME_MATCHER.i [0]), 
            .I3(GND_net), .O(n78));
    defparam i2_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [5]), 
            .O(n52188));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [6]), 
            .O(n52189));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1874 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [7]), 
            .O(n52190));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1874.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47859 (.I0(n9582), .I1(n420), .I2(current[15]), 
            .I3(duty[23]), .O(n62829));
    defparam n9582_bdd_4_lut_47859.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1875 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5817));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1875.LUT_INIT = 16'h6666;
    SB_LUT4 i14275_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [6]), 
            .O(n27981));   // verilog/coms.v(130[12] 305[6])
    defparam i14275_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [0]), 
            .O(n52191));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5798), .I3(n45751), .O(displacement_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n45751), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5798), .CO(n45752));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5797), .I3(n45750), .O(displacement_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n45750), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5797), .CO(n45751));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5786), .I3(n45749), .O(displacement_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1877 (.I0(\data_in_frame[2] [0]), .I1(n25713), 
            .I2(n25768), .I3(rx_data[0]), .O(n51681));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1877.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52424), .O(n52427));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [1]), 
            .O(n52192));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [2]), 
            .O(n52193));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n45749), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5786), .CO(n45750));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [3]), 
            .O(n52194));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5785), .I3(n45748), .O(displacement_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n45748), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5785), .CO(n45749));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5784), .I3(n45747), .O(displacement_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n45747), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5784), .CO(n45748));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5783), .I3(n45746), .O(displacement_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [4]), 
            .O(n52195));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [5]), 
            .O(n52196));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n45746), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5783), .CO(n45747));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5782), .I3(n45745), .O(displacement_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [6]), 
            .O(n52197));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 i13037_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n25761), 
            .I3(GND_net), .O(n26743));   // verilog/coms.v(130[12] 305[6])
    defparam i13037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n62829_bdd_4_lut (.I0(n62829), .I1(duty[21]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam n62829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[24] [7]), 
            .O(n52198));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 i24561_2_lut_2_lut (.I0(duty[10]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5047));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24561_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n45745), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5782), .CO(n45746));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5780), .I3(n45744), .O(displacement_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n45744), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5780), .CO(n45745));
    SB_LUT4 add_156_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n45525), .O(n1266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5779), .I3(n45743), .O(displacement_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n45743), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5779), .CO(n45744));
    SB_LUT4 dti_counter_1928_add_4_9_lut (.I0(n59312), .I1(n37855), .I2(dti_counter[7]), 
            .I3(n46065), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 dti_counter_1928_add_4_8_lut (.I0(n59311), .I1(n37855), .I2(dti_counter[6]), 
            .I3(n46064), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1928_add_4_8 (.CI(n46064), .I0(n37855), .I1(dti_counter[6]), 
            .CO(n46065));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5763), .I3(n45742), .O(displacement_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_237_15 (.CI(n45498), .I0(duty[16]), .I1(n62401), .CO(n45499));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n45742), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5763), .CO(n45743));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [0]), 
            .O(n52199));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5762), .I3(n45741), .O(displacement_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1928_add_4_7_lut (.I0(n59310), .I1(n37855), .I2(dti_counter[5]), 
            .I3(n46063), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1928_add_4_7 (.CI(n46063), .I0(n37855), .I1(dti_counter[5]), 
            .CO(n46064));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n45741), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5762), .CO(n45742));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5761), .I3(VCC_net), .O(displacement_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_237_14_lut (.I0(current[15]), .I1(duty[15]), .I2(n62401), 
            .I3(n45497), .O(n258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_237_14_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5761), .CO(n45741));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [1]), 
            .O(n52200));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 dti_counter_1928_add_4_6_lut (.I0(n59309), .I1(n37855), .I2(dti_counter[4]), 
            .I3(n46062), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1928_add_4_6 (.CI(n46062), .I0(n37855), .I1(dti_counter[4]), 
            .CO(n46063));
    SB_LUT4 dti_counter_1928_add_4_5_lut (.I0(n59308), .I1(n37855), .I2(dti_counter[3]), 
            .I3(n46061), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1928_add_4_5 (.CI(n46061), .I0(n37855), .I1(dti_counter[3]), 
            .CO(n46062));
    SB_LUT4 dti_counter_1928_add_4_4_lut (.I0(n59307), .I1(n37855), .I2(dti_counter[2]), 
            .I3(n46060), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1928_add_4_4 (.CI(n46060), .I0(n37855), .I1(dti_counter[2]), 
            .CO(n46061));
    SB_CARRY add_237_14 (.CI(n45497), .I0(duty[15]), .I1(n62401), .CO(n45498));
    SB_LUT4 dti_counter_1928_add_4_3_lut (.I0(n59306), .I1(n37855), .I2(dti_counter[1]), 
            .I3(n46059), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY add_156_21 (.CI(n45525), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n45526));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [2]), 
            .O(n52201));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_CARRY dti_counter_1928_add_4_3 (.CI(n46059), .I0(n37855), .I1(dti_counter[1]), 
            .CO(n46060));
    SB_LUT4 add_156_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n45524), .O(n1267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1928_add_4_2_lut (.I0(n59279), .I1(n2916), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1928_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_1928_add_4_2 (.CI(VCC_net), .I0(n2916), .I1(dti_counter[0]), 
            .CO(n46059));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [3]), 
            .O(n52202));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_CARRY add_156_20 (.CI(n45524), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n45525));
    SB_LUT4 add_156_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n45523), .O(n1268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_156_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [4]), 
            .O(n52203));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47854 (.I0(n9582), .I1(n421), .I2(current[15]), 
            .I3(duty[23]), .O(n62823));
    defparam n9582_bdd_4_lut_47854.LUT_INIT = 16'he4aa;
    SB_LUT4 i14066_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n52435), 
            .I3(GND_net), .O(n27772));   // verilog/coms.v(130[12] 305[6])
    defparam i14066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [5]), 
            .O(n52204));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [6]), 
            .O(n52205));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_CARRY add_237_6 (.CI(n45489), .I0(duty[7]), .I1(n62401), .CO(n45490));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[25] [7]), 
            .O(n52206));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[3] [1]), 
            .O(n52207));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[3] [3]), 
            .O(n52208));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[3] [4]), 
            .O(n52209));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[3] [6]), 
            .O(n52210));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 n62823_bdd_4_lut (.I0(n62823), .I1(duty[20]), .I2(n250), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam n62823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[3] [7]), 
            .O(n52211));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [0]), 
            .O(n52212));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [1]), 
            .O(n26215));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [2]), 
            .O(n52213));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [3]), 
            .O(n26213));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [4]), 
            .O(n52214));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [5]), 
            .O(n52215));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 mux_15_i1_3_lut (.I0(current[0]), .I1(n1788), .I2(n209), .I3(GND_net), 
            .O(n270));   // verilog/TinyFPGA_B.v(112[16] 114[10])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [6]), 
            .O(n26207));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i24562_2_lut_2_lut (.I0(duty[9]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5048));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24562_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [7]), 
            .O(n52216));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47759 (.I0(n9582), .I1(n440), .I2(current[1]), 
            .I3(duty[23]), .O(n62709));
    defparam n9582_bdd_4_lut_47759.LUT_INIT = 16'he4aa;
    SB_LUT4 i24544_2_lut_2_lut (.I0(duty[23]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5034));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24544_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i41925_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56825));
    defparam i41925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41926_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56826));
    defparam i41926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [0]), 
            .O(n52300));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i41689_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56589));
    defparam i41689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41688_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56588));
    defparam i41688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[0] [4]), 
            .O(n52299));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [1]), 
            .O(n52298));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [2]), 
            .O(n52297));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [3]), 
            .O(n52296));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_67[19]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13486_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n54720), .I3(GND_net), .O(n27192));   // verilog/coms.v(130[12] 305[6])
    defparam i13486_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_252_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_67[20]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [4]), 
            .O(n52295));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [5]), 
            .O(n26402));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [6]), 
            .O(n52294));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 mux_250_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_67[21]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [7]), 
            .O(n26400));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 mux_252_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_67[14]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [0]), 
            .O(n26399));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [1]), 
            .O(n52293));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 i24565_2_lut_2_lut (.I0(duty[8]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5049));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24565_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mux_252_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22453_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_67[22]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(n9_adj_5816));
    defparam i22453_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1917 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [2]), 
            .O(n52292));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1917.LUT_INIT = 16'h2300;
    SB_LUT4 i24569_2_lut_2_lut (.I0(duty[7]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5050));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24569_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24570_2_lut_2_lut (.I0(duty[6]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5051));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24570_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [3]), 
            .O(n52291));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5761));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [4]), 
            .O(n52290));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5762));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5763));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [5]), 
            .O(n52289));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [6]), 
            .O(n52288));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h2300;
    SB_LUT4 i24267_2_lut (.I0(n20251), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n37855));
    defparam i24267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5779));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_252_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_67[23]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5780));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [7]), 
            .O(n52287));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [0]), 
            .O(n26391));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5782));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i44665_3_lut_4_lut (.I0(r_Clock_Count_adj_5934[3]), .I1(o_Rx_DV_N_3464[3]), 
            .I2(o_Rx_DV_N_3464[2]), .I3(r_Clock_Count_adj_5934[2]), .O(n59565));   // verilog/uart_tx.v(117[17:57])
    defparam i44665_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5783));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5784));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5785));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13034_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n25761), 
            .I3(GND_net), .O(n26740));   // verilog/coms.v(130[12] 305[6])
    defparam i13034_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1071_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5934[3]), 
            .I1(o_Rx_DV_N_3464[3]), .I2(o_Rx_DV_N_3464[2]), .I3(GND_net), 
            .O(n6_adj_5820));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1071_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i13031_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n25761), 
            .I3(GND_net), .O(n26737));   // verilog/coms.v(130[12] 305[6])
    defparam i13031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5786));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5797));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13028_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n25761), 
            .I3(GND_net), .O(n26734));   // verilog/coms.v(130[12] 305[6])
    defparam i13028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5798));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [1]), 
            .O(n26390));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [2]), 
            .O(n52286));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 i13025_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n25761), 
            .I3(GND_net), .O(n26731));   // verilog/coms.v(130[12] 305[6])
    defparam i13025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [3]), 
            .O(n52285));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5799));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(duty[7]), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(duty[6]), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(duty[9]), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(duty[8]), .I1(n338), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i7_2_lut (.I0(duty[3]), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(duty[4]), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(duty[5]), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i5_2_lut (.I0(duty[2]), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45267_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n60167));
    defparam i45267_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n342), .I1(n338), .I2(n17), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i6_3_lut (.I0(n344), .I1(n343), .I2(n7), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n8), .I1(n337), .I2(n19), .I3(GND_net), 
            .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41414_3_lut (.I0(duty[19]), .I1(duty[21]), .I2(n330), .I3(GND_net), 
            .O(n56302));
    defparam i41414_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i41418_3_lut (.I0(duty[14]), .I1(duty[17]), .I2(n330), .I3(GND_net), 
            .O(n56306));
    defparam i41418_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i41572_4_lut (.I0(duty[20]), .I1(n56302), .I2(duty[22]), .I3(n330), 
            .O(n56463));
    defparam i41572_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 LessThan_20_i4_3_lut (.I0(n59198), .I1(n345), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [4]), 
            .O(n52284));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h2300;
    SB_LUT4 i46703_3_lut (.I0(n4), .I1(n341), .I2(n11), .I3(GND_net), 
            .O(n61603));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i46703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46704_3_lut (.I0(n61603), .I1(n340), .I2(n13), .I3(GND_net), 
            .O(n61604));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i46704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45254_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n60167), 
            .O(n60154));
    defparam i45254_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47035_4_lut (.I0(n16), .I1(n6), .I2(n19), .I3(n60152), 
            .O(n61935));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i47035_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45555_3_lut (.I0(n61604), .I1(n339), .I2(n15), .I3(GND_net), 
            .O(n60455));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i45555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47202_4_lut (.I0(n60455), .I1(n61935), .I2(n19), .I3(n60154), 
            .O(n62102));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i47202_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47203_3_lut (.I0(n62102), .I1(n336), .I2(duty[10]), .I3(GND_net), 
            .O(n62103));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i47203_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47186_3_lut (.I0(n62103), .I1(n335), .I2(duty[11]), .I3(GND_net), 
            .O(n62086));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i47186_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_20_i26_3_lut (.I0(n62086), .I1(n334), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7_4_lut_adj_1928 (.I0(duty[18]), .I1(n26), .I2(n330), .I3(duty[23]), 
            .O(n20_adj_5859));
    defparam i7_4_lut_adj_1928.LUT_INIT = 16'h2100;
    SB_LUT4 i11_4_lut (.I0(n330), .I1(n56463), .I2(n56306), .I3(duty[13]), 
            .O(n24_adj_5858));
    defparam i11_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i44752_4_lut (.I0(duty[16]), .I1(n20_adj_5859), .I2(duty[15]), 
            .I3(n330), .O(n59349));
    defparam i44752_4_lut.LUT_INIT = 16'h8004;
    SB_LUT4 i14_4_lut_adj_1929 (.I0(n59349), .I1(pwm_setpoint_23__N_183), 
            .I2(n296), .I3(n24_adj_5858), .O(n9582));
    defparam i14_4_lut_adj_1929.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [5]), 
            .O(n52283));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1931 (.I0(n33996), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n125));
    defparam i1_2_lut_adj_1931.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1932 (.I0(n33996), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n198));
    defparam i1_2_lut_adj_1932.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [6]), 
            .O(n52282));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1934 (.I0(n33996), .I1(Ki[3]), .I2(GND_net), 
            .I3(GND_net), .O(n271));
    defparam i1_2_lut_adj_1934.LUT_INIT = 16'h8888;
    SB_LUT4 i47296_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n37857), .I3(GND_net), .O(n25013));
    defparam i47296_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i1_2_lut_adj_1935 (.I0(n33996), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5832));
    defparam i1_2_lut_adj_1935.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [7]), 
            .O(n26384));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1937 (.I0(n33996), .I1(Ki[5]), .I2(GND_net), 
            .I3(GND_net), .O(n417));
    defparam i1_2_lut_adj_1937.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [0]), 
            .O(n52281));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 i44676_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n59196));
    defparam i44676_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i24381_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n37857), .I3(GND_net), .O(n37969));
    defparam i24381_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1939 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(delay_counter[14]), .O(n4_adj_5840));
    defparam i1_2_lut_4_lut_adj_1939.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52434), .O(n52435));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut_adj_1940.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1941 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52430), .O(n52432));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut_adj_1941.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_1942 (.I0(n33996), .I1(Ki[6]), .I2(GND_net), 
            .I3(GND_net), .O(n490));
    defparam i1_2_lut_adj_1942.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5800));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5801));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5803));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5804));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5805));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5806));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5807));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5808));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9582_bdd_4_lut_47849 (.I0(n9582), .I1(n422), .I2(current[15]), 
            .I3(duty[23]), .O(n62817));
    defparam n9582_bdd_4_lut_47849.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5764));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5765));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5767));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n22887), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5728));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5717));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5716));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n62817_bdd_4_lut (.I0(n62817), .I1(duty[19]), .I2(n251), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[19]));
    defparam n62817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5711));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5710));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1943 (.I0(control_mode[0]), .I1(n22887), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_5727));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_3_lut_adj_1943.LUT_INIT = 16'hfefe;
    SB_LUT4 i14273_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [4]), 
            .O(n27979));   // verilog/coms.v(130[12] 305[6])
    defparam i14273_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5709));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5708));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(duty[0]), .I1(duty[23]), .I2(duty[1]), .I3(duty[2]), 
            .O(n211));   // verilog/TinyFPGA_B.v(111[25:31])
    defparam i14_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5707));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5706));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_1_lut (.I0(current[15]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5705));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9582_bdd_4_lut_47844 (.I0(n9582), .I1(n423), .I2(current[15]), 
            .I3(duty[23]), .O(n62811));
    defparam n9582_bdd_4_lut_47844.LUT_INIT = 16'he4aa;
    SB_LUT4 i13547_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[3]), 
            .I2(counter_adj_5947[0]), .I3(n22918), .O(n27253));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13547_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13549_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[4]), 
            .I2(counter_adj_5947[0]), .I3(n22915), .O(n27255));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13549_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13550_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[5]), 
            .I2(counter_adj_5947[0]), .I3(n22915), .O(n27256));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13550_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[5] [7]), .I3(n10_adj_5729), .O(n1513));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13551_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[6]), 
            .I2(counter_adj_5947[0]), .I3(n22907), .O(n27257));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13551_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [0]), .O(n23427));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1944 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[12] [5]), .I3(\data_out_frame[14] [7]), 
            .O(n53122));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1944.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5704));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13553_4_lut (.I0(state_7__N_4100[3]), .I1(data_adj_5912[7]), 
            .I2(counter_adj_5947[0]), .I3(n22907), .O(n27259));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13553_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_3_lut_adj_1945 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(n52979), .I3(GND_net), .O(n8_adj_5720));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1945.LUT_INIT = 16'h9696;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1088_i1_4_lut (.I0(n59192), .I1(duty[0]), .I2(n296), .I3(n356), 
            .O(n5057));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam mux_1088_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i5_3_lut_4_lut_adj_1946 (.I0(\data_out_frame[7] [1]), .I1(n10_adj_5845), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [2]), 
            .O(n47380));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1946.LUT_INIT = 16'h6996;
    SB_LUT4 i24575_2_lut (.I0(duty[1]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5056));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24575_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13621_3_lut_4_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(rx_data[7]), 
            .I2(reset), .I3(n78), .O(n27327));   // verilog/coms.v(130[12] 305[6])
    defparam i13621_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i13615_3_lut_4_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n78), .O(n27321));   // verilog/coms.v(130[12] 305[6])
    defparam i13615_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i13_4_lut_adj_1947 (.I0(\data_in_frame[11] [7]), .I1(n10_adj_5778), 
            .I2(n25750), .I3(n52362), .O(n51551));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1947.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1948 (.I0(\data_in_frame[11] [6]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[6]), .O(n51553));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1948.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1949 (.I0(\data_in_frame[11] [5]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[5]), .O(n51555));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1949.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1950 (.I0(\data_in_frame[11] [4]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[4]), .O(n51557));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1950.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1951 (.I0(\data_in_frame[11] [3]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[3]), .O(n51559));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1951.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_1952 (.I0(\data_in_frame[11] [2]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[2]), .O(n51561));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1952.LUT_INIT = 16'h3a0a;
    SB_LUT4 i11_4_lut_adj_1953 (.I0(\data_in_frame[11] [1]), .I1(n38310), 
            .I2(n25750), .I3(rx_data[1]), .O(n51585));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1953.LUT_INIT = 16'hca0a;
    SB_LUT4 i13606_3_lut_4_lut_4_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), 
            .I2(reset), .I3(n78), .O(n27312));   // verilog/coms.v(130[12] 305[6])
    defparam i13606_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i13_4_lut_adj_1954 (.I0(\data_in_frame[11] [0]), .I1(n53300), 
            .I2(n25750), .I3(rx_data[0]), .O(n51563));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1954.LUT_INIT = 16'h3a0a;
    SB_LUT4 i47501_1_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n54039), 
            .I3(n54035), .O(n62401));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i47501_1_lut_4_lut.LUT_INIT = 16'h4c5d;
    SB_LUT4 i1_4_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n54039), 
            .I3(n54035), .O(n209));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb3a2;
    SB_LUT4 i2_3_lut_adj_1955 (.I0(\FRAME_MATCHER.i [0]), .I1(n38306), .I2(n10_adj_5778), 
            .I3(GND_net), .O(n25707));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_adj_1955.LUT_INIT = 16'hfbfb;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5747));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i4900_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_331));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i4900_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i4902_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_348));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i4902_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i4904_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_353));
    defparam i4904_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i4906_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_362));
    defparam i4906_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i24545_2_lut_2_lut (.I0(duty[22]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5035));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24545_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i44907_2_lut_4_lut (.I0(current[8]), .I1(duty[8]), .I2(current[4]), 
            .I3(duty[4]), .O(n59807));
    defparam i44907_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5745));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13081_3_lut_4_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26787));   // verilog/coms.v(130[12] 305[6])
    defparam i13081_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13080_3_lut_4_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26786));   // verilog/coms.v(130[12] 305[6])
    defparam i13080_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13076_3_lut_4_lut (.I0(deadband[0]), .I1(\data_in_frame[16] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26782));   // verilog/coms.v(130[12] 305[6])
    defparam i13076_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n62811_bdd_4_lut (.I0(n62811), .I1(duty[18]), .I2(n252), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[18]));
    defparam n62811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14272_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[22] [3]), 
            .O(n27978));   // verilog/coms.v(130[12] 305[6])
    defparam i14272_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_252_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(motor_state_23__N_67[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_252_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_250_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_67[15]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13063_3_lut_4_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26769));   // verilog/coms.v(130[12] 305[6])
    defparam i13063_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13062_3_lut_4_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26768));   // verilog/coms.v(130[12] 305[6])
    defparam i13062_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_4_lut_adj_1956 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n37857), .O(n50941));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_4_lut_4_lut_adj_1956.LUT_INIT = 16'hb1f1;
    SB_LUT4 i2_3_lut_adj_1957 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_192));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_3_lut_adj_1957.LUT_INIT = 16'h0202;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5862));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1958 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_184[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1958.LUT_INIT = 16'h1414;
    SB_LUT4 i14264_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [3]), 
            .O(n27970));   // verilog/coms.v(130[12] 305[6])
    defparam i14264_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14262_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[21] [1]), 
            .O(n27968));   // verilog/coms.v(130[12] 305[6])
    defparam i14262_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38451_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n38306), 
            .I2(n10_adj_5778), .I3(GND_net), .O(n53300));
    defparam i38451_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i12464_2_lut (.I0(n24962), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n26176));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i12464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47258_4_lut (.I0(commutation_state[1]), .I1(n20251), .I2(dti), 
            .I3(commutation_state[2]), .O(n24962));
    defparam i47258_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i41764_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56664));
    defparam i41764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41763_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56663));
    defparam i41763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41765_4_lut (.I0(n56664), .I1(n62472), .I2(n47529), .I3(n47509), 
            .O(n56665));
    defparam i41765_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 n9582_bdd_4_lut_47839 (.I0(n9582), .I1(n424), .I2(current[15]), 
            .I3(duty[23]), .O(n62805));
    defparam n9582_bdd_4_lut_47839.LUT_INIT = 16'he4aa;
    SB_LUT4 i13430_3_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(n25739), .I3(GND_net), .O(n27136));   // verilog/coms.v(130[12] 305[6])
    defparam i13430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n62805_bdd_4_lut (.I0(n62805), .I1(duty[17]), .I2(n253), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[17]));
    defparam n62805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9582_bdd_4_lut_47834 (.I0(n9582), .I1(n425), .I2(current[15]), 
            .I3(duty[23]), .O(n62799));
    defparam n9582_bdd_4_lut_47834.LUT_INIT = 16'he4aa;
    SB_LUT4 i45252_2_lut_4_lut (.I0(duty[8]), .I1(n338), .I2(duty[4]), 
            .I3(n342), .O(n60152));
    defparam i45252_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i13423_3_lut_4_lut (.I0(deadband[1]), .I1(\data_in_frame[16] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27129));   // verilog/coms.v(130[12] 305[6])
    defparam i13423_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13422_3_lut_4_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27128));   // verilog/coms.v(130[12] 305[6])
    defparam i13422_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n62799_bdd_4_lut (.I0(n62799), .I1(duty[16]), .I2(n254), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[16]));
    defparam n62799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13421_3_lut_4_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27127));   // verilog/coms.v(130[12] 305[6])
    defparam i13421_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13420_3_lut_4_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27126));   // verilog/coms.v(130[12] 305[6])
    defparam i13420_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i30968_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5724), .I3(n15_adj_5728), .O(n3_adj_5841));
    defparam i30968_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14256_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [3]), 
            .O(n27962));   // verilog/coms.v(130[12] 305[6])
    defparam i14256_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30969_3_lut (.I0(encoder0_position_scaled[16]), .I1(n3_adj_5841), 
            .I2(n15_adj_5727), .I3(GND_net), .O(n5_adj_5839));
    defparam i30969_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i24268_1_lut_2_lut (.I0(n20251), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n2916));
    defparam i24268_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i14254_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[20] [1]), 
            .O(n27960));   // verilog/coms.v(130[12] 305[6])
    defparam i14254_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_4_lut_adj_1959 (.I0(reset), .I1(n25705), .I2(\data_in_frame[0] [7]), 
            .I3(rx_data[7]), .O(n51817));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut_adj_1959.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13427_3_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(n25739), .I3(GND_net), .O(n27133));   // verilog/coms.v(130[12] 305[6])
    defparam i13427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24574_2_lut (.I0(duty[2]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5055));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24574_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24573_2_lut (.I0(duty[3]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5054));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24573_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13747_3_lut (.I0(current[10]), .I1(data_adj_5920[10]), .I2(n25021), 
            .I3(GND_net), .O(n27453));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13748_3_lut (.I0(current[9]), .I1(data_adj_5920[9]), .I2(n25021), 
            .I3(GND_net), .O(n27454));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9582_bdd_4_lut_47829 (.I0(n9582), .I1(n426), .I2(current[15]), 
            .I3(duty[23]), .O(n62793));
    defparam n9582_bdd_4_lut_47829.LUT_INIT = 16'he4aa;
    SB_LUT4 i13749_3_lut (.I0(current[8]), .I1(data_adj_5920[8]), .I2(n25021), 
            .I3(GND_net), .O(n27455));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13750_3_lut (.I0(current[7]), .I1(data_adj_5920[7]), .I2(n25021), 
            .I3(GND_net), .O(n27456));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13751_3_lut (.I0(current[6]), .I1(data_adj_5920[6]), .I2(n25021), 
            .I3(GND_net), .O(n27457));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13752_3_lut (.I0(current[5]), .I1(data_adj_5920[5]), .I2(n25021), 
            .I3(GND_net), .O(n27458));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13753_3_lut (.I0(current[4]), .I1(data_adj_5920[4]), .I2(n25021), 
            .I3(GND_net), .O(n27459));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13754_3_lut (.I0(current[3]), .I1(data_adj_5920[3]), .I2(n25021), 
            .I3(GND_net), .O(n27460));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13755_3_lut (.I0(current[2]), .I1(data_adj_5920[2]), .I2(n25021), 
            .I3(GND_net), .O(n27461));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13756_3_lut (.I0(current[1]), .I1(data_adj_5920[1]), .I2(n25021), 
            .I3(GND_net), .O(n27462));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13757_3_lut (.I0(baudrate[31]), .I1(data_adj_5912[7]), .I2(n25293), 
            .I3(GND_net), .O(n27463));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13758_3_lut (.I0(baudrate[30]), .I1(data_adj_5912[6]), .I2(n25293), 
            .I3(GND_net), .O(n27464));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13759_3_lut (.I0(baudrate[29]), .I1(data_adj_5912[5]), .I2(n25293), 
            .I3(GND_net), .O(n27465));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n62793_bdd_4_lut (.I0(n62793), .I1(duty[15]), .I2(n255), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[15]));
    defparam n62793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9582_bdd_4_lut_47824 (.I0(n9582), .I1(n427), .I2(current[15]), 
            .I3(duty[23]), .O(n62787));
    defparam n9582_bdd_4_lut_47824.LUT_INIT = 16'he4aa;
    SB_LUT4 i13760_3_lut (.I0(baudrate[28]), .I1(data_adj_5912[4]), .I2(n25293), 
            .I3(GND_net), .O(n27466));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13761_3_lut (.I0(baudrate[27]), .I1(data_adj_5912[3]), .I2(n25293), 
            .I3(GND_net), .O(n27467));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13762_3_lut (.I0(baudrate[26]), .I1(data_adj_5912[2]), .I2(n25293), 
            .I3(GND_net), .O(n27468));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13763_3_lut (.I0(baudrate[25]), .I1(data_adj_5912[1]), .I2(n25293), 
            .I3(GND_net), .O(n27469));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13764_3_lut (.I0(baudrate[24]), .I1(data_adj_5912[0]), .I2(n25293), 
            .I3(GND_net), .O(n27470));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n62787_bdd_4_lut (.I0(n62787), .I1(duty[14]), .I2(n256), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[14]));
    defparam n62787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9582_bdd_4_lut_47819 (.I0(n9582), .I1(n428), .I2(current[15]), 
            .I3(duty[23]), .O(n62781));
    defparam n9582_bdd_4_lut_47819.LUT_INIT = 16'he4aa;
    SB_LUT4 i13776_3_lut (.I0(baudrate[12]), .I1(data_adj_5912[4]), .I2(n25295), 
            .I3(GND_net), .O(n27482));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13777_3_lut (.I0(baudrate[11]), .I1(data_adj_5912[3]), .I2(n25295), 
            .I3(GND_net), .O(n27483));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13778_3_lut (.I0(baudrate[10]), .I1(data_adj_5912[2]), .I2(n25295), 
            .I3(GND_net), .O(n27484));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13779_3_lut (.I0(baudrate[9]), .I1(data_adj_5912[1]), .I2(n25295), 
            .I3(GND_net), .O(n27485));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13780_3_lut (.I0(baudrate[8]), .I1(data_adj_5912[0]), .I2(n25295), 
            .I3(GND_net), .O(n27486));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24572_2_lut (.I0(duty[4]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5053));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24572_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 n62781_bdd_4_lut (.I0(n62781), .I1(duty[13]), .I2(n257), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[13]));
    defparam n62781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13418_3_lut_4_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27124));   // verilog/coms.v(130[12] 305[6])
    defparam i13418_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13417_3_lut_4_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27123));   // verilog/coms.v(130[12] 305[6])
    defparam i13417_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13416_3_lut_4_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27122));   // verilog/coms.v(130[12] 305[6])
    defparam i13416_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13415_3_lut_4_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27121));   // verilog/coms.v(130[12] 305[6])
    defparam i13415_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13414_3_lut_4_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27120));   // verilog/coms.v(130[12] 305[6])
    defparam i13414_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_250_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_67[17]), 
            .I2(n15_adj_5727), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_250_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5742));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5741));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5738));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5739));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5746));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5744));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5743));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i5_2_lut (.I0(current[2]), .I1(duty[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5748));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24546_2_lut_2_lut (.I0(duty[21]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5036));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24546_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i44936_4_lut (.I0(n11_adj_5743), .I1(n9_adj_5744), .I2(n7_adj_5746), 
            .I3(n5_adj_5748), .O(n59836));
    defparam i44936_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i4910_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_376));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i4910_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i4908_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_367));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i4908_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5745), .I1(duty[9]), .I2(n19_adj_5738), 
            .I3(GND_net), .O(n16_adj_5740));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 n9582_bdd_4_lut_47814 (.I0(n9582), .I1(n429), .I2(current[15]), 
            .I3(duty[23]), .O(n62775));
    defparam n9582_bdd_4_lut_47814.LUT_INIT = 16'he4aa;
    SB_LUT4 i46691_3_lut (.I0(n4_adj_5749), .I1(duty[5]), .I2(n11_adj_5743), 
            .I3(GND_net), .O(n61591));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i46691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n62775_bdd_4_lut (.I0(n62775), .I1(duty[12]), .I2(n258), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[12]));
    defparam n62775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46692_3_lut (.I0(n61591), .I1(duty[6]), .I2(n13_adj_5742), 
            .I3(GND_net), .O(n61592));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i46692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44909_4_lut (.I0(n17_adj_5739), .I1(n15_adj_5741), .I2(n13_adj_5742), 
            .I3(n59836), .O(n59809));
    defparam i44909_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46799_4_lut (.I0(n16_adj_5740), .I1(n6_adj_5747), .I2(n19_adj_5738), 
            .I3(n59807), .O(n61699));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i46799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45571_3_lut (.I0(n61592), .I1(duty[7]), .I2(n15_adj_5741), 
            .I3(GND_net), .O(n60471));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i45571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47120_4_lut (.I0(n60471), .I1(n61699), .I2(n19_adj_5738), 
            .I3(n59809), .O(n62020));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i47120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47121_3_lut (.I0(n62020), .I1(duty[10]), .I2(current[10]), 
            .I3(GND_net), .O(n62021));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i47121_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47054_3_lut (.I0(n62021), .I1(duty[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5737));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i47054_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut_adj_1960 (.I0(duty[14]), .I1(n24_adj_5737), .I2(duty[12]), 
            .I3(duty[13]), .O(n54842));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1960.LUT_INIT = 16'hfffe;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i3_4_lut_adj_1961 (.I0(duty[14]), .I1(n24_adj_5737), .I2(duty[12]), 
            .I3(duty[13]), .O(n54861));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1961.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1962 (.I0(duty[15]), .I1(current[15]), .I2(n54861), 
            .I3(n54842), .O(n32));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1962.LUT_INIT = 16'hb3a2;
    SB_LUT4 i24613_2_lut_2_lut (.I0(n296), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n5010));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i24613_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i45345_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n59279));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i45345_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i44853_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n59306));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44853_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i3_4_lut_adj_1963 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n55011));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1963.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1964 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n55054));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1964.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1965 (.I0(duty[19]), .I1(current[15]), .I2(n55054), 
            .I3(n55011), .O(n40_adj_5736));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1965.LUT_INIT = 16'hb3a2;
    SB_LUT4 i44738_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n59307));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44738_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i44687_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n59308));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44687_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i44878_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n59309));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44878_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i3_4_lut_adj_1966 (.I0(duty[22]), .I1(n40_adj_5736), .I2(duty[20]), 
            .I3(duty[21]), .O(n54035));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1966.LUT_INIT = 16'hfffe;
    SB_LUT4 i13438_3_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(n25739), .I3(GND_net), .O(n27144));   // verilog/coms.v(130[12] 305[6])
    defparam i13438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1967 (.I0(duty[22]), .I1(n40_adj_5736), .I2(duty[20]), 
            .I3(duty[21]), .O(n54039));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1967.LUT_INIT = 16'h8000;
    SB_LUT4 i44737_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n59310));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44737_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 n9582_bdd_4_lut_47809 (.I0(n9582), .I1(n430), .I2(current[11]), 
            .I3(duty[23]), .O(n62769));
    defparam n9582_bdd_4_lut_47809.LUT_INIT = 16'he4aa;
    SB_LUT4 i44736_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n59311));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44736_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_3_lut_adj_1968 (.I0(n38306), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n10), .I3(GND_net), .O(n25713));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1968.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n78), .I2(GND_net), .I3(GND_net), 
            .O(n25768));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 n62769_bdd_4_lut (.I0(n62769), .I1(duty[11]), .I2(n259), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[11]));
    defparam n62769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1969 (.I0(\data_out_frame[12] [7]), .I1(n53113), 
            .I2(n52939), .I3(n52584), .O(n23594));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1969.LUT_INIT = 16'h6996;
    SB_LUT4 i13494_3_lut (.I0(\data_in_frame[18] [1]), .I1(rx_data[1]), 
            .I2(n54720), .I3(GND_net), .O(n27200));   // verilog/coms.v(130[12] 305[6])
    defparam i13494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13497_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n54720), .I3(GND_net), .O(n27203));   // verilog/coms.v(130[12] 305[6])
    defparam i13497_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(100[12:26])
    defparam i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1970 (.I0(n68), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n10), .O(n25766));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_adj_1970.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_adj_1971 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53092));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1971.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1972 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5857));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1972.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n53092), .I1(n52922), .I2(n53125), .I3(n6_adj_5857), 
            .O(n52564));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1973 (.I0(n10), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n38306), .I3(GND_net), .O(n25709));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1973.LUT_INIT = 16'hbfbf;
    SB_LUT4 i4_4_lut_adj_1974 (.I0(\data_out_frame[9] [2]), .I1(n1130), 
            .I2(n52741), .I3(n23531), .O(n10_adj_5815));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1974.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1975 (.I0(n23427), .I1(n10_adj_5815), .I2(\data_out_frame[6] [6]), 
            .I3(GND_net), .O(n53035));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1975.LUT_INIT = 16'h9696;
    SB_LUT4 i13413_3_lut_4_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27119));   // verilog/coms.v(130[12] 305[6])
    defparam i13413_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i24901104_i1_3_lut (.I0(n62568), .I1(n62418), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n41));
    defparam i24901104_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13412_3_lut_4_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27118));   // verilog/coms.v(130[12] 305[6])
    defparam i13412_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n62709_bdd_4_lut (.I0(n62709), .I1(duty[1]), .I2(n269), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n62709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1976 (.I0(\data_out_frame[8] [7]), .I1(n23531), 
            .I2(n32_adj_5818), .I3(n23688), .O(n52842));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1976.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1977 (.I0(n52842), .I1(n22594), .I2(\data_out_frame[13] [4]), 
            .I3(n53069), .O(n10_adj_5845));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1977.LUT_INIT = 16'h6996;
    SB_LUT4 i46103_3_lut (.I0(n62658), .I1(n62532), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n61003));
    defparam i46103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1978 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53069));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1978.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1979 (.I0(\data_out_frame[6] [0]), .I1(n52496), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n52922));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1979.LUT_INIT = 16'h9696;
    SB_LUT4 i41767_3_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n56667));
    defparam i41767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41766_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[6] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n56666));
    defparam i41766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14239_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[18] [2]), 
            .O(n27945));   // verilog/coms.v(130[12] 305[6])
    defparam i14239_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i41768_4_lut (.I0(n56667), .I1(n25356), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n56668));
    defparam i41768_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i13411_3_lut_4_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27117));   // verilog/coms.v(130[12] 305[6])
    defparam i13411_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_1980 (.I0(\data_out_frame[8] [3]), .I1(n53161), 
            .I2(GND_net), .I3(GND_net), .O(n52584));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1980.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [5]), 
            .I2(n52584), .I3(\data_out_frame[10] [6]), .O(n12_adj_5719));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13410_3_lut_4_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27116));   // verilog/coms.v(130[12] 305[6])
    defparam i13410_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13409_3_lut_4_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27115));   // verilog/coms.v(130[12] 305[6])
    defparam i13409_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13408_3_lut_4_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27114));   // verilog/coms.v(130[12] 305[6])
    defparam i13408_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_3_lut_adj_1981 (.I0(\data_out_frame[13] [1]), .I1(n23945), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n53113));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1981.LUT_INIT = 16'h9696;
    SB_LUT4 i41773_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56673));
    defparam i41773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41774_4_lut (.I0(n56673), .I1(n25346), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n56674));
    defparam i41774_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i13407_3_lut_4_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27113));   // verilog/coms.v(130[12] 305[6])
    defparam i13407_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13406_3_lut_4_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27112));   // verilog/coms.v(130[12] 305[6])
    defparam i13406_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13405_3_lut_4_lut (.I0(deadband[19]), .I1(\data_in_frame[14] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27111));   // verilog/coms.v(130[12] 305[6])
    defparam i13405_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i41772_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56672));
    defparam i41772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13404_3_lut_4_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27110));   // verilog/coms.v(130[12] 305[6])
    defparam i13404_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i44735_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n59312));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i44735_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_4_lut_adj_1982 (.I0(commutation_state[0]), .I1(n4_adj_5846), 
            .I2(commutation_state_prev[0]), .I3(dti_N_380), .O(n24938));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_1982.LUT_INIT = 16'hdeff;
    SB_LUT4 i13507_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n54720), .I3(GND_net), .O(n27213));   // verilog/coms.v(130[12] 305[6])
    defparam i13507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13276_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n52427), .I3(GND_net), .O(n26982));   // verilog/coms.v(130[12] 305[6])
    defparam i13276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13273_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n52427), .I3(GND_net), .O(n26979));   // verilog/coms.v(130[12] 305[6])
    defparam i13273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1983 (.I0(n10_adj_5755), .I1(n3543), .I2(n35696), 
            .I3(GND_net), .O(n52409));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_adj_1983.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1984 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52641));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1984.LUT_INIT = 16'h6666;
    SB_LUT4 n9582_bdd_4_lut_47804 (.I0(n9582), .I1(n431), .I2(current[10]), 
            .I3(duty[23]), .O(n62763));
    defparam n9582_bdd_4_lut_47804.LUT_INIT = 16'he4aa;
    SB_LUT4 i13512_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n54720), .I3(GND_net), .O(n27218));   // verilog/coms.v(130[12] 305[6])
    defparam i13512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n62763_bdd_4_lut (.I0(n62763), .I1(duty[10]), .I2(n260), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[10]));
    defparam n62763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13266_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n52427), .I3(GND_net), .O(n26972));   // verilog/coms.v(130[12] 305[6])
    defparam i13266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13516_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[1]), .I2(n5_adj_5754), 
            .I3(n4_adj_5848), .O(n27222));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13516_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i38449_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n38306), 
            .I2(n10_adj_5755), .I3(GND_net), .O(n53298));
    defparam i38449_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13517_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[2]), .I2(n6_adj_5725), 
            .I3(n22880), .O(n27223));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13517_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_3_lut_adj_1985 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n52513));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1985.LUT_INIT = 16'h9696;
    SB_LUT4 i13518_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[3]), .I2(n6_adj_5725), 
            .I3(n22870), .O(n27224));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13518_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13263_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n52427), .I3(GND_net), .O(n26969));   // verilog/coms.v(130[12] 305[6])
    defparam i13263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13403_3_lut_4_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27109));   // verilog/coms.v(130[12] 305[6])
    defparam i13403_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13402_3_lut_4_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27108));   // verilog/coms.v(130[12] 305[6])
    defparam i13402_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_1986 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52928));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1986.LUT_INIT = 16'h6666;
    SB_LUT4 bit_ctr_0__bdd_4_lut_47664_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n62589));
    defparam bit_ctr_0__bdd_4_lut_47664_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i4_4_lut_adj_1987 (.I0(n52928), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(n53098), .O(n10_adj_5729));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1987.LUT_INIT = 16'h6996;
    SB_LUT4 i13520_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[4]), .I2(n5_adj_5809), 
            .I3(n22893), .O(n27226));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13520_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [1]), 
            .O(n52280));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i13398_3_lut_4_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27104));   // verilog/coms.v(130[12] 305[6])
    defparam i13398_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i24547_2_lut_2_lut (.I0(duty[20]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5037));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24547_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [2]), 
            .O(n52279));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i13521_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[5]), .I2(n5_adj_5754), 
            .I3(n22893), .O(n27227));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13521_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [5]), 
            .O(n52310));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [3]), 
            .O(n52278));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [6]), 
            .O(n52309));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.i [0]), .I1(n35706), 
            .I2(n38302), .I3(n10_adj_5778), .O(n25699));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1993.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [6]), 
            .O(n52308));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [7]), 
            .O(n52307));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47799 (.I0(n9582), .I1(n432), .I2(current[9]), 
            .I3(duty[23]), .O(n62757));
    defparam n9582_bdd_4_lut_47799.LUT_INIT = 16'he4aa;
    SB_LUT4 n62757_bdd_4_lut (.I0(n62757), .I1(duty[9]), .I2(n261), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n62757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [7]), 
            .O(n52306));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [0]), 
            .O(n26691));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [1]), 
            .O(n52154));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [2]), 
            .O(n52305));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i24548_2_lut_2_lut (.I0(duty[19]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5038));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24548_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [3]), 
            .O(n52304));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [4]), 
            .O(n52318));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [5]), 
            .O(n52303));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47794 (.I0(n9582), .I1(n433), .I2(current[8]), 
            .I3(duty[23]), .O(n62751));
    defparam n9582_bdd_4_lut_47794.LUT_INIT = 16'he4aa;
    SB_LUT4 n62751_bdd_4_lut (.I0(n62751), .I1(duty[8]), .I2(n262), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n62751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13522_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[6]), .I2(n6_adj_5753), 
            .I3(n22880), .O(n27228));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13522_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4192_4_lut (.I0(n22774), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5766));
    defparam i4192_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5766), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n54312));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [6]), 
            .O(n52158));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_2004 (.I0(n54312), .I1(delay_counter[18]), .I2(n22771), 
            .I3(GND_net), .O(n54562));
    defparam i2_3_lut_adj_2004.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_2005 (.I0(delay_counter[23]), .I1(n54562), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5722));
    defparam i2_4_lut_adj_2005.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_2006 (.I0(n7_adj_5722), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n22765), .O(n62));
    defparam i4_4_lut_adj_2006.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_2007 (.I0(delay_counter[24]), .I1(delay_counter[27]), 
            .I2(delay_counter[28]), .I3(delay_counter[29]), .O(n12_adj_5831));
    defparam i5_4_lut_adj_2007.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [4]), 
            .O(n52156));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [5]), 
            .O(n52277));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i6_4_lut_adj_2010 (.I0(delay_counter[26]), .I1(n12_adj_5831), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n22765));
    defparam i6_4_lut_adj_2010.LUT_INIT = 16'hfffe;
    SB_LUT4 i13356_3_lut_4_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27062));   // verilog/coms.v(130[12] 305[6])
    defparam i13356_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i5_3_lut_adj_2011 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_5853));
    defparam i5_3_lut_adj_2011.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_2012 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5852));
    defparam i6_4_lut_adj_2012.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_2013 (.I0(n15_adj_5852), .I1(delay_counter[2]), 
            .I2(n14_adj_5853), .I3(delay_counter[6]), .O(n22774));
    defparam i8_4_lut_adj_2013.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2014 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n22771));
    defparam i2_3_lut_adj_2014.LUT_INIT = 16'hfefe;
    SB_LUT4 i4184_3_lut (.I0(delay_counter[9]), .I1(delay_counter[10]), 
            .I2(n22774), .I3(GND_net), .O(n22));
    defparam i4184_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13355_3_lut_4_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27061));   // verilog/coms.v(130[12] 305[6])
    defparam i13355_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4183_4_lut (.I0(n22), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(n28));
    defparam i4183_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47565 (.I0(byte_transmit_counter[1]), 
            .I1(n56588), .I2(n56589), .I3(byte_transmit_counter[2]), .O(n62463));
    defparam byte_transmit_counter_1__bdd_4_lut_47565.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [6]), 
            .O(n52276));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 i13351_3_lut_4_lut (.I0(n1840), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3803), .O(n27057));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13351_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2016 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[10] [7]), 
            .O(n52275));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2016.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2017 (.I0(delay_counter[21]), .I1(delay_counter[20]), 
            .I2(delay_counter[23]), .I3(delay_counter[22]), .O(n4_adj_5781));
    defparam i1_4_lut_adj_2017.LUT_INIT = 16'h8000;
    SB_LUT4 i3166_4_lut (.I0(n28), .I1(delay_counter[19]), .I2(delay_counter[18]), 
            .I3(n4_adj_5840), .O(n40));
    defparam i3166_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i24347_4_lut (.I0(n40), .I1(delay_counter[31]), .I2(n22765), 
            .I3(n4_adj_5781), .O(n1365));   // verilog/TinyFPGA_B.v(382[14:38])
    defparam i24347_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i6_4_lut_adj_2018 (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5837));   // verilog/TinyFPGA_B.v(380[12:17])
    defparam i6_4_lut_adj_2018.LUT_INIT = 16'hfffe;
    SB_LUT4 i13350_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n27056));   // verilog/coms.v(130[12] 305[6])
    defparam i13350_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13349_3_lut_4_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27055));   // verilog/coms.v(130[12] 305[6])
    defparam i13349_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i5_4_lut_adj_2019 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5838));   // verilog/TinyFPGA_B.v(380[12:17])
    defparam i5_4_lut_adj_2019.LUT_INIT = 16'hfffe;
    SB_LUT4 i13348_3_lut_4_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27054));   // verilog/coms.v(130[12] 305[6])
    defparam i13348_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13347_3_lut_4_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27053));   // verilog/coms.v(130[12] 305[6])
    defparam i13347_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13346_3_lut_4_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27052));   // verilog/coms.v(130[12] 305[6])
    defparam i13346_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i24269_4_lut (.I0(n13_adj_5838), .I1(baudrate[0]), .I2(n14_adj_5837), 
            .I3(n22878), .O(n37857));
    defparam i24269_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2020 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [0]), 
            .O(n52274));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2020.LUT_INIT = 16'h2300;
    SB_LUT4 i13424_3_lut (.I0(\data_in_frame[16] [2]), .I1(rx_data[2]), 
            .I2(n25739), .I3(GND_net), .O(n27130));   // verilog/coms.v(130[12] 305[6])
    defparam i13424_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [1]), 
            .O(n52273));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47789 (.I0(n9582), .I1(n434), .I2(current[7]), 
            .I3(duty[23]), .O(n62745));
    defparam n9582_bdd_4_lut_47789.LUT_INIT = 16'he4aa;
    SB_LUT4 n62745_bdd_4_lut (.I0(n62745), .I1(duty[7]), .I2(n263), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n62745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9582_bdd_4_lut_47754 (.I0(n9582), .I1(n441), .I2(current[0]), 
            .I3(duty[23]), .O(n62703));
    defparam n9582_bdd_4_lut_47754.LUT_INIT = 16'he4aa;
    SB_LUT4 i14229_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[17] [0]), 
            .O(n27935));   // verilog/coms.v(130[12] 305[6])
    defparam i14229_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n62463_bdd_4_lut (.I0(n62463), .I1(n56826), .I2(n56825), .I3(byte_transmit_counter[2]), 
            .O(n62466));
    defparam n62463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [2]), 
            .O(n52272));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i13345_3_lut_4_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27051));   // verilog/coms.v(130[12] 305[6])
    defparam i13345_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13344_3_lut_4_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27050));   // verilog/coms.v(130[12] 305[6])
    defparam i13344_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13343_3_lut_4_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27049));   // verilog/coms.v(130[12] 305[6])
    defparam i13343_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13342_3_lut_4_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27048));   // verilog/coms.v(130[12] 305[6])
    defparam i13342_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13341_3_lut_4_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27047));   // verilog/coms.v(130[12] 305[6])
    defparam i13341_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13789_3_lut (.I0(ID[7]), .I1(data_adj_5912[7]), .I2(n25014), 
            .I3(GND_net), .O(n27495));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13790_3_lut (.I0(ID[6]), .I1(data_adj_5912[6]), .I2(n25014), 
            .I3(GND_net), .O(n27496));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44977_2_lut (.I0(n62586), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n59364));
    defparam i44977_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13791_3_lut (.I0(ID[5]), .I1(data_adj_5912[5]), .I2(n25014), 
            .I3(GND_net), .O(n27497));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24402_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_385));   // verilog/TinyFPGA_B.v(368[12:35])
    defparam i24402_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13340_3_lut_4_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27046));   // verilog/coms.v(130[12] 305[6])
    defparam i13340_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13792_3_lut (.I0(ID[4]), .I1(data_adj_5912[4]), .I2(n25014), 
            .I3(GND_net), .O(n27498));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12978_4_lut (.I0(n25013), .I1(n1365), .I2(n59196), .I3(n37969), 
            .O(n26655));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i12978_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5733));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13339_3_lut_4_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27045));   // verilog/coms.v(130[12] 305[6])
    defparam i13339_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2023 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [3]), 
            .O(n52271));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2023.LUT_INIT = 16'h2300;
    SB_LUT4 i45180_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n60080));
    defparam i45180_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5731));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [4]), 
            .O(n52270));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24571_2_lut (.I0(duty[5]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5052));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24571_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13338_3_lut_4_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27044));   // verilog/coms.v(130[12] 305[6])
    defparam i13338_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13337_3_lut_4_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27043));   // verilog/coms.v(130[12] 305[6])
    defparam i13337_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13336_3_lut_4_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27042));   // verilog/coms.v(130[12] 305[6])
    defparam i13336_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13793_3_lut (.I0(ID[3]), .I1(data_adj_5912[3]), .I2(n25014), 
            .I3(GND_net), .O(n27499));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13794_3_lut (.I0(ID[2]), .I1(data_adj_5912[2]), .I2(n25014), 
            .I3(GND_net), .O(n27500));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13795_3_lut (.I0(ID[1]), .I1(data_adj_5912[1]), .I2(n25014), 
            .I3(GND_net), .O(n27501));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13796_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3691 [23]), 
            .I2(control_update), .I3(GND_net), .O(n27502));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13335_3_lut_4_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27041));   // verilog/coms.v(130[12] 305[6])
    defparam i13335_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13334_3_lut_4_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27040));   // verilog/coms.v(130[12] 305[6])
    defparam i13334_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13333_3_lut_4_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27039));   // verilog/coms.v(130[12] 305[6])
    defparam i13333_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13524_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[7]), .I2(n6_adj_5753), 
            .I3(n22870), .O(n27230));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13332_3_lut_4_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27038));   // verilog/coms.v(130[12] 305[6])
    defparam i13332_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13525_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[8]), .I2(n5_adj_5809), 
            .I3(n22896), .O(n27231));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13525_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13526_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[9]), .I2(n5_adj_5754), 
            .I3(n22896), .O(n27232));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13526_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13797_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3691 [22]), 
            .I2(control_update), .I3(GND_net), .O(n27503));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13322_3_lut_4_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27028));   // verilog/coms.v(130[12] 305[6])
    defparam i13322_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13798_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3691 [21]), 
            .I2(control_update), .I3(GND_net), .O(n27504));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9582_bdd_4_lut_47784 (.I0(n9582), .I1(n435), .I2(current[6]), 
            .I3(duty[23]), .O(n62739));
    defparam n9582_bdd_4_lut_47784.LUT_INIT = 16'he4aa;
    SB_LUT4 i13527_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[10]), .I2(n6_adj_5752), 
            .I3(n22880), .O(n27233));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13527_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [5]), 
            .O(n52269));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h2300;
    SB_LUT4 i13799_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3691 [20]), 
            .I2(control_update), .I3(GND_net), .O(n27505));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [6]), 
            .O(n52268));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h2300;
    SB_LUT4 i13528_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[11]), .I2(n6_adj_5752), 
            .I3(n22870), .O(n27234));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13528_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13908_3_lut_4_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27614));   // verilog/coms.v(130[12] 305[6])
    defparam i13908_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n62739_bdd_4_lut (.I0(n62739), .I1(duty[6]), .I2(n264), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n62739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[11] [7]), 
            .O(n52267));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h2300;
    SB_LUT4 i13442_3_lut (.I0(\data_in_frame[16] [7]), .I1(rx_data[7]), 
            .I2(n25739), .I3(GND_net), .O(n27148));   // verilog/coms.v(130[12] 305[6])
    defparam i13442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13907_3_lut_4_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27613));   // verilog/coms.v(130[12] 305[6])
    defparam i13907_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13906_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27612));   // verilog/coms.v(130[12] 305[6])
    defparam i13906_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13254_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n52427), .I3(GND_net), .O(n26960));   // verilog/coms.v(130[12] 305[6])
    defparam i13254_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13800_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(\PID_CONTROLLER.integral_23__N_3691 [19]), 
            .I2(control_update), .I3(GND_net), .O(n27506));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5698));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13801_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(\PID_CONTROLLER.integral_23__N_3691 [18]), 
            .I2(control_update), .I3(GND_net), .O(n27507));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20330_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n33996), 
            .I2(control_update), .I3(GND_net), .O(n27508));   // verilog/motorControl.v(20[7:21])
    defparam i20330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5703));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13803_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3691 [16]), 
            .I2(control_update), .I3(GND_net), .O(n27509));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13804_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3691 [15]), 
            .I2(control_update), .I3(GND_net), .O(n27510));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13805_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3691 [14]), 
            .I2(control_update), .I3(GND_net), .O(n27511));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13806_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3691 [13]), 
            .I2(control_update), .I3(GND_net), .O(n27512));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13530_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[12]), .I2(n5_adj_5809), 
            .I3(n4_adj_5726), .O(n27236));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13530_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [0]), 
            .O(n52266));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47779 (.I0(n9582), .I1(n436), .I2(current[5]), 
            .I3(duty[23]), .O(n62733));
    defparam n9582_bdd_4_lut_47779.LUT_INIT = 16'he4aa;
    SB_LUT4 n62733_bdd_4_lut (.I0(n62733), .I1(duty[5]), .I2(n265), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n62733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [1]), 
            .O(n52265));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h2300;
    SB_LUT4 i13903_3_lut_4_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27609));   // verilog/coms.v(130[12] 305[6])
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [2]), 
            .O(n52264));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i13531_4_lut (.I0(CS_MISO_c), .I1(data_adj_5920[15]), .I2(n37991), 
            .I3(n22870), .O(n27237));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13531_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_adj_2031 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n52352));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_2031.LUT_INIT = 16'h2222;
    SB_LUT4 i12055_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n35706), 
            .I2(n52412), .I3(reset), .O(n25761));   // verilog/coms.v(158[12:15])
    defparam i12055_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [3]), 
            .O(n52263));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i13902_3_lut_4_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27608));   // verilog/coms.v(130[12] 305[6])
    defparam i13902_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13807_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3691 [12]), 
            .I2(control_update), .I3(GND_net), .O(n27513));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20035_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .I2(control_update), .I3(GND_net), .O(n27514));   // verilog/motorControl.v(20[7:21])
    defparam i20035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13809_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3691 [10]), 
            .I2(control_update), .I3(GND_net), .O(n27515));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13810_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3691 [9]), 
            .I2(control_update), .I3(GND_net), .O(n27516));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13811_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3691 [8]), 
            .I2(control_update), .I3(GND_net), .O(n27517));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13812_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3691 [7]), 
            .I2(control_update), .I3(GND_net), .O(n27518));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13317_3_lut_4_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27023));   // verilog/coms.v(130[12] 305[6])
    defparam i13317_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13813_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3691 [6]), 
            .I2(control_update), .I3(GND_net), .O(n27519));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13814_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3691 [5]), 
            .I2(control_update), .I3(GND_net), .O(n27520));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13815_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3691 [4]), 
            .I2(control_update), .I3(GND_net), .O(n27521));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13316_3_lut_4_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27022));   // verilog/coms.v(130[12] 305[6])
    defparam i13316_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[6] [7]), 
            .O(n52302));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h2300;
    SB_LUT4 i13816_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3691 [3]), 
            .I2(control_update), .I3(GND_net), .O(n27522));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47528 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n62427));
    defparam byte_transmit_counter_0__bdd_4_lut_47528.LUT_INIT = 16'he4aa;
    SB_LUT4 n62427_bdd_4_lut (.I0(n62427), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n62430));
    defparam n62427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n62703_bdd_4_lut (.I0(n62703), .I1(duty[0]), .I2(n270), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n62703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13315_3_lut_4_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27021));   // verilog/coms.v(130[12] 305[6])
    defparam i13315_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n62685_bdd_4_lut (.I0(n62685), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n62688));
    defparam n62685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13314_3_lut_4_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27020));   // verilog/coms.v(130[12] 305[6])
    defparam i13314_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2034 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [0]), 
            .O(n26705));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2034.LUT_INIT = 16'h2300;
    SB_LUT4 i13251_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n52427), .I3(GND_net), .O(n26957));   // verilog/coms.v(130[12] 305[6])
    defparam i13251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13313_3_lut_4_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27019));   // verilog/coms.v(130[12] 305[6])
    defparam i13313_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [0]), 
            .O(n52317));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h2300;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47523 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[2]), .O(n62415));
    defparam byte_transmit_counter_0__bdd_4_lut_47523.LUT_INIT = 16'he4aa;
    SB_LUT4 n62415_bdd_4_lut (.I0(n62415), .I1(\data_out_frame[11] [2]), 
            .I2(\data_out_frame[10] [2]), .I3(byte_transmit_counter[2]), 
            .O(n62418));
    defparam n62415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13817_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3691 [2]), 
            .I2(control_update), .I3(GND_net), .O(n27523));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13818_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3691 [1]), 
            .I2(control_update), .I3(GND_net), .O(n27524));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13312_3_lut_4_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27018));   // verilog/coms.v(130[12] 305[6])
    defparam i13312_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n9582_bdd_4_lut_47774 (.I0(n9582), .I1(n437), .I2(current[4]), 
            .I3(duty[23]), .O(n62727));
    defparam n9582_bdd_4_lut_47774.LUT_INIT = 16'he4aa;
    SB_LUT4 n62727_bdd_4_lut (.I0(n62727), .I1(duty[4]), .I2(n266), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n62727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13901_3_lut_4_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27607));   // verilog/coms.v(130[12] 305[6])
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [1]), 
            .O(n52316));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 i13_4_lut_adj_2037 (.I0(\data_in_frame[19] [5]), .I1(n53298), 
            .I2(n25734), .I3(rx_data[5]), .O(n51565));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2037.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13900_3_lut_4_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27606));   // verilog/coms.v(130[12] 305[6])
    defparam i13900_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13899_3_lut_4_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27605));   // verilog/coms.v(130[12] 305[6])
    defparam i13899_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13898_3_lut_4_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27604));   // verilog/coms.v(130[12] 305[6])
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [1]), 
            .O(n52315));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i13897_3_lut_4_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27603));   // verilog/coms.v(130[12] 305[6])
    defparam i13897_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13896_3_lut_4_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27602));   // verilog/coms.v(130[12] 305[6])
    defparam i13896_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 color_bit_N_478_1__bdd_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[5]), .I3(neopxl_color[7]), .O(n62637));
    defparam color_bit_N_478_1__bdd_4_lut_4_lut.LUT_INIT = 16'he6a2;
    SB_LUT4 i13895_3_lut_4_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27601));   // verilog/coms.v(130[12] 305[6])
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13894_3_lut_4_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27600));   // verilog/coms.v(130[12] 305[6])
    defparam i13894_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [2]), 
            .O(n52314));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h2300;
    SB_LUT4 i44860_4_lut (.I0(n7_adj_5718), .I1(n47509), .I2(n47529), 
            .I3(bit_ctr[0]), .O(n59353));   // verilog/neopixel.v(34[12] 116[6])
    defparam i44860_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i26_4_lut (.I0(n20312), .I1(n59353), .I2(state[1]), .I3(n4_adj_5814), 
            .O(n51153));   // verilog/neopixel.v(34[12] 116[6])
    defparam i26_4_lut.LUT_INIT = 16'hf5c5;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [3]), 
            .O(n52313));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h2300;
    SB_LUT4 i13893_3_lut_4_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27599));   // verilog/coms.v(130[12] 305[6])
    defparam i13893_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13892_3_lut_4_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27598));   // verilog/coms.v(130[12] 305[6])
    defparam i13892_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13311_3_lut_4_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27017));   // verilog/coms.v(130[12] 305[6])
    defparam i13311_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13310_3_lut_4_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27016));   // verilog/coms.v(130[12] 305[6])
    defparam i13310_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i41584_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56475));
    defparam i41584_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47446_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6543), .I2(n56475), 
            .I3(n25_adj_5851), .O(n17_adj_5850));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i47446_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i13891_3_lut_4_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27597));   // verilog/coms.v(130[12] 305[6])
    defparam i13891_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13889_3_lut_4_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27595));   // verilog/coms.v(130[12] 305[6])
    defparam i13889_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13888_3_lut_4_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27594));   // verilog/coms.v(130[12] 305[6])
    defparam i13888_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13887_3_lut_4_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27593));   // verilog/coms.v(130[12] 305[6])
    defparam i13887_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47744 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n62685));
    defparam byte_transmit_counter_0__bdd_4_lut_47744.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2041 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[1] [3]), 
            .O(n52312));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2041.LUT_INIT = 16'h2300;
    SB_LUT4 i20049_3_lut_4_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27015));
    defparam i20049_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [4]), 
            .O(n52311));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[5] [5]), 
            .O(n52157));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_4_lut_adj_2044 (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5723));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i2_3_lut_4_lut_adj_2044.LUT_INIT = 16'h2022;
    SB_LUT4 i1847_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1365), .I3(n37857), .O(n6543));   // verilog/TinyFPGA_B.v(364[5] 390[12])
    defparam i1847_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[0] [2]), 
            .O(n52218));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_2046 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1365), .I3(n37857), .O(n24_adj_5849));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_adj_2046.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[0] [3]), 
            .O(n52301));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2048 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [4]), 
            .O(n52262));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2048.LUT_INIT = 16'h2300;
    SB_LUT4 n9582_bdd_4_lut_47749 (.I0(n9582), .I1(n418), .I2(current[15]), 
            .I3(duty[23]), .O(n62403));
    defparam n9582_bdd_4_lut_47749.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2049 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [5]), 
            .O(n52261));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2049.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2050 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [6]), 
            .O(n52260));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2050.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[12] [7]), 
            .O(n52259));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 i13534_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n55734), 
            .I3(n27), .O(n27240));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13534_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2052 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [0]), 
            .O(n52258));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2052.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [1]), 
            .O(n52257));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2054 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [2]), 
            .O(n52256));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2054.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [3]), 
            .O(n52255));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h2300;
    coms neopxl_color_23__I_0 (.GND_net(GND_net), .\byte_transmit_counter[4] (byte_transmit_counter[4]), 
         .\byte_transmit_counter[0] (byte_transmit_counter[0]), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .\byte_transmit_counter[1] (byte_transmit_counter[1]), .\byte_transmit_counter[3] (byte_transmit_counter[3]), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .clk16MHz(clk16MHz), 
         .n2978(n2978), .\data_out_frame[10] ({\data_out_frame[10] }), .n52280(n52280), 
         .n52279(n52279), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n52310(n52310), .n52278(n52278), .tx_active(tx_active), .n26953(n26953), 
         .\data_in_frame[13] ({Open_3, Open_4, Open_5, Open_6, Open_7, 
         \data_in_frame[13] [2:0]}), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\FRAME_MATCHER.i_31__N_2485 (\FRAME_MATCHER.i_31__N_2485 ), .encoder0_position_scaled({encoder0_position_scaled}), 
         .n52309(n52309), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .n52308(n52308), .control_mode({control_mode}), .n3543(n3543), 
         .n52307(n52307), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n52306(n52306), .n26957(n26957), .n26691(n26691), .n52154(n52154), 
         .n52305(n52305), .n26960(n26960), .n52304(n52304), .n52318(n52318), 
         .n52303(n52303), .n52158(n52158), .n26969(n26969), .\data_in_frame[13][4] (\data_in_frame[13] [4]), 
         .n26972(n26972), .\data_in_frame[13][5] (\data_in_frame[13] [5]), 
         .n27218(n27218), .VCC_net(VCC_net), .\data_in_frame[18] ({Open_8, 
         Open_9, \data_in_frame[18] [5:0]}), .n26979(n26979), .\data_in_frame[13][6] (\data_in_frame[13] [6]), 
         .n26982(n26982), .\data_in_frame[13][7] (\data_in_frame[13] [7]), 
         .n27213(n27213), .\data_in_frame[14] ({\data_in_frame[14] }), .n27203(n27203), 
         .n27200(n27200), .encoder1_position_scaled({encoder1_position_scaled}), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .setpoint({setpoint}), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n52156(n52156), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n62658(n62658), .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .Kp_23__N_1724(Kp_23__N_1724), 
         .reset(reset), .n27192(n27192), .n52277(n52277), .n52276(n52276), 
         .n52275(n52275), .n52274(n52274), .n52273(n52273), .n52272(n52272), 
         .n52271(n52271), .n52270(n52270), .n52269(n52269), .n52268(n52268), 
         .n52267(n52267), .n52266(n52266), .n52265(n52265), .n52264(n52264), 
         .rx_data_ready(rx_data_ready), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .\FRAME_MATCHER.i[1] (\FRAME_MATCHER.i [1]), .\FRAME_MATCHER.i[2] (\FRAME_MATCHER.i [2]), 
         .n35706(n35706), .n27101(n27101), .\data_in_frame[16] ({\data_in_frame[16] [7:6], 
         Open_10, Open_11, \data_in_frame[16] [3:0]}), .n27105(n27105), 
         .\data_in_frame[2] ({Open_12, Open_13, \data_in_frame[2] [5:0]}), 
         .\Kp[5] (Kp[5]), .n30905(n30905), .n27148(n27148), .n27130(n27130), 
         .ID({ID}), .\data_in_frame[0][7] (\data_in_frame[0] [7]), .n27144(n27144), 
         .n27133(n27133), .n52263(n52263), .n27136(n27136), .\data_in_frame[16][4] (\data_in_frame[16] [4]), 
         .n27129(n27129), .deadband({deadband}), .n27128(n27128), .n27127(n27127), 
         .n27126(n27126), .n26731(n26731), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n26734(n26734), .n26737(n26737), .n26740(n26740), .n51817(n51817), 
         .n27772(n27772), .\data_in_frame[4] ({\data_in_frame[4] }), .n27124(n27124), 
         .n27123(n27123), .n27122(n27122), .n27121(n27121), .n27120(n27120), 
         .n26743(n26743), .n51681(n51681), .n51677(n51677), .n27312(n27312), 
         .n27317(n27317), .n51673(n51673), .n27321(n27321), .n26746(n26746), 
         .n26749(n26749), .n27327(n27327), .\data_in_frame[2][7] (\data_in_frame[2] [7]), 
         .n27331(n27331), .\data_in_frame[3][0] (\data_in_frame[3] [0]), 
         .n27757(n27757), .\data_in_frame[6][1] (\data_in_frame[6] [1]), 
         .n51669(n51669), .\data_in_frame[3][1] (\data_in_frame[3] [1]), 
         .n51667(n51667), .\data_in_frame[3][2] (\data_in_frame[3] [2]), 
         .n51663(n51663), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .n51659(n51659), .\data_in_frame[3][4] (\data_in_frame[3] [4]), 
         .n27119(n27119), .n27118(n27118), .n27117(n27117), .n27116(n27116), 
         .n27115(n27115), .n27114(n27114), .n27113(n27113), .n27112(n27112), 
         .n27111(n27111), .n27110(n27110), .n51655(n51655), .\data_in_frame[3][7] (\data_in_frame[3] [7]), 
         .n27365(n27365), .n27370(n27370), .n27375(n27375), .n27379(n27379), 
         .n27387(n27387), .n27391(n27391), .n27430(n27430), .\data_in_frame[18][7] (\data_in_frame[18] [7]), 
         .n27433(n27433), .n51579(n51579), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .n27439(n27439), .n27109(n27109), .n27108(n27108), .n27104(n27104), 
         .n27100(n27100), .neopxl_color({neopxl_color}), .n27099(n27099), 
         .n27097(n27097), .n27096(n27096), .n27095(n27095), .n27094(n27094), 
         .n27093(n27093), .n27092(n27092), .n27091(n27091), .n27662(n27662), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .n27659(n27659), .n20140(n20140), 
         .n27090(n27090), .n27089(n27089), .n27088(n27088), .n27087(n27087), 
         .n27086(n27086), .n27085(n27085), .n27084(n27084), .n27083(n27083), 
         .n27082(n27082), .n27081(n27081), .n27080(n27080), .n27656(n27656), 
         .n27653(n27653), .n27650(n27650), .n27647(n27647), .n27644(n27644), 
         .n27079(n27079), .n27078(n27078), .n51577(n51577), .n51575(n51575), 
         .\data_in_frame[6][2] (\data_in_frame[6] [2]), .\data_in_frame[6][3] (\data_in_frame[6] [3]), 
         .n27637(n27637), .n27062(n27062), .IntegralLimit({IntegralLimit}), 
         .n27061(n27061), .n27056(n27056), .n27055(n27055), .n27054(n27054), 
         .n27053(n27053), .\Ki[15] (Ki[15]), .n27052(n27052), .current_limit({current_limit}), 
         .n27051(n27051), .\Ki[13] (Ki[13]), .n27050(n27050), .n27049(n27049), 
         .\Ki[11] (Ki[11]), .n27048(n27048), .\Ki[10] (Ki[10]), .n27047(n27047), 
         .\Ki[9] (Ki[9]), .n27046(n27046), .\Ki[8] (Ki[8]), .n27045(n27045), 
         .\Ki[7] (Ki[7]), .n27044(n27044), .\Ki[6] (Ki[6]), .n27043(n27043), 
         .\Ki[5] (Ki[5]), .n27042(n27042), .\Ki[4] (Ki[4]), .n27041(n27041), 
         .\Ki[3] (Ki[3]), .n27040(n27040), .\Ki[2] (Ki[2]), .n27039(n27039), 
         .n27038(n27038), .\Ki[1] (Ki[1]), .n27028(n27028), .\Kp[15] (Kp[15]), 
         .\Kp[14] (Kp[14]), .n27614(n27614), .PWMLimit({PWMLimit}), .n27613(n27613), 
         .n27612(n27612), .n27611(n27611), .n27609(n27609), .n27608(n27608), 
         .n27023(n27023), .\Kp[13] (Kp[13]), .n27022(n27022), .\Kp[12] (Kp[12]), 
         .n27021(n27021), .\Kp[11] (Kp[11]), .n27020(n27020), .\Kp[10] (Kp[10]), 
         .n27019(n27019), .n27018(n27018), .\Ki[14] (Ki[14]), .n27607(n27607), 
         .n27606(n27606), .n27605(n27605), .n27604(n27604), .n27603(n27603), 
         .n27602(n27602), .n27601(n27601), .n27600(n27600), .n27599(n27599), 
         .n27598(n27598), .n27017(n27017), .\Ki[12] (Ki[12]), .n27016(n27016), 
         .n27597(n27597), .n27595(n27595), .n27594(n27594), .n27593(n27593), 
         .n27590(n27590), .\data_in_frame[6][4] (\data_in_frame[6] [4]), 
         .n27015(n27015), .n27014(n27014), .n27010(n27010), .\data_in_frame[6][6] (\data_in_frame[6] [6]), 
         .n52302(n52302), .n26986(n26986), .n26985(n26985), .\data_in_frame[6][7] (\data_in_frame[6] [7]), 
         .n51567(n51567), .n51549(n51549), .n27551(n27551), .n26978(n26978), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n26977(n26977), .n26976(n26976), .n26705(n26705), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n52317(n52317), .n52316(n52316), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n52315(n52315), .n52314(n52314), .n52313(n52313), .n52312(n52312), 
         .n52311(n52311), .n52157(n52157), .n26975(n26975), .n26968(n26968), 
         .n26956(n26956), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n52218(n52218), .n52301(n52301), .n26946(n26946), .n26944(n26944), 
         .n26930(n26930), .\Kp[1] (Kp[1]), .n26929(n26929), .\Kp[2] (Kp[2]), 
         .n26925(n26925), .\Kp[3] (Kp[3]), .n26924(n26924), .\Kp[4] (Kp[4]), 
         .n26920(n26920), .n26916(n26916), .\Ki[0] (Ki[0]), .n26915(n26915), 
         .\Kp[0] (Kp[0]), .n52262(n52262), .\motor_state_23__N_67[13] (motor_state_23__N_67[13]), 
         .n15(n15_adj_5727), .n9(n9_adj_5843), .n52261(n52261), .n52260(n52260), 
         .n52259(n52259), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n52258(n52258), .n52257(n52257), .n52256(n52256), .n52255(n52255), 
         .n52254(n52254), .n52160(n52160), .n52253(n52253), .n52252(n52252), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n52251(n52251), 
         .n52250(n52250), .n52249(n52249), .n52248(n52248), .n26347(n26347), 
         .n52247(n52247), .n52246(n52246), .n52217(n52217), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n52245(n52245), .n52244(n52244), .n52243(n52243), .n52242(n52242), 
         .n27549(n27549), .\data_in_frame[8] ({Open_14, Open_15, Open_16, 
         Open_17, Open_18, \data_in_frame[8] [2:0]}), .\data_in_frame[8][4] (\data_in_frame[8] [4]), 
         .\data_in_frame[8][5] (\data_in_frame[8] [5]), .\data_in_frame[8][6] (\data_in_frame[8] [6]), 
         .\data_in_frame[8][7] (\data_in_frame[8] [7]), .n51565(n51565), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .n52409(n52409), .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), 
         .n62586(n62586), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n52430(n52430), .rx_data({rx_data}), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n62532(n62532), 
         .n52241(n52241), .n52240(n52240), .n52239(n52239), .n52223(n52223), 
         .n52238(n52238), .n52237(n52237), .n52236(n52236), .n52235(n52235), 
         .n52234(n52234), .n52233(n52233), .n52232(n52232), .n52231(n52231), 
         .n27935(n27935), .n26327(n26327), .n52230(n52230), .n52229(n52229), 
         .n52228(n52228), .n52227(n52227), .n52226(n52226), .n52225(n52225), 
         .n52155(n52155), .n26319(n26319), .n52220(n52220), .n59364(n59364), 
         .n62466(n62466), .n27945(n27945), .n26317(n26317), .n52221(n52221), 
         .n52222(n52222), .n52224(n52224), .n52159(n52159), .n52219(n52219), 
         .n52161(n52161), .n52162(n52162), .n52163(n52163), .n52164(n52164), 
         .n52165(n52165), .n52166(n52166), .n52167(n52167), .n52168(n52168), 
         .n52169(n52169), .n27960(n27960), .n26302(n26302), .n52170(n52170), 
         .n27962(n27962), .n26300(n26300), .n52171(n52171), .n52172(n52172), 
         .n52173(n52173), .n52174(n52174), .n52175(n52175), .n27968(n27968), 
         .n26294(n26294), .n52176(n52176), .n27970(n27970), .n26292(n26292), 
         .n52177(n52177), .n52178(n52178), .n52179(n52179), .n52180(n52180), 
         .n52181(n52181), .n52182(n52182), .n52183(n52183), .n27978(n27978), 
         .n26284(n26284), .n27979(n27979), .n26283(n26283), .n52184(n52184), 
         .n27981(n27981), .n26281(n26281), .n52185(n52185), .n52186(n52186), 
         .n52187(n52187), .n27985(n27985), .n26277(n26277), .n27986(n27986), 
         .n26276(n26276), .n54720(n54720), .n27987(n27987), .n26275(n26275), 
         .n52188(n52188), .n52189(n52189), .n52190(n52190), .n52191(n52191), 
         .n52192(n52192), .n52193(n52193), .n52194(n52194), .n52195(n52195), 
         .n52196(n52196), .n52197(n52197), .n52198(n52198), .n52199(n52199), 
         .n52200(n52200), .n52201(n52201), .n52202(n52202), .n52203(n52203), 
         .n52204(n52204), .n52205(n52205), .n52206(n52206), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n4(n4_adj_5750), .\data_in_frame[10] ({Open_19, \data_in_frame[10] [6], 
         Open_20, Open_21, Open_22, Open_23, Open_24, Open_25}), 
         .\data_out_frame[26][2] (\data_out_frame[26] [2]), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
         .\data_out_frame[27][2] (\data_out_frame[27] [2]), .n23375(n23375), 
         .Kp_23__N_645(Kp_23__N_645), .n52455(n52455), .\Kp[6] (Kp[6]), 
         .n52656(n52656), .n26787(n26787), .\Kp[7] (Kp[7]), .n26786(n26786), 
         .n25709(n25709), .n25766(n25766), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n52207(n52207), .n52208(n52208), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .n52209(n52209), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .n52210(n52210), .\data_out_frame[3][7] (\data_out_frame[3] [7]), 
         .n52211(n52211), .n52212(n52212), .n26782(n26782), .n28044(n28044), 
         .n26215(n26215), .n52213(n52213), .n28046(n28046), .n26213(n26213), 
         .n52214(n52214), .n52215(n52215), .n28052(n28052), .n26207(n26207), 
         .LED_c(LED_c), .n52216(n52216), .DE_c(DE_c), .n26769(n26769), 
         .\Kp[8] (Kp[8]), .n26768(n26768), .\Kp[9] (Kp[9]), .n52300(n52300), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n52299(n52299), 
         .n52298(n52298), .n52297(n52297), .n52296(n52296), .n52295(n52295), 
         .n28093(n28093), .n26402(n26402), .n52294(n52294), .n28095(n28095), 
         .n26400(n26400), .n28096(n28096), .n26399(n26399), .n52293(n52293), 
         .n52292(n52292), .n52291(n52291), .n52290(n52290), .n52289(n52289), 
         .n52288(n52288), .n52287(n52287), .n26391(n26391), .n28105(n28105), 
         .n26390(n26390), .n52286(n52286), .\data_in_frame[10][0] (\data_in_frame[10] [0]), 
         .\data_in_frame[10][1] (\data_in_frame[10] [1]), .\data_in_frame[10][2] (\data_in_frame[10] [2]), 
         .\data_in_frame[10][3] (\data_in_frame[10] [3]), .\data_in_frame[10][4] (\data_in_frame[10] [4]), 
         .n51563(n51563), .n51585(n51585), .n51561(n51561), .n51559(n51559), 
         .n51557(n51557), .n51555(n51555), .n51553(n51553), .n51551(n51551), 
         .n52285(n52285), .n52284(n52284), .n52283(n52283), .n52282(n52282), 
         .n28111(n28111), .n26384(n26384), .n22568(n22568), .n23824(n23824), 
         .n53055(n53055), .n52281(n52281), .n10(n10), .n38306(n38306), 
         .n25768(n25768), .n47452(n47452), .n52831(n52831), .n52848(n52848), 
         .n23338(n23338), .n47989(n47989), .n16(n16_adj_5847), .n53140(n53140), 
         .n52878(n52878), .Kp_23__N_969(Kp_23__N_969), .Kp_23__N_675(Kp_23__N_675), 
         .n3(n3_adj_5751), .n375(n375), .n11(n11_adj_5813), .n53137(n53137), 
         .n11_adj_8(n11_adj_5812), .n52925(n52925), .n13(n13_adj_5817), 
         .n52424(n52424), .n38302(n38302), .n52412(n52412), .n10_adj_9(n10_adj_5755), 
         .n25739(n25739), .n23958(n23958), .n1513(n1513), .n52564(n52564), 
         .n35696(n35696), .n53098(n53098), .n25705(n25705), .n52842(n52842), 
         .n47380(n47380), .n23427(n23427), .n53035(n53035), .n25707(n25707), 
         .n23531(n23531), .n22594(n22594), .n23688(n23688), .n1130(n1130), 
         .n23945(n23945), .n32(n32_adj_5818), .n53161(n53161), .n56674(n56674), 
         .n56672(n56672), .n52053(n52053), .n151(n151), .n203(n203), 
         .n181(n181), .n155(n155), .\PID_CONTROLLER.integral_23__N_3691[3] (\PID_CONTROLLER.integral_23__N_3691 [3]), 
         .\current[11] (current[11]), .\data[11] (data_adj_5920[11]), .n25021(n25021), 
         .n27452(n27452), .displacement({displacement}), .n15_adj_10(n15_adj_5724), 
         .n15_adj_11(n15_adj_5728), .\motor_state_23__N_67[17] (motor_state_23__N_67[17]), 
         .n2076(n2076), .n52979(n52979), .n52928(n52928), .n23594(n23594), 
         .n53122(n53122), .n68(n68), .n62598(n62598), .n59386(n59386), 
         .n25356(n25356), .n52922(n52922), .n52641(n52641), .n56668(n56668), 
         .n56666(n56666), .n53069(n53069), .n52513(n52513), .n12(n12_adj_5719), 
         .n8(n8_adj_5720), .n52434(n52434), .n25346(n25346), .n52939(n52939), 
         .n52741(n52741), .n25699(n25699), .n204(n204), .n6(n6_adj_5811), 
         .n152(n152), .n60212(n60212), .n53113(n53113), .n53125(n53125), 
         .n52496(n52496), .n25734(n25734), .n10_adj_12(n10_adj_5778), 
         .n25750(n25750), .n35727(n35727), .\current[7] (current[7]), 
         .\current[6] (current[6]), .\current[5] (current[5]), .\current[4] (current[4]), 
         .\current[3] (current[3]), .\current[2] (current[2]), .\current[1] (current[1]), 
         .\current[0] (current[0]), .\current[15] (current[15]), .\current[10] (current[10]), 
         .\current[9] (current[9]), .\current[8] (current[8]), .n62688(n62688), 
         .n62430(n62430), .pwm_setpoint({pwm_setpoint}), .n52427(n52427), 
         .n62840(n62840), .r_SM_Main({r_SM_Main_adj_5933}), .r_Clock_Count({r_Clock_Count_adj_5934}), 
         .tx_o(tx_o), .n26943(n26943), .\tx_data[2] (tx_data[2]), .n23(n23_adj_5854), 
         .\o_Rx_DV_N_3464[12] (o_Rx_DV_N_3464[12]), .n4858(n4858), .\o_Rx_DV_N_3464[24] (o_Rx_DV_N_3464[24]), 
         .n27(n27), .n29(n29), .n6_adj_13(n6_adj_5842), .tx_enable(tx_enable), 
         .n27247(n27247), .baudrate({baudrate}), .n55830(n55830), .n27246(n27246), 
         .n27245(n27245), .n27243(n27243), .n27242(n27242), .\o_Rx_DV_N_3464[8] (o_Rx_DV_N_3464[8]), 
         .n4855(n4855), .n52352(n52352), .\r_SM_Main[1]_adj_14 (r_SM_Main[1]), 
         .n25039(n25039), .n27241(n27241), .n27240(n27240), .\r_SM_Main[2]_adj_15 (r_SM_Main[2]), 
         .n55782(n55782), .r_Clock_Count_adj_24({r_Clock_Count}), .n55798(n55798), 
         .n55750(n55750), .n55766(n55766), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
         .n22878(n22878), .\o_Rx_DV_N_3464[7] (o_Rx_DV_N_3464[7]), .\o_Rx_DV_N_3464[6] (o_Rx_DV_N_3464[6]), 
         .\o_Rx_DV_N_3464[5] (o_Rx_DV_N_3464[5]), .\o_Rx_DV_N_3464[4] (o_Rx_DV_N_3464[4]), 
         .\o_Rx_DV_N_3464[3] (o_Rx_DV_N_3464[3]), .\o_Rx_DV_N_3464[2] (o_Rx_DV_N_3464[2]), 
         .\o_Rx_DV_N_3464[1] (o_Rx_DV_N_3464[1]), .\o_Rx_DV_N_3464[0] (o_Rx_DV_N_3464[0]), 
         .n25264(n25264), .n27583(n27583), .n48661(n48661), .n27579(n27579), 
         .\r_Bit_Index[0] (r_Bit_Index[0]), .n53350(n53350), .n55734(n55734), 
         .n55846(n55846), .n55814(n55814)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [4]), 
            .O(n52254));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h2300;
    SB_LUT4 n62403_bdd_3_lut (.I0(n62403), .I1(duty[23]), .I2(n249), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam n62403_bdd_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 i13535_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n55846), 
            .I3(n27), .O(n27241));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13535_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [5]), 
            .O(n52160));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    \quadrature_decoder(1)_U0  quad_counter0 (.\a_new[1] (a_new[1]), .b_prev(b_prev), 
            .GND_net(GND_net), .ENCODER0_B_N_keep(ENCODER0_B_N), .n1884(clk16MHz), 
            .ENCODER0_A_N_keep(ENCODER0_A_N), .n1842(n1842), .n1844(n1844), 
            .n1846(n1846), .n1848(n1848), .n1850(n1850), .n1852(n1852), 
            .n1854(n1854), .n1856(n1856), .\encoder0_position[23] (encoder0_position[23]), 
            .\encoder0_position[22] (encoder0_position[22]), .\encoder0_position[21] (encoder0_position[21]), 
            .\encoder0_position[20] (encoder0_position[20]), .\encoder0_position[19] (encoder0_position[19]), 
            .position_31__N_3803(position_31__N_3803), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .n27057(n27057), 
            .n1840(n1840), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[49] 310[6])
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n25039), .O(n48661));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [6]), 
            .O(n52253));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h2300;
    SB_LUT4 i13216_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3691 [0]), 
            .I2(control_update), .I3(GND_net), .O(n26922));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9582_bdd_4_lut_47769 (.I0(n9582), .I1(n438), .I2(current[3]), 
            .I3(duty[23]), .O(n62721));
    defparam n9582_bdd_4_lut_47769.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[13] [7]), 
            .O(n52252));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h2300;
    SB_LUT4 i13308_3_lut_4_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27014));   // verilog/coms.v(130[12] 305[6])
    defparam i13308_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13304_3_lut_4_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27010));   // verilog/coms.v(130[12] 305[6])
    defparam i13304_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13217_3_lut (.I0(ID[0]), .I1(data_adj_5912[0]), .I2(n25014), 
            .I3(GND_net), .O(n26923));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13536_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n55814), 
            .I3(n27), .O(n27242));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13536_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_4_lut_adj_2060 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_385), .I3(n2925), .O(n25_adj_5851));   // verilog/TinyFPGA_B.v(379[7:11])
    defparam i1_4_lut_4_lut_adj_2060.LUT_INIT = 16'h5450;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [0]), 
            .O(n52251));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h2300;
    SB_LUT4 i13226_3_lut (.I0(current[0]), .I1(data_adj_5920[0]), .I2(n25021), 
            .I3(GND_net), .O(n26932));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24549_2_lut_2_lut (.I0(duty[18]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5039));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24549_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13228_3_lut (.I0(CS_c), .I1(state_adj_5922[0]), .I2(state_adj_5922[1]), 
            .I3(GND_net), .O(n26934));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13228_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i47493_4_lut (.I0(n15_adj_5756), .I1(clk_out), .I2(state_adj_5922[0]), 
            .I3(state_adj_5922[1]), .O(n9_adj_5855));   // verilog/tli4970.v(35[10] 68[6])
    defparam i47493_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i24550_2_lut_2_lut (.I0(duty[17]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5040));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24550_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 n62721_bdd_4_lut (.I0(n62721), .I1(duty[3]), .I2(n267), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n62721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13303_3_lut_4_lut (.I0(n1889), .I1(b_prev_adj_5759), .I2(a_new_adj_5900[1]), 
            .I3(position_31__N_3803_adj_5760), .O(n27009));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13303_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i10_1_lut_adj_2062 (.I0(duty[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_setpoint_23__N_183));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut_adj_2062.LUT_INIT = 16'h5555;
    SB_LUT4 i24551_2_lut_2_lut (.I0(duty[16]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5041));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24551_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [1]), 
            .O(n52250));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i14405_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [7]), 
            .O(n28111));   // verilog/coms.v(130[12] 305[6])
    defparam i14405_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14399_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[9] [1]), 
            .O(n28105));   // verilog/coms.v(130[12] 305[6])
    defparam i14399_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2064 (.I0(hall1), .I1(commutation_state[2]), .I2(hall3), 
            .I3(hall2), .O(n51937));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_2064.LUT_INIT = 16'hd054;
    SB_LUT4 i14390_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[8] [0]), 
            .O(n28096));   // verilog/coms.v(130[12] 305[6])
    defparam i14390_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14389_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [7]), 
            .O(n28095));   // verilog/coms.v(130[12] 305[6])
    defparam i14389_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13280_3_lut_4_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26986));   // verilog/coms.v(130[12] 305[6])
    defparam i13280_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i14387_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[7] [5]), 
            .O(n28093));   // verilog/coms.v(130[12] 305[6])
    defparam i14387_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14346_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [6]), 
            .O(n28052));   // verilog/coms.v(130[12] 305[6])
    defparam i14346_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5697));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13279_3_lut_4_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26985));   // verilog/coms.v(130[12] 305[6])
    defparam i13279_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [2]), 
            .O(n52249));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 i14340_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [3]), 
            .O(n28046));   // verilog/coms.v(130[12] 305[6])
    defparam i14340_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [3]), 
            .O(n52248));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2067 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [4]), 
            .O(n26347));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2067.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_adj_2068 (.I0(rx_data[7]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n38306), .I3(GND_net), .O(n52362));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_2068.LUT_INIT = 16'h8080;
    SB_LUT4 i13272_3_lut_4_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26978));   // verilog/coms.v(130[12] 305[6])
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [5]), 
            .O(n52247));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2070 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [6]), 
            .O(n52246));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2070.LUT_INIT = 16'h2300;
    SB_LUT4 i14338_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[4] [1]), 
            .O(n28044));   // verilog/coms.v(130[12] 305[6])
    defparam i14338_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24552_2_lut_2_lut (.I0(duty[15]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5042));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i24552_2_lut_2_lut.LUT_INIT = 16'h4444;
    TLI4970 tli (.clk_out(clk_out), .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), 
            .GND_net(GND_net), .n27237(n27237), .\data[15] (data_adj_5920[15]), 
            .n27236(n27236), .\data[12] (data_adj_5920[12]), .n27234(n27234), 
            .\data[11] (data_adj_5920[11]), .n27233(n27233), .\data[10] (data_adj_5920[10]), 
            .n27232(n27232), .\data[9] (data_adj_5920[9]), .n27231(n27231), 
            .\data[8] (data_adj_5920[8]), .n27230(n27230), .\data[7] (data_adj_5920[7]), 
            .n27228(n27228), .\data[6] (data_adj_5920[6]), .n27227(n27227), 
            .\data[5] (data_adj_5920[5]), .n27226(n27226), .\data[4] (data_adj_5920[4]), 
            .n27224(n27224), .\data[3] (data_adj_5920[3]), .n27223(n27223), 
            .\data[2] (data_adj_5920[2]), .n27222(n27222), .\data[1] (data_adj_5920[1]), 
            .clk16MHz(clk16MHz), .\state[1] (state_adj_5922[1]), .\state[0] (state_adj_5922[0]), 
            .n27584(n27584), .\data[0] (data_adj_5920[0]), .n9(n9_adj_5855), 
            .n26934(n26934), .n26932(n26932), .\current[0] (current[0]), 
            .n25021(n25021), .\current[15] (current[15]), .n27462(n27462), 
            .\current[1] (current[1]), .n27461(n27461), .\current[2] (current[2]), 
            .n27460(n27460), .\current[3] (current[3]), .n27459(n27459), 
            .\current[4] (current[4]), .n27458(n27458), .\current[5] (current[5]), 
            .n27457(n27457), .\current[6] (current[6]), .n27456(n27456), 
            .\current[7] (current[7]), .n27455(n27455), .\current[8] (current[8]), 
            .n27454(n27454), .\current[9] (current[9]), .n27453(n27453), 
            .\current[10] (current[10]), .n27452(n27452), .\current[11] (current[11]), 
            .VCC_net(VCC_net), .n15(n15_adj_5756), .n4(n4_adj_5726), .n22896(n22896), 
            .n22893(n22893), .n4_adj_3(n4_adj_5848), .n22870(n22870), 
            .n22880(n22880), .state_7__N_4293(state_7__N_4293), .n6(n6_adj_5725), 
            .n6_adj_4(n6_adj_5753), .n5(n5_adj_5754), .n6_adj_5(n6_adj_5752), 
            .n5_adj_6(n5_adj_5809), .n37991(n37991), .n11(n11_adj_5757)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(407[11] 413[4])
    EEPROM eeprom (.GND_net(GND_net), .clk16MHz(clk16MHz), .\state_7__N_3892[0] (state_7__N_3892[0]), 
           .enable_slow_N_4187(enable_slow_N_4187), .data_ready(data_ready), 
           .n26923(n26923), .ID({ID}), .n27501(n27501), .n27500(n27500), 
           .n27499(n27499), .n27498(n27498), .n27497(n27497), .n27496(n27496), 
           .n27495(n27495), .baudrate({baudrate}), .n27486(n27486), .n27485(n27485), 
           .n27484(n27484), .n27483(n27483), .n27482(n27482), .n27470(n27470), 
           .n27469(n27469), .n27468(n27468), .n27467(n27467), .n27466(n27466), 
           .n27465(n27465), .n27464(n27464), .n27463(n27463), .n25014(n25014), 
           .n25295(n25295), .n25293(n25293), .\state[0] (state_adj_5946[0]), 
           .data({data_adj_5912}), .\state_7__N_4084[0] (state_7__N_4084[0]), 
           .n27252(n27252), .n27251(n27251), .sda_enable(sda_enable), 
           .sda_out(sda_out), .\counter[0] (counter_adj_5947[0]), .n37902(n37902), 
           .n6352(n6352), .scl_enable(scl_enable), .VCC_net(VCC_net), 
           .n27572(n27572), .n8(n8_adj_5856), .n27259(n27259), .n27257(n27257), 
           .n27256(n27256), .n27255(n27255), .n27253(n27253), .n22915(n22915), 
           .scl(scl), .\state_7__N_4100[3] (state_7__N_4100[3]), .n22875(n22875), 
           .n6(n6_adj_5721), .n22907(n22907), .n22918(n22918)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(393[10] 405[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2071 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[14] [7]), 
            .O(n52217));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2071.LUT_INIT = 16'h2300;
    SB_LUT4 i14281_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [4]), 
            .O(n27987));   // verilog/coms.v(130[12] 305[6])
    defparam i14281_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20343_3_lut_4_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26977));
    defparam i20343_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    motorControl control (.\Kp[3] (Kp[3]), .GND_net(GND_net), .\Ki[15] (Ki[15]), 
            .\PID_CONTROLLER.integral_23__N_3691[7] (\PID_CONTROLLER.integral_23__N_3691 [7]), 
            .\Kp[5] (Kp[5]), .\Kp[4] (Kp[4]), .PWMLimit({PWMLimit}), .\Kp[0] (Kp[0]), 
            .\Kp[1] (Kp[1]), .control_update(control_update), .duty({duty}), 
            .clk16MHz(clk16MHz), .reset(reset), .setpoint({setpoint}), 
            .\motor_state[18] (motor_state[18]), .n35(n35), .\Kp[6] (Kp[6]), 
            .n181(n181), .IntegralLimit({IntegralLimit}), .n155(n155), 
            .\Ki[6] (Ki[6]), .\PID_CONTROLLER.integral_23__N_3691[12] (\PID_CONTROLLER.integral_23__N_3691 [12]), 
            .\Ki[1] (Ki[1]), .\PID_CONTROLLER.integral_23__N_3691[6] (\PID_CONTROLLER.integral_23__N_3691 [6]), 
            .\Ki[0] (Ki[0]), .\Kp[2] (Kp[2]), .\Ki[7] (Ki[7]), .\Kp[12] (Kp[12]), 
            .\Kp[7] (Kp[7]), .\Ki[2] (Ki[2]), .n11(n11_adj_5812), .\Ki[3] (Ki[3]), 
            .\Ki[8] (Ki[8]), .\Kp[13] (Kp[13]), .\Ki[14] (Ki[14]), .\PID_CONTROLLER.integral_23__N_3691[15] (\PID_CONTROLLER.integral_23__N_3691 [15]), 
            .\PID_CONTROLLER.integral_23__N_3691[14] (\PID_CONTROLLER.integral_23__N_3691 [14]), 
            .n375(n375), .\PID_CONTROLLER.integral_23__N_3691[3] (\PID_CONTROLLER.integral_23__N_3691 [3]), 
            .\Ki[9] (Ki[9]), .\Ki[4] (Ki[4]), .n214(n214), .\PID_CONTROLLER.integral_23__N_3691[16] (\PID_CONTROLLER.integral_23__N_3691 [16]), 
            .\PID_CONTROLLER.integral_23__N_3691[4] (\PID_CONTROLLER.integral_23__N_3691 [4]), 
            .\Kp[8] (Kp[8]), .\PID_CONTROLLER.integral_23__N_3691[0] (\PID_CONTROLLER.integral_23__N_3691 [0]), 
            .\Ki[12] (Ki[12]), .\Kp[14] (Kp[14]), .\Ki[5] (Ki[5]), .\Kp[15] (Kp[15]), 
            .deadband({deadband}), .\motor_state[17] (motor_state[17]), 
            .\PID_CONTROLLER.integral_23__N_3691[11] (\PID_CONTROLLER.integral_23__N_3691 [11]), 
            .\Ki[10] (Ki[10]), .n5(n5_adj_5839), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .n9(n9_adj_5843), .\Ki[11] (Ki[11]), 
            .\motor_state[12] (motor_state[12]), .n545(n545), .n143(n143), 
            .n220(n220), .\motor_state[11] (motor_state[11]), .\motor_state[10] (motor_state[10]), 
            .VCC_net(VCC_net), .n472(n472), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .\PID_CONTROLLER.integral_23__N_3691[10] (\PID_CONTROLLER.integral_23__N_3691 [10]), 
            .n399(n399), .n326(n326), .n253(n253_adj_5833), .n180(n180), 
            .\motor_state[7] (motor_state[7]), .n53(n53_adj_5836), .\motor_state[6] (motor_state[6]), 
            .n107(n107), .\motor_state[5] (motor_state[5]), .n203(n203), 
            .\motor_state[4] (motor_state[4]), .n204(n204), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .\Kp[11] (Kp[11]), .\motor_state[1] (motor_state[1]), 
            .\Kp[9] (Kp[9]), .\motor_state[0] (motor_state[0]), .\PID_CONTROLLER.integral_23__N_3691[1] (\PID_CONTROLLER.integral_23__N_3691 [1]), 
            .\Kp[10] (Kp[10]), .\PID_CONTROLLER.integral_23__N_3691[13] (\PID_CONTROLLER.integral_23__N_3691 [13]), 
            .\Ki[13] (Ki[13]), .n26922(n26922), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .n27524(n27524), .n27523(n27523), .n27522(n27522), .n27521(n27521), 
            .n27520(n27520), .n27519(n27519), .n27518(n27518), .n27517(n27517), 
            .n27516(n27516), .n27515(n27515), .n27514(n27514), .n27513(n27513), 
            .n27512(n27512), .n27511(n27511), .n27510(n27510), .n27509(n27509), 
            .n27508(n27508), .n27507(n27507), .n27506(n27506), .n27505(n27505), 
            .n27504(n27504), .n27503(n27503), .n27502(n27502), .n23(n23_adj_5810), 
            .n53137(n53137), .\data_in_frame[9][6] (\data_in_frame[9] [6]), 
            .\data_in_frame[11][3] (\data_in_frame[11] [3]), .Kp_23__N_969(Kp_23__N_969), 
            .n53140(n53140), .Kp_23__N_645(Kp_23__N_645), .\data_in_frame[11][4] (\data_in_frame[11] [4]), 
            .\data_in_frame[12][3] (\data_in_frame[12] [3]), .n23958(n23958), 
            .\data_in_frame[12][5] (\data_in_frame[12] [5]), .n23338(n23338), 
            .\data_in_frame[12][1] (\data_in_frame[12] [1]), .Kp_23__N_675(Kp_23__N_675), 
            .n52656(n52656), .n52455(n52455), .n52831(n52831), .n52848(n52848), 
            .n52925(n52925), .n22568(n22568), .n151(n151), .n152(n152), 
            .n490(n490), .n417(n417), .n344(n344_adj_5832), .n271(n271), 
            .n198(n198), .n125(n125), .\motor_state[23] (motor_state[23]), 
            .n9_adj_1(n9_adj_5816), .\motor_state[21] (motor_state[21]), 
            .\PID_CONTROLLER.integral_23__N_3691[23] (\PID_CONTROLLER.integral_23__N_3691 [23]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .n60212(n60212), .n6(n6_adj_5811), .\PID_CONTROLLER.integral_23__N_3691[2] (\PID_CONTROLLER.integral_23__N_3691 [2]), 
            .\PID_CONTROLLER.integral_23__N_3691[5] (\PID_CONTROLLER.integral_23__N_3691 [5]), 
            .\PID_CONTROLLER.integral_23__N_3691[9] (\PID_CONTROLLER.integral_23__N_3691 [9]), 
            .\PID_CONTROLLER.integral_23__N_3691[8] (\PID_CONTROLLER.integral_23__N_3691 [8]), 
            .\PID_CONTROLLER.integral_23__N_3691[18] (\PID_CONTROLLER.integral_23__N_3691 [18]), 
            .\PID_CONTROLLER.integral_23__N_3691[20] (\PID_CONTROLLER.integral_23__N_3691 [20]), 
            .\PID_CONTROLLER.integral_23__N_3691[22] (\PID_CONTROLLER.integral_23__N_3691 [22]), 
            .\PID_CONTROLLER.integral_23__N_3691[19] (\PID_CONTROLLER.integral_23__N_3691 [19]), 
            .\PID_CONTROLLER.integral_23__N_3691[21] (\PID_CONTROLLER.integral_23__N_3691 [21]), 
            .n11_adj_2(n11_adj_5813), .n4(n4_adj_5750), .n3(n3_adj_5751), 
            .\data_in_frame[10][4] (\data_in_frame[10] [4]), .n23375(n23375), 
            .n23824(n23824), .n53055(n53055), .n47989(n47989), .\data_in_frame[9][5] (\data_in_frame[9] [5]), 
            .\data_in_frame[11][6] (\data_in_frame[11] [6]), .n47452(n47452), 
            .n16(n16_adj_5847), .n52878(n52878), .Kp_23__N_1724(Kp_23__N_1724), 
            .n30905(n30905), .n27611(n27611)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    SB_LUT4 i14280_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [3]), 
            .O(n27986));   // verilog/coms.v(130[12] 305[6])
    defparam i14280_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14279_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[23] [2]), 
            .O(n27985));   // verilog/coms.v(130[12] 305[6])
    defparam i14279_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9582_bdd_4_lut_47764 (.I0(n9582), .I1(n439), .I2(current[2]), 
            .I3(duty[23]), .O(n62715));
    defparam n9582_bdd_4_lut_47764.LUT_INIT = 16'he4aa;
    SB_LUT4 i24257_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i24257_2_lut.LUT_INIT = 16'h8888;
    \quadrature_decoder(1)  quad_counter1 (.b_prev(b_prev_adj_5759), .GND_net(GND_net), 
            .a_new({a_new_adj_5900[1], Open_26}), .position_31__N_3803(position_31__N_3803_adj_5760), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1884(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .n27009(n27009), .n1889(n1889), .\encoder1_position[0] (encoder1_position[0]), 
            .\encoder1_position[1] (encoder1_position[1]), .\encoder1_position[2] (encoder1_position[2]), 
            .\encoder1_position[3] (encoder1_position[3]), .\encoder1_position[4] (encoder1_position[4]), 
            .\encoder1_position[5] (encoder1_position[5]), .\encoder1_position[6] (encoder1_position[6]), 
            .\encoder1_position[7] (encoder1_position[7]), .\encoder1_position[8] (encoder1_position[8]), 
            .\encoder1_position[9] (encoder1_position[9]), .\encoder1_position[10] (encoder1_position[10]), 
            .\encoder1_position[11] (encoder1_position[11]), .\encoder1_position[12] (encoder1_position[12]), 
            .\encoder1_position[13] (encoder1_position[13]), .\encoder1_position[14] (encoder1_position[14]), 
            .\encoder1_position[15] (encoder1_position[15]), .\encoder1_position[16] (encoder1_position[16]), 
            .\encoder1_position[17] (encoder1_position[17]), .\encoder1_position[18] (encoder1_position[18]), 
            .\encoder1_position[19] (encoder1_position[19]), .\encoder1_position[20] (encoder1_position[20]), 
            .\encoder1_position[21] (encoder1_position[21]), .\encoder1_position[22] (encoder1_position[22]), 
            .\encoder1_position[23] (encoder1_position[23]), .n1905(n1905), 
            .n1903(n1903), .n1901(n1901), .n1899(n1899), .n1897(n1897), 
            .n1895(n1895), .n1893(n1893), .n1891(n1891), .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[49] 318[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2072 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [0]), 
            .O(n52245));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2072.LUT_INIT = 16'h2300;
    SB_LUT4 i13270_3_lut_4_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26976));   // verilog/coms.v(130[12] 305[6])
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[15] [1]), 
            .O(n52244));   // verilog/TinyFPGA_B.v(361[10] 391[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    pwm PWM (.n2978(n2978), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .pwm_setpoint({pwm_setpoint}), 
        .GND_net(GND_net), .reset(reset), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, GND_net, state, 
            VCC_net, n20312, bit_ctr, n7, \neopxl_color[9] , \neopxl_color[8] , 
            \color_bit_N_478[1] , n27543, n51153, n25081, \bit_ctr[3] , 
            \bit_ctr[4] , NEOPXL_c, \neopxl_color[16] , \neopxl_color[17] , 
            \neopxl_color[18] , \neopxl_color[19] , \neopxl_color[22] , 
            \neopxl_color[23] , \neopxl_color[20] , \neopxl_color[21] , 
            LED_c, n38354, n47529, n56665, n56663, n62592, n62640, 
            \neopxl_color[10] , \neopxl_color[11] , n62472, n47509) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    input GND_net;
    output [1:0]state;
    input VCC_net;
    output n20312;
    output [4:0]bit_ctr;
    output n7;
    input \neopxl_color[9] ;
    input \neopxl_color[8] ;
    output \color_bit_N_478[1] ;
    input n27543;
    input n51153;
    output n25081;
    output \bit_ctr[3] ;
    output \bit_ctr[4] ;
    output NEOPXL_c;
    input \neopxl_color[16] ;
    input \neopxl_color[17] ;
    input \neopxl_color[18] ;
    input \neopxl_color[19] ;
    input \neopxl_color[22] ;
    input \neopxl_color[23] ;
    input \neopxl_color[20] ;
    input \neopxl_color[21] ;
    input LED_c;
    output n38354;
    output n47529;
    input n56665;
    input n56663;
    input n62592;
    input n62640;
    input \neopxl_color[10] ;
    input \neopxl_color[11] ;
    output n62472;
    output n47509;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_492 , n52360, \neo_pixel_transmitter.done , 
        start_N_483, n7_c, start, n7_adj_5672, n7_adj_5673, n38427, 
        n38365, n18, n21, n4;
    wire [10:0]one_wire_N_455;
    
    wire n38346, n22780, n46958, n4_adj_5674, n38431, n59356, n53268, 
        n12, n53302, n27183;
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n56405, n12_adj_5675, n56507, n39, n55225, n27182, n27181, 
        n27180, n27179, n27178, n27177, n27176, n27175;
    wire [10:0]n13;
    
    wire n27174;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n45571, n4_adj_5677, n45570, n45569, n45568, n45567, n45566, 
        n45565, n45564, n45563, n45562;
    wire [5:0]color_bit_N_478;
    
    wire n62601, n62604;
    wire [10:0]n49;
    
    wire n26964;
    wire [31:0]n137;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(17[11:18])
    
    wire n26268, n1, n25091, n26180;
    wire [1:0]state_1__N_416;
    
    wire n24980, n26270, \neo_pixel_transmitter.done_N_500 , n61376, 
        n55243, n46075, n46074, n46073, n46072, n46071, n46070, 
        n46069, n46068, n46067, n46066, n56696, n56697, n56715, 
        n56714, n57_adj_5681, n38419, n6822, n22859, n22860, n57827, 
        n4_adj_5682, n4_adj_5683, n59360, n53406, n53418, n61375, 
        n2943, n56592, n56591, n56593, n62469, n6_adj_5684;
    
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n52360), .D(\neo_pixel_transmitter.done_N_492 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7_c), .D(start_N_483));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i2_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5672));
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut (.I0(n7_adj_5673), .I1(n7_adj_5672), .I2(n38427), 
            .I3(n38365), .O(n18));
    defparam i1_4_lut.LUT_INIT = 16'h7350;
    SB_LUT4 i47259_4_lut (.I0(state[1]), .I1(state[0]), .I2(n21), .I3(n18), 
            .O(n4));
    defparam i47259_4_lut.LUT_INIT = 16'h5410;
    SB_LUT4 i24755_3_lut (.I0(one_wire_N_455[8]), .I1(one_wire_N_455[10]), 
            .I2(one_wire_N_455[9]), .I3(GND_net), .O(n38346));
    defparam i24755_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i38377_4_lut (.I0(n22780), .I1(n46958), .I2(n4_adj_5674), 
            .I3(state[0]), .O(n38431));   // verilog/neopixel.v(35[4] 115[11])
    defparam i38377_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i44920_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n59356));
    defparam i44920_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i38419_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n38431), .I3(GND_net), .O(n53268));
    defparam i38419_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut (.I0(n53268), .I1(n59356), .I2(state[1]), .I3(n38346), 
            .O(n7_c));
    defparam i15_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i47392_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_483));   // verilog/neopixel.v(35[4] 115[11])
    defparam i47392_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut_adj_1767 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5673));
    defparam i2_2_lut_adj_1767.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(one_wire_N_455[7]), .I1(one_wire_N_455[9]), .I2(one_wire_N_455[4]), 
            .I3(one_wire_N_455[6]), .O(n12));   // verilog/neopixel.v(61[15:42])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_455[8]), .I1(n12), .I2(one_wire_N_455[5]), 
            .I3(one_wire_N_455[10]), .O(n22780));   // verilog/neopixel.v(61[15:42])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i38453_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n53302));
    defparam i38453_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24833_2_lut (.I0(n22780), .I1(n46958), .I2(GND_net), .I3(GND_net), 
            .O(n38427));
    defparam i24833_2_lut.LUT_INIT = 16'heeee;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n27183));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i1_2_lut (.I0(one_wire_N_455[2]), .I1(one_wire_N_455[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5674));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41515_2_lut (.I0(one_wire_N_455[4]), .I1(n4_adj_5674), .I2(GND_net), 
            .I3(GND_net), .O(n56405));
    defparam i41515_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(one_wire_N_455[10]), 
            .I2(state[0]), .I3(GND_net), .O(n12_adj_5675));
    defparam i3_3_lut.LUT_INIT = 16'h2121;
    SB_LUT4 i41616_4_lut (.I0(one_wire_N_455[6]), .I1(one_wire_N_455[9]), 
            .I2(one_wire_N_455[8]), .I3(n56405), .O(n56507));
    defparam i41616_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i65_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(one_wire_N_455[7]), .I1(n56507), .I2(n12_adj_5675), 
            .I3(one_wire_N_455[5]), .O(n55225));
    defparam i8_4_lut.LUT_INIT = 16'h0010;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n27182));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i47484_4_lut (.I0(n38427), .I1(n53302), .I2(n55225), .I3(n39), 
            .O(n52360));
    defparam i47484_4_lut.LUT_INIT = 16'hcecf;
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n27181));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n27180));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n27179));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n27178));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n27177));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n27176));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n27175));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n27174));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n45571), .O(one_wire_N_455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1768 (.I0(one_wire_N_455[3]), .I1(one_wire_N_455[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5677));
    defparam i1_2_lut_adj_1768.LUT_INIT = 16'h8888;
    SB_LUT4 sub_67_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n13[9]), 
            .I3(n45570), .O(one_wire_N_455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_67_add_2_11 (.CI(n45570), .I0(timer[9]), .I1(n13[9]), 
            .CO(n45571));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n45569), .O(one_wire_N_455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n45569), .I0(timer[8]), .I1(n13[8]), 
            .CO(n45570));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n45568), .O(one_wire_N_455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n45568), .I0(timer[7]), .I1(n13[7]), 
            .CO(n45569));
    SB_LUT4 sub_67_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n13[6]), 
            .I3(n45567), .O(one_wire_N_455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_8 (.CI(n45567), .I0(timer[6]), .I1(n13[6]), 
            .CO(n45568));
    SB_LUT4 sub_67_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n13[5]), 
            .I3(n45566), .O(one_wire_N_455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_67_add_2_7 (.CI(n45566), .I0(timer[5]), .I1(n13[5]), 
            .CO(n45567));
    SB_LUT4 sub_67_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n45565), .O(one_wire_N_455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_67_add_2_6 (.CI(n45565), .I0(timer[4]), .I1(n13[4]), 
            .CO(n45566));
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n45564), .O(one_wire_N_455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n45564), .I0(timer[3]), .I1(n13[3]), 
            .CO(n45565));
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n45563), .O(one_wire_N_455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_4 (.CI(n45563), .I0(timer[2]), .I1(n13[2]), 
            .CO(n45564));
    SB_LUT4 sub_67_add_2_3_lut (.I0(n4_adj_5677), .I1(timer[1]), .I2(n13[1]), 
            .I3(n45562), .O(n46958)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_67_add_2_3 (.CI(n45562), .I0(timer[1]), .I1(n13[1]), 
            .CO(n45563));
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n45562));
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(n38431), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n20312));   // verilog/neopixel.v(35[4] 115[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(color_bit_N_478[2]), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hf6f6;
    SB_LUT4 n62601_bdd_4_lut (.I0(n62601), .I1(\neopxl_color[9] ), .I2(\neopxl_color[8] ), 
            .I3(\color_bit_N_478[1] ), .O(n62604));
    defparam n62601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF timer_1929__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n26964));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(VCC_net), .D(n27543));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n51153));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n25081), 
            .D(n137[2]), .R(n26268));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(\bit_ctr[3] ), .C(clk16MHz), .E(n25081), 
            .D(n137[3]), .R(n26268));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n25081), 
            .D(n137[4]), .R(n26268));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n25091), .D(n1), 
            .R(n26180));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n24980), .D(state_1__N_416[0]), 
            .S(n26270));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n61376), .D(\neo_pixel_transmitter.done_N_500 ), 
            .R(n55243));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1929__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1929__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 timer_1929_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n46075), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1929_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n46074), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_11 (.CI(n46074), .I0(GND_net), .I1(timer[9]), 
            .CO(n46075));
    SB_LUT4 timer_1929_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n46073), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_10 (.CI(n46073), .I0(GND_net), .I1(timer[8]), 
            .CO(n46074));
    SB_LUT4 timer_1929_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n46072), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_9 (.CI(n46072), .I0(GND_net), .I1(timer[7]), 
            .CO(n46073));
    SB_LUT4 timer_1929_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n46071), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_8 (.CI(n46071), .I0(GND_net), .I1(timer[6]), 
            .CO(n46072));
    SB_LUT4 timer_1929_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n46070), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_7 (.CI(n46070), .I0(GND_net), .I1(timer[5]), 
            .CO(n46071));
    SB_LUT4 timer_1929_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n46069), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_6 (.CI(n46069), .I0(GND_net), .I1(timer[4]), 
            .CO(n46070));
    SB_LUT4 timer_1929_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n46068), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_5 (.CI(n46068), .I0(GND_net), .I1(timer[3]), 
            .CO(n46069));
    SB_LUT4 timer_1929_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n46067), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_4 (.CI(n46067), .I0(GND_net), .I1(timer[2]), 
            .CO(n46068));
    SB_LUT4 timer_1929_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n46066), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_3 (.CI(n46066), .I0(GND_net), .I1(timer[1]), 
            .CO(n46067));
    SB_LUT4 timer_1929_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1929_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1929_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n46066));
    SB_LUT4 i41796_3_lut (.I0(\neopxl_color[16] ), .I1(\neopxl_color[17] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56696));
    defparam i41796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41797_3_lut (.I0(\neopxl_color[18] ), .I1(\neopxl_color[19] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56697));
    defparam i41797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41815_3_lut (.I0(\neopxl_color[22] ), .I1(\neopxl_color[23] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56715));
    defparam i41815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41814_3_lut (.I0(\neopxl_color[20] ), .I1(\neopxl_color[21] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n56714));
    defparam i41814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5681), .I2(LED_c), 
            .I3(state[1]), .O(n25091));   // verilog/neopixel.v(35[4] 115[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i12474_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5681), .I2(LED_c), 
            .I3(state[1]), .O(n26180));   // verilog/neopixel.v(35[4] 115[11])
    defparam i12474_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_adj_1769 (.I0(\bit_ctr[3] ), .I1(n38354), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n47529));
    defparam i1_2_lut_3_lut_adj_1769.LUT_INIT = 16'h7878;
    SB_LUT4 i24824_2_lut_3_lut (.I0(\bit_ctr[3] ), .I1(n38354), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n38419));
    defparam i24824_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1770 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(color_bit_N_478[2]));
    defparam i1_2_lut_3_lut_adj_1770.LUT_INIT = 16'h1e1e;
    SB_LUT4 i24763_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n38354));
    defparam i24763_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1771 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_478[1] ));
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'h6666;
    SB_LUT4 i2085_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2085_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2099_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n6822), .I2(\bit_ctr[3] ), 
            .I3(\bit_ctr[4] ), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2099_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i1_2_lut_4_lut_adj_1772 (.I0(n22780), .I1(n46958), .I2(start), 
            .I3(\neo_pixel_transmitter.done ), .O(n22859));   // verilog/neopixel.v(78[18] 98[12])
    defparam i1_2_lut_4_lut_adj_1772.LUT_INIT = 16'hf1ff;
    SB_LUT4 i1_2_lut_3_lut_adj_1773 (.I0(n38365), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n22860));   // verilog/neopixel.v(51[18] 71[12])
    defparam i1_2_lut_3_lut_adj_1773.LUT_INIT = 16'hdfdf;
    SB_LUT4 i42927_2_lut_3_lut (.I0(n47529), .I1(\bit_ctr[3] ), .I2(n38354), 
            .I3(GND_net), .O(n57827));   // verilog/neopixel.v(21[26:38])
    defparam i42927_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i1_2_lut_3_lut_adj_1774 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n38431), .I3(GND_net), .O(n4_adj_5682));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut_adj_1774.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_1775 (.I0(n22780), .I1(start), .I2(state[1]), 
            .I3(GND_net), .O(n4_adj_5683));
    defparam i1_2_lut_3_lut_adj_1775.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n38346), .I1(state[1]), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n55243));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i44955_2_lut (.I0(n22780), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n59360));
    defparam i44955_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51_4_lut (.I0(n59360), .I1(n38346), .I2(state[1]), .I3(n4_adj_5674), 
            .O(n53406));
    defparam i51_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i50_3_lut (.I0(n46958), .I1(n4_adj_5674), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n53418));
    defparam i50_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46475_4_lut (.I0(n53406), .I1(n53302), .I2(\neo_pixel_transmitter.done ), 
            .I3(n38427), .O(n61375));
    defparam i46475_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i46476_4_lut (.I0(n61375), .I1(n53418), .I2(state[0]), .I3(n4_adj_5683), 
            .O(n61376));
    defparam i46476_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i2_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_500 ));
    defparam i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i609_2_lut (.I0(n38346), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n2943));   // verilog/neopixel.v(102[9] 110[12])
    defparam i609_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1776 (.I0(n4_adj_5682), .I1(state[0]), .I2(state[1]), 
            .I3(n2943), .O(n26270));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15_4_lut_adj_1776.LUT_INIT = 16'h0a3a;
    SB_LUT4 i20_4_lut (.I0(n4_adj_5682), .I1(n2943), .I2(state[1]), .I3(state[0]), 
            .O(n24980));
    defparam i20_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i41692_4_lut (.I0(n56665), .I1(n56663), .I2(n47529), .I3(\color_bit_N_478[1] ), 
            .O(n56592));
    defparam i41692_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i41691_3_lut (.I0(n62592), .I1(n62640), .I2(color_bit_N_478[2]), 
            .I3(GND_net), .O(n56591));
    defparam i41691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41693_4_lut (.I0(n56592), .I1(n62604), .I2(n47529), .I3(color_bit_N_478[2]), 
            .O(n56593));
    defparam i41693_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i24272_4_lut (.I0(n56593), .I1(n57_adj_5681), .I2(n56591), 
            .I3(n57827), .O(state_1__N_416[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i24272_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n22859), .I1(n22860), .I2(state[0]), 
            .I3(bit_ctr[0]), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 i2092_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(\bit_ctr[3] ), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2092_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(\neopxl_color[10] ), 
            .I2(\neopxl_color[11] ), .I3(bit_ctr[1]), .O(n62601));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 color_bit_N_478_1__bdd_4_lut_47694 (.I0(\color_bit_N_478[1] ), 
            .I1(n56714), .I2(n56715), .I3(color_bit_N_478[2]), .O(n62469));
    defparam color_bit_N_478_1__bdd_4_lut_47694.LUT_INIT = 16'he4aa;
    SB_LUT4 i2080_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6822));   // verilog/neopixel.v(68[23:32])
    defparam i2080_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n62469_bdd_4_lut (.I0(n62469), .I1(n56697), .I2(n56696), .I3(color_bit_N_478[2]), 
            .O(n62472));
    defparam n62469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 state_1__I_0_i3_3_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_492 ));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_i3_3_lut_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i13477_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[1]), 
            .I3(\neo_pixel_transmitter.t0 [1]), .O(n27183));
    defparam i13477_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13468_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[10]), 
            .I3(\neo_pixel_transmitter.t0 [10]), .O(n27174));
    defparam i13468_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13469_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[9]), 
            .I3(\neo_pixel_transmitter.t0 [9]), .O(n27175));
    defparam i13469_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13470_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[8]), 
            .I3(\neo_pixel_transmitter.t0 [8]), .O(n27176));
    defparam i13470_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13471_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[7]), 
            .I3(\neo_pixel_transmitter.t0 [7]), .O(n27177));
    defparam i13471_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13472_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[6]), 
            .I3(\neo_pixel_transmitter.t0 [6]), .O(n27178));
    defparam i13472_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13473_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[5]), 
            .I3(\neo_pixel_transmitter.t0 [5]), .O(n27179));
    defparam i13473_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13474_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[4]), 
            .I3(\neo_pixel_transmitter.t0 [4]), .O(n27180));
    defparam i13474_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13475_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[3]), 
            .I3(\neo_pixel_transmitter.t0 [3]), .O(n27181));
    defparam i13475_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13476_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[2]), 
            .I3(\neo_pixel_transmitter.t0 [2]), .O(n27182));
    defparam i13476_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13258_3_lut_4_lut (.I0(start_N_483), .I1(n4), .I2(timer[0]), 
            .I3(\neo_pixel_transmitter.t0 [0]), .O(n26964));
    defparam i13258_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1777 (.I0(\bit_ctr[3] ), .I1(n38354), .I2(GND_net), 
            .I3(GND_net), .O(n47509));
    defparam i1_2_lut_adj_1777.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1778 (.I0(n47529), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5684));
    defparam i1_2_lut_adj_1778.LUT_INIT = 16'hdddd;
    SB_LUT4 i1060_4_lut (.I0(n7), .I1(n38419), .I2(n47509), .I3(n6_adj_5684), 
            .O(n57_adj_5681));   // verilog/neopixel.v(21[26:38])
    defparam i1060_4_lut.LUT_INIT = 16'h3323;
    SB_LUT4 i1_3_lut (.I0(n25091), .I1(n20312), .I2(state[1]), .I3(GND_net), 
            .O(n25081));
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i12563_2_lut (.I0(n25081), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n26268));   // verilog/neopixel.v(34[12] 116[6])
    defparam i12563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n38365), .I3(n38427), .O(n21));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5410;
    SB_LUT4 i2_2_lut_3_lut_adj_1779 (.I0(n22780), .I1(one_wire_N_455[2]), 
            .I2(one_wire_N_455[3]), .I3(GND_net), .O(n38365));
    defparam i2_2_lut_3_lut_adj_1779.LUT_INIT = 16'hfefe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (GND_net, \byte_transmit_counter[4] , \byte_transmit_counter[0] , 
            \byte_transmit_counter[2] , \byte_transmit_counter[1] , \byte_transmit_counter[3] , 
            \data_in_frame[12] , clk16MHz, n2978, \data_out_frame[10] , 
            n52280, n52279, \data_out_frame[1][5] , n52310, n52278, 
            tx_active, n26953, \data_in_frame[13] , \data_out_frame[0][3] , 
            \data_out_frame[1][3] , \data_out_frame[3][3] , \data_out_frame[6] , 
            \data_out_frame[7] , \data_out_frame[4] , \data_out_frame[5] , 
            \FRAME_MATCHER.i_31__N_2485 , encoder0_position_scaled, n52309, 
            \data_out_frame[1][6] , n52308, control_mode, n3543, n52307, 
            \data_out_frame[1][7] , n52306, n26957, n26691, n52154, 
            n52305, n26960, n52304, n52318, n52303, n52158, n26969, 
            \data_in_frame[13][4] , n26972, \data_in_frame[13][5] , n27218, 
            VCC_net, \data_in_frame[18] , n26979, \data_in_frame[13][6] , 
            n26982, \data_in_frame[13][7] , n27213, \data_in_frame[14] , 
            n27203, n27200, encoder1_position_scaled, \data_out_frame[12] , 
            setpoint, \data_out_frame[11] , \data_out_frame[18] , \data_out_frame[19] , 
            n52156, \data_out_frame[17] , \data_out_frame[16] , n62658, 
            \data_out_frame[9] , \data_out_frame[8] , \data_in_frame[15] , 
            Kp_23__N_1724, reset, n27192, n52277, n52276, n52275, 
            n52274, n52273, n52272, n52271, n52270, n52269, n52268, 
            n52267, n52266, n52265, n52264, rx_data_ready, \FRAME_MATCHER.rx_data_ready_prev , 
            \FRAME_MATCHER.i[1] , \FRAME_MATCHER.i[2] , n35706, n27101, 
            \data_in_frame[16] , n27105, \data_in_frame[2] , \Kp[5] , 
            n30905, n27148, n27130, ID, \data_in_frame[0][7] , n27144, 
            n27133, n52263, n27136, \data_in_frame[16][4] , n27129, 
            deadband, n27128, n27127, n27126, n26731, \data_in_frame[5] , 
            n26734, n26737, n26740, n51817, n27772, \data_in_frame[4] , 
            n27124, n27123, n27122, n27121, n27120, n26743, n51681, 
            n51677, n27312, n27317, n51673, n27321, n26746, n26749, 
            n27327, \data_in_frame[2][7] , n27331, \data_in_frame[3][0] , 
            n27757, \data_in_frame[6][1] , n51669, \data_in_frame[3][1] , 
            n51667, \data_in_frame[3][2] , n51663, \data_in_frame[3][3] , 
            n51659, \data_in_frame[3][4] , n27119, n27118, n27117, 
            n27116, n27115, n27114, n27113, n27112, n27111, n27110, 
            n51655, \data_in_frame[3][7] , n27365, n27370, n27375, 
            n27379, n27387, n27391, n27430, \data_in_frame[18][7] , 
            n27433, n51579, \data_in_frame[19] , n27439, n27109, n27108, 
            n27104, n27100, neopxl_color, n27099, n27097, n27096, 
            n27095, n27094, n27093, n27092, n27091, n27662, \data_in_frame[20] , 
            n27659, n20140, n27090, n27089, n27088, n27087, n27086, 
            n27085, n27084, n27083, n27082, n27081, n27080, n27656, 
            n27653, n27650, n27647, n27644, n27079, n27078, n51577, 
            n51575, \data_in_frame[6][2] , \data_in_frame[6][3] , n27637, 
            n27062, IntegralLimit, n27061, n27056, n27055, n27054, 
            n27053, \Ki[15] , n27052, current_limit, n27051, \Ki[13] , 
            n27050, n27049, \Ki[11] , n27048, \Ki[10] , n27047, 
            \Ki[9] , n27046, \Ki[8] , n27045, \Ki[7] , n27044, \Ki[6] , 
            n27043, \Ki[5] , n27042, \Ki[4] , n27041, \Ki[3] , n27040, 
            \Ki[2] , n27039, n27038, \Ki[1] , n27028, \Kp[15] , 
            \Kp[14] , n27614, PWMLimit, n27613, n27612, n27611, 
            n27609, n27608, n27023, \Kp[13] , n27022, \Kp[12] , 
            n27021, \Kp[11] , n27020, \Kp[10] , n27019, n27018, 
            \Ki[14] , n27607, n27606, n27605, n27604, n27603, n27602, 
            n27601, n27600, n27599, n27598, n27017, \Ki[12] , n27016, 
            n27597, n27595, n27594, n27593, n27590, \data_in_frame[6][4] , 
            n27015, n27014, n27010, \data_in_frame[6][6] , n52302, 
            n26986, n26985, \data_in_frame[6][7] , n51567, n51549, 
            n27551, n26978, \data_out_frame[25] , \data_out_frame[24] , 
            n26977, n26976, n26705, \data_out_frame[1][0] , n52317, 
            n52316, \data_out_frame[1][1] , n52315, n52314, n52313, 
            n52312, n52311, n52157, n26975, n26968, n26956, \data_out_frame[0][2] , 
            n52218, n52301, n26946, n26944, n26930, \Kp[1] , n26929, 
            \Kp[2] , n26925, \Kp[3] , n26924, \Kp[4] , n26920, n26916, 
            \Ki[0] , n26915, \Kp[0] , n52262, \motor_state_23__N_67[13] , 
            n15, n9, n52261, n52260, n52259, \data_out_frame[13] , 
            n52258, n52257, n52256, n52255, n52254, n52160, n52253, 
            n52252, \data_out_frame[14] , n52251, n52250, n52249, 
            n52248, n26347, n52247, n52246, n52217, \data_out_frame[15] , 
            n52245, n52244, n52243, n52242, n27549, \data_in_frame[8] , 
            \data_in_frame[8][4] , \data_in_frame[8][5] , \data_in_frame[8][6] , 
            \data_in_frame[8][7] , n51565, \data_in_frame[9] , n52409, 
            \FRAME_MATCHER.i[0] , n62586, \FRAME_MATCHER.state[3] , n52430, 
            rx_data, \data_out_frame[22] , \data_out_frame[23] , \data_out_frame[21] , 
            \data_out_frame[20] , n62532, n52241, n52240, n52239, 
            n52223, n52238, n52237, n52236, n52235, n52234, n52233, 
            n52232, n52231, n27935, n26327, n52230, n52229, n52228, 
            n52227, n52226, n52225, n52155, n26319, n52220, n59364, 
            n62466, n27945, n26317, n52221, n52222, n52224, n52159, 
            n52219, n52161, n52162, n52163, n52164, n52165, n52166, 
            n52167, n52168, n52169, n27960, n26302, n52170, n27962, 
            n26300, n52171, n52172, n52173, n52174, n52175, n27968, 
            n26294, n52176, n27970, n26292, n52177, n52178, n52179, 
            n52180, n52181, n52182, n52183, n27978, n26284, n27979, 
            n26283, n52184, n27981, n26281, n52185, n52186, n52187, 
            n27985, n26277, n27986, n26276, n54720, n27987, n26275, 
            n52188, n52189, n52190, n52191, n52192, n52193, n52194, 
            n52195, n52196, n52197, n52198, n52199, n52200, n52201, 
            n52202, n52203, n52204, n52205, n52206, \data_in_frame[11] , 
            n4, \data_in_frame[10] , \data_out_frame[26][2] , \data_in_frame[10][7] , 
            \data_out_frame[27][2] , n23375, Kp_23__N_645, n52455, \Kp[6] , 
            n52656, n26787, \Kp[7] , n26786, n25709, n25766, \data_out_frame[3][1] , 
            n52207, n52208, \data_out_frame[3][4] , n52209, \data_out_frame[3][6] , 
            n52210, \data_out_frame[3][7] , n52211, n52212, n26782, 
            n28044, n26215, n52213, n28046, n26213, n52214, n52215, 
            n28052, n26207, LED_c, n52216, DE_c, n26769, \Kp[8] , 
            n26768, \Kp[9] , n52300, \data_out_frame[0][4] , n52299, 
            n52298, n52297, n52296, n52295, n28093, n26402, n52294, 
            n28095, n26400, n28096, n26399, n52293, n52292, n52291, 
            n52290, n52289, n52288, n52287, n26391, n28105, n26390, 
            n52286, \data_in_frame[10][0] , \data_in_frame[10][1] , \data_in_frame[10][2] , 
            \data_in_frame[10][3] , \data_in_frame[10][4] , n51563, n51585, 
            n51561, n51559, n51557, n51555, n51553, n51551, n52285, 
            n52284, n52283, n52282, n28111, n26384, n22568, n23824, 
            n53055, n52281, n10, n38306, n25768, n47452, n52831, 
            n52848, n23338, n47989, n16, n53140, n52878, Kp_23__N_969, 
            Kp_23__N_675, n3, n375, n11, n53137, n11_adj_8, n52925, 
            n13, n52424, n38302, n52412, n10_adj_9, n25739, n23958, 
            n1513, n52564, n35696, n53098, n25705, n52842, n47380, 
            n23427, n53035, n25707, n23531, n22594, n23688, n1130, 
            n23945, n32, n53161, n56674, n56672, n52053, n151, 
            n203, n181, n155, \PID_CONTROLLER.integral_23__N_3691[3] , 
            \current[11] , \data[11] , n25021, n27452, displacement, 
            n15_adj_10, n15_adj_11, \motor_state_23__N_67[17] , n2076, 
            n52979, n52928, n23594, n53122, n68, n62598, n59386, 
            n25356, n52922, n52641, n56668, n56666, n53069, n52513, 
            n12, n8, n52434, n25346, n52939, n52741, n25699, n204, 
            n6, n152, n60212, n53113, n53125, n52496, n25734, 
            n10_adj_12, n25750, n35727, \current[7] , \current[6] , 
            \current[5] , \current[4] , \current[3] , \current[2] , 
            \current[1] , \current[0] , \current[15] , \current[10] , 
            \current[9] , \current[8] , n62688, n62430, pwm_setpoint, 
            n52427, n62840, r_SM_Main, r_Clock_Count, tx_o, n26943, 
            \tx_data[2] , n23, \o_Rx_DV_N_3464[12] , n4858, \o_Rx_DV_N_3464[24] , 
            n27, n29, n6_adj_13, tx_enable, n27247, baudrate, n55830, 
            n27246, n27245, n27243, n27242, \o_Rx_DV_N_3464[8] , n4855, 
            n52352, \r_SM_Main[1]_adj_14 , n25039, n27241, n27240, 
            \r_SM_Main[2]_adj_15 , n55782, r_Clock_Count_adj_24, n55798, 
            n55750, n55766, r_Rx_Data, RX_N_2, n22878, \o_Rx_DV_N_3464[7] , 
            \o_Rx_DV_N_3464[6] , \o_Rx_DV_N_3464[5] , \o_Rx_DV_N_3464[4] , 
            \o_Rx_DV_N_3464[3] , \o_Rx_DV_N_3464[2] , \o_Rx_DV_N_3464[1] , 
            \o_Rx_DV_N_3464[0] , n25264, n27583, n48661, n27579, \r_Bit_Index[0] , 
            n53350, n55734, n55846, n55814) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \byte_transmit_counter[4] ;
    output \byte_transmit_counter[0] ;
    output \byte_transmit_counter[2] ;
    output \byte_transmit_counter[1] ;
    output \byte_transmit_counter[3] ;
    output [7:0]\data_in_frame[12] ;
    input clk16MHz;
    input n2978;
    output [7:0]\data_out_frame[10] ;
    input n52280;
    input n52279;
    output \data_out_frame[1][5] ;
    input n52310;
    input n52278;
    output tx_active;
    input n26953;
    output [7:0]\data_in_frame[13] ;
    output \data_out_frame[0][3] ;
    output \data_out_frame[1][3] ;
    output \data_out_frame[3][3] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output \FRAME_MATCHER.i_31__N_2485 ;
    input [23:0]encoder0_position_scaled;
    input n52309;
    output \data_out_frame[1][6] ;
    input n52308;
    output [7:0]control_mode;
    output n3543;
    input n52307;
    output \data_out_frame[1][7] ;
    input n52306;
    input n26957;
    input n26691;
    input n52154;
    input n52305;
    input n26960;
    input n52304;
    input n52318;
    input n52303;
    input n52158;
    input n26969;
    output \data_in_frame[13][4] ;
    input n26972;
    output \data_in_frame[13][5] ;
    input n27218;
    input VCC_net;
    output [7:0]\data_in_frame[18] ;
    input n26979;
    output \data_in_frame[13][6] ;
    input n26982;
    output \data_in_frame[13][7] ;
    input n27213;
    output [7:0]\data_in_frame[14] ;
    input n27203;
    input n27200;
    input [23:0]encoder1_position_scaled;
    output [7:0]\data_out_frame[12] ;
    output [23:0]setpoint;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    input n52156;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[16] ;
    output n62658;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_in_frame[15] ;
    output Kp_23__N_1724;
    input reset;
    input n27192;
    input n52277;
    input n52276;
    input n52275;
    input n52274;
    input n52273;
    input n52272;
    input n52271;
    input n52270;
    input n52269;
    input n52268;
    input n52267;
    input n52266;
    input n52265;
    input n52264;
    output rx_data_ready;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output \FRAME_MATCHER.i[1] ;
    output \FRAME_MATCHER.i[2] ;
    output n35706;
    input n27101;
    output [7:0]\data_in_frame[16] ;
    input n27105;
    output [7:0]\data_in_frame[2] ;
    output \Kp[5] ;
    output n30905;
    input n27148;
    input n27130;
    input [7:0]ID;
    output \data_in_frame[0][7] ;
    input n27144;
    input n27133;
    input n52263;
    input n27136;
    output \data_in_frame[16][4] ;
    input n27129;
    output [23:0]deadband;
    input n27128;
    input n27127;
    input n27126;
    input n26731;
    output [7:0]\data_in_frame[5] ;
    input n26734;
    input n26737;
    input n26740;
    input n51817;
    input n27772;
    output [7:0]\data_in_frame[4] ;
    input n27124;
    input n27123;
    input n27122;
    input n27121;
    input n27120;
    input n26743;
    input n51681;
    input n51677;
    input n27312;
    input n27317;
    input n51673;
    input n27321;
    input n26746;
    input n26749;
    input n27327;
    output \data_in_frame[2][7] ;
    input n27331;
    output \data_in_frame[3][0] ;
    input n27757;
    output \data_in_frame[6][1] ;
    input n51669;
    output \data_in_frame[3][1] ;
    input n51667;
    output \data_in_frame[3][2] ;
    input n51663;
    output \data_in_frame[3][3] ;
    input n51659;
    output \data_in_frame[3][4] ;
    input n27119;
    input n27118;
    input n27117;
    input n27116;
    input n27115;
    input n27114;
    input n27113;
    input n27112;
    input n27111;
    input n27110;
    input n51655;
    output \data_in_frame[3][7] ;
    input n27365;
    input n27370;
    input n27375;
    input n27379;
    input n27387;
    input n27391;
    input n27430;
    output \data_in_frame[18][7] ;
    input n27433;
    input n51579;
    output [7:0]\data_in_frame[19] ;
    input n27439;
    input n27109;
    input n27108;
    input n27104;
    input n27100;
    output [23:0]neopxl_color;
    input n27099;
    input n27097;
    input n27096;
    input n27095;
    input n27094;
    input n27093;
    input n27092;
    input n27091;
    input n27662;
    output [7:0]\data_in_frame[20] ;
    input n27659;
    output n20140;
    input n27090;
    input n27089;
    input n27088;
    input n27087;
    input n27086;
    input n27085;
    input n27084;
    input n27083;
    input n27082;
    input n27081;
    input n27080;
    input n27656;
    input n27653;
    input n27650;
    input n27647;
    input n27644;
    input n27079;
    input n27078;
    input n51577;
    input n51575;
    output \data_in_frame[6][2] ;
    output \data_in_frame[6][3] ;
    input n27637;
    input n27062;
    output [23:0]IntegralLimit;
    input n27061;
    input n27056;
    input n27055;
    input n27054;
    input n27053;
    output \Ki[15] ;
    input n27052;
    output [15:0]current_limit;
    input n27051;
    output \Ki[13] ;
    input n27050;
    input n27049;
    output \Ki[11] ;
    input n27048;
    output \Ki[10] ;
    input n27047;
    output \Ki[9] ;
    input n27046;
    output \Ki[8] ;
    input n27045;
    output \Ki[7] ;
    input n27044;
    output \Ki[6] ;
    input n27043;
    output \Ki[5] ;
    input n27042;
    output \Ki[4] ;
    input n27041;
    output \Ki[3] ;
    input n27040;
    output \Ki[2] ;
    input n27039;
    input n27038;
    output \Ki[1] ;
    input n27028;
    output \Kp[15] ;
    output \Kp[14] ;
    input n27614;
    output [23:0]PWMLimit;
    input n27613;
    input n27612;
    input n27611;
    input n27609;
    input n27608;
    input n27023;
    output \Kp[13] ;
    input n27022;
    output \Kp[12] ;
    input n27021;
    output \Kp[11] ;
    input n27020;
    output \Kp[10] ;
    input n27019;
    input n27018;
    output \Ki[14] ;
    input n27607;
    input n27606;
    input n27605;
    input n27604;
    input n27603;
    input n27602;
    input n27601;
    input n27600;
    input n27599;
    input n27598;
    input n27017;
    output \Ki[12] ;
    input n27016;
    input n27597;
    input n27595;
    input n27594;
    input n27593;
    input n27590;
    output \data_in_frame[6][4] ;
    input n27015;
    input n27014;
    input n27010;
    output \data_in_frame[6][6] ;
    input n52302;
    input n26986;
    input n26985;
    output \data_in_frame[6][7] ;
    input n51567;
    input n51549;
    input n27551;
    input n26978;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    input n26977;
    input n26976;
    input n26705;
    output \data_out_frame[1][0] ;
    input n52317;
    input n52316;
    output \data_out_frame[1][1] ;
    input n52315;
    input n52314;
    input n52313;
    input n52312;
    input n52311;
    input n52157;
    input n26975;
    input n26968;
    input n26956;
    output \data_out_frame[0][2] ;
    input n52218;
    input n52301;
    input n26946;
    input n26944;
    input n26930;
    output \Kp[1] ;
    input n26929;
    output \Kp[2] ;
    input n26925;
    output \Kp[3] ;
    input n26924;
    output \Kp[4] ;
    input n26920;
    input n26916;
    output \Ki[0] ;
    input n26915;
    output \Kp[0] ;
    input n52262;
    input \motor_state_23__N_67[13] ;
    input n15;
    output n9;
    input n52261;
    input n52260;
    input n52259;
    output [7:0]\data_out_frame[13] ;
    input n52258;
    input n52257;
    input n52256;
    input n52255;
    input n52254;
    input n52160;
    input n52253;
    input n52252;
    output [7:0]\data_out_frame[14] ;
    input n52251;
    input n52250;
    input n52249;
    input n52248;
    input n26347;
    input n52247;
    input n52246;
    input n52217;
    output [7:0]\data_out_frame[15] ;
    input n52245;
    input n52244;
    input n52243;
    input n52242;
    input n27549;
    output [7:0]\data_in_frame[8] ;
    output \data_in_frame[8][4] ;
    output \data_in_frame[8][5] ;
    output \data_in_frame[8][6] ;
    output \data_in_frame[8][7] ;
    input n51565;
    output [7:0]\data_in_frame[9] ;
    input n52409;
    output \FRAME_MATCHER.i[0] ;
    output n62586;
    output \FRAME_MATCHER.state[3] ;
    output n52430;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[21] ;
    output [7:0]\data_out_frame[20] ;
    output n62532;
    input n52241;
    input n52240;
    input n52239;
    input n52223;
    input n52238;
    input n52237;
    input n52236;
    input n52235;
    input n52234;
    input n52233;
    input n52232;
    input n52231;
    input n27935;
    input n26327;
    input n52230;
    input n52229;
    input n52228;
    input n52227;
    input n52226;
    input n52225;
    input n52155;
    input n26319;
    input n52220;
    input n59364;
    input n62466;
    input n27945;
    input n26317;
    input n52221;
    input n52222;
    input n52224;
    input n52159;
    input n52219;
    input n52161;
    input n52162;
    input n52163;
    input n52164;
    input n52165;
    input n52166;
    input n52167;
    input n52168;
    input n52169;
    input n27960;
    input n26302;
    input n52170;
    input n27962;
    input n26300;
    input n52171;
    input n52172;
    input n52173;
    input n52174;
    input n52175;
    input n27968;
    input n26294;
    input n52176;
    input n27970;
    input n26292;
    input n52177;
    input n52178;
    input n52179;
    input n52180;
    input n52181;
    input n52182;
    input n52183;
    input n27978;
    input n26284;
    input n27979;
    input n26283;
    input n52184;
    input n27981;
    input n26281;
    input n52185;
    input n52186;
    input n52187;
    input n27985;
    input n26277;
    input n27986;
    input n26276;
    output n54720;
    input n27987;
    input n26275;
    input n52188;
    input n52189;
    input n52190;
    input n52191;
    input n52192;
    input n52193;
    input n52194;
    input n52195;
    input n52196;
    input n52197;
    input n52198;
    input n52199;
    input n52200;
    input n52201;
    input n52202;
    input n52203;
    input n52204;
    input n52205;
    input n52206;
    output [7:0]\data_in_frame[11] ;
    output n4;
    output [7:0]\data_in_frame[10] ;
    output \data_out_frame[26][2] ;
    output \data_in_frame[10][7] ;
    output \data_out_frame[27][2] ;
    input n23375;
    output Kp_23__N_645;
    output n52455;
    output \Kp[6] ;
    output n52656;
    input n26787;
    output \Kp[7] ;
    input n26786;
    input n25709;
    input n25766;
    output \data_out_frame[3][1] ;
    input n52207;
    input n52208;
    output \data_out_frame[3][4] ;
    input n52209;
    output \data_out_frame[3][6] ;
    input n52210;
    output \data_out_frame[3][7] ;
    input n52211;
    input n52212;
    input n26782;
    input n28044;
    input n26215;
    input n52213;
    input n28046;
    input n26213;
    input n52214;
    input n52215;
    input n28052;
    input n26207;
    output LED_c;
    input n52216;
    output DE_c;
    input n26769;
    output \Kp[8] ;
    input n26768;
    output \Kp[9] ;
    input n52300;
    output \data_out_frame[0][4] ;
    input n52299;
    input n52298;
    input n52297;
    input n52296;
    input n52295;
    input n28093;
    input n26402;
    input n52294;
    input n28095;
    input n26400;
    input n28096;
    input n26399;
    input n52293;
    input n52292;
    input n52291;
    input n52290;
    input n52289;
    input n52288;
    input n52287;
    input n26391;
    input n28105;
    input n26390;
    input n52286;
    output \data_in_frame[10][0] ;
    output \data_in_frame[10][1] ;
    output \data_in_frame[10][2] ;
    output \data_in_frame[10][3] ;
    output \data_in_frame[10][4] ;
    input n51563;
    input n51585;
    input n51561;
    input n51559;
    input n51557;
    input n51555;
    input n51553;
    input n51551;
    input n52285;
    input n52284;
    input n52283;
    input n52282;
    input n28111;
    input n26384;
    input n22568;
    output n23824;
    output n53055;
    input n52281;
    output n10;
    output n38306;
    input n25768;
    output n47452;
    output n52831;
    output n52848;
    output n23338;
    output n47989;
    input n16;
    output n53140;
    output n52878;
    output Kp_23__N_969;
    output Kp_23__N_675;
    output n3;
    input n375;
    output n11;
    output n53137;
    output n11_adj_8;
    output n52925;
    input n13;
    output n52424;
    output n38302;
    output n52412;
    output n10_adj_9;
    output n25739;
    output n23958;
    input n1513;
    input n52564;
    output n35696;
    output n53098;
    output n25705;
    input n52842;
    input n47380;
    input n23427;
    input n53035;
    input n25707;
    output n23531;
    output n22594;
    output n23688;
    output n1130;
    output n23945;
    output n32;
    output n53161;
    input n56674;
    input n56672;
    output n52053;
    input n151;
    input n203;
    input n181;
    input n155;
    output \PID_CONTROLLER.integral_23__N_3691[3] ;
    input \current[11] ;
    input \data[11] ;
    input n25021;
    output n27452;
    input [23:0]displacement;
    input n15_adj_10;
    input n15_adj_11;
    output \motor_state_23__N_67[17] ;
    input n2076;
    output n52979;
    input n52928;
    input n23594;
    input n53122;
    output n68;
    input n62598;
    output n59386;
    output n25356;
    input n52922;
    input n52641;
    input n56668;
    input n56666;
    input n53069;
    input n52513;
    input n12;
    input n8;
    output n52434;
    output n25346;
    output n52939;
    output n52741;
    input n25699;
    input n204;
    output n6;
    input n152;
    output n60212;
    input n53113;
    output n53125;
    output n52496;
    output n25734;
    output n10_adj_12;
    output n25750;
    output n35727;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input n62688;
    input n62430;
    input [23:0]pwm_setpoint;
    input n52427;
    input n62840;
    output [2:0]r_SM_Main;
    output [8:0]r_Clock_Count;
    output tx_o;
    input n26943;
    input \tx_data[2] ;
    output n23;
    output \o_Rx_DV_N_3464[12] ;
    input n4858;
    output \o_Rx_DV_N_3464[24] ;
    output n27;
    output n29;
    output n6_adj_13;
    output tx_enable;
    input n27247;
    input [31:0]baudrate;
    output n55830;
    input n27246;
    input n27245;
    input n27243;
    input n27242;
    output \o_Rx_DV_N_3464[8] ;
    input n4855;
    input n52352;
    output \r_SM_Main[1]_adj_14 ;
    output n25039;
    input n27241;
    input n27240;
    output \r_SM_Main[2]_adj_15 ;
    output n55782;
    output [7:0]r_Clock_Count_adj_24;
    output n55798;
    output n55750;
    output n55766;
    output r_Rx_Data;
    input RX_N_2;
    output n22878;
    output \o_Rx_DV_N_3464[7] ;
    output \o_Rx_DV_N_3464[6] ;
    output \o_Rx_DV_N_3464[5] ;
    output \o_Rx_DV_N_3464[4] ;
    output \o_Rx_DV_N_3464[3] ;
    output \o_Rx_DV_N_3464[2] ;
    output \o_Rx_DV_N_3464[1] ;
    output \o_Rx_DV_N_3464[0] ;
    output n25264;
    input n27583;
    input n48661;
    input n27579;
    output \r_Bit_Index[0] ;
    output n53350;
    output n55734;
    output n55846;
    output n55814;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.i_31__N_2483 , n59174;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n4_c, n4_adj_5254, n61019, n59363, n62679, n26947, n26950, 
        n59173, n2, n2_adj_5255, n2_adj_5256, n2_adj_5257, n59172, 
        n38421;
    wire [2:0]r_SM_Main_2__N_3521;
    
    wire n37879, n59171, n1, n59217, n5, n26, n59170;
    wire [31:0]\FRAME_MATCHER.state_31__N_2588 ;
    
    wire n2_adj_5258, n59169, n2_adj_5259, n2_adj_5260, n59168, n59167, 
        n25674, n2_adj_5261, n2_adj_5262, n2_adj_5263, n2_adj_5264, 
        n2_adj_5265, n2_adj_5266, n2_adj_5267, n2_adj_5268, n2_adj_5269, 
        n26965;
    wire [7:0]\data_in_frame[13]_c ;   // verilog/coms.v(99[12:25])
    
    wire n26987, n62490, n7;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n61017, n59337, n62673, n62484, n7_adj_5270, n26990, n26993, 
        n26996, n26999, n27005, n27011, n62574, n2_adj_5271, n2_adj_5272, 
        n2_adj_5273, n2_adj_5274, n2_adj_5275, n2_adj_5276, n2_adj_5277, 
        n2_adj_5278, n2_adj_5279, n2_adj_5280, n2_adj_5281, n2_adj_5282, 
        n2_adj_5283, n2_adj_5284, n60999, n59336, n62661, n14, n7_adj_5285, 
        n27024, n62655, n2_adj_5286, n62544, n62460, n62649, n62652, 
        n4_adj_5287, n13_c, n62643, n27029, n59216, n59215, n56617, 
        n2173, n27032, n27035;
    wire [23:0]n4757;
    
    wire n25059, n27189;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    
    wire n27063, n27066, n27069, n27072, n27075, n161, n27171, 
        n27167, n27164, n52332, n45647, n52326, n52333, n45646, 
        n52334, n45645, n52331, n45644, n52330, n45643, n52329, 
        n45642, n27160, n27157, n52328, n45641, n52327, tx_transmit_N_3392, 
        n27154;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n23706, n51701;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n26921, n8_c, n7_adj_5288, n9_c, n27142;
    wire [7:0]\data_in_frame[16]_c ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5289, n1_adj_5290, n9_adj_5291, n25, n52472, n27260, 
        n27263, n27266, n51825, n51823, n27275, n27281;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    
    wire n27284, n27287, n27291, n27294, n27297, n27125, n27300, 
        n27303, n51693;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(99[12:25])
    
    wire n51805;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    
    wire n26758, n51691, n51695, n27394;
    wire [7:0]\data_in_frame[18]_c ;   // verilog/coms.v(99[12:25])
    
    wire n27734;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n27731, n52689, n27728, n27725, n27722, n27719, n27716, 
        n27713, n27710;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n27707, n27704, n27701, n27698, n27695, n27692, n27098, 
        n27689, n27686;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    
    wire n27683, n27680, n27677, n51803, n27671, n27668, n27665, 
        n52463, Kp_23__N_724, n26761, n26764, n27636, n27635, n27634, 
        n27633, n27632, n23149, n27060, n27631, n27630, n27629, 
        n27628, n27627, n27626, n27625, n27624, n27623, n27622, 
        n27621, n27620, n27619, n27027, n27618, n27617, n27616, 
        n27615, n27610, n27596, n51791, n51797, n27569, n25455, 
        n46136, n25453, n46135, n25451, n46134, n26776, n52611, 
        n25449, n46133, n52561, n26779, n62631, n26783;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n26788, n26791, n26794, n56626;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n62625, n62628, n62619, n62622, n25447, n46132, n62613, 
        n62616, n62607, n62610, n25445, n46131, n25443, n46130, 
        n25441, n46129, n25439, n46128, n59183, n10_c, n2_adj_5292, 
        n2_adj_5293, n2_adj_5294, n2_adj_5295, n2_adj_5296, n2_adj_5297, 
        n2_adj_5298, n2_adj_5299, n2_adj_5300, n2_adj_5301, n2_adj_5302, 
        n26945;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n26919, n26918, n26917, n2_adj_5303, n25437, n46127, n59187, 
        n2_adj_5305, n2_adj_5306, n2_adj_5307, n2_adj_5308, n2_adj_5309, 
        n2_adj_5310, n2_adj_5311, n2_adj_5312, n2_adj_5313, n2_adj_5314, 
        n2_adj_5315, n2_adj_5316, n2_adj_5317, n2_adj_5318, n2_adj_5319, 
        n2_adj_5320, n2_adj_5321, n2_adj_5322, n6_c, n2_adj_5323, 
        n2_adj_5324, n2_adj_5325, n2_adj_5326, n2_adj_5327, n26798, 
        n26801, n26804, n26807, n26810, n26813, n26816, n26819;
    wire [7:0]\data_in_frame[8]_c ;   // verilog/coms.v(99[12:25])
    
    wire n26822, n26825, n26828, n26831, n26834, n26837, n25685, 
        n25435, n46126, n59188, n55166, n25433, n46125, n59189, 
        n25384, n62844, n25431, n46124, n59280, n25429, n46123, 
        n59281, n62583, n62577, n62580, n25427, n46122, n59282, 
        n24380, \FRAME_MATCHER.i_31__N_2484 , n2153, n2154, n18397, 
        \FRAME_MATCHER.i_31__N_2487 , n51443, \FRAME_MATCHER.i_31__N_2488 , 
        n2165, \FRAME_MATCHER.i_31__N_2489 , n24602, \FRAME_MATCHER.i_31__N_2490 , 
        n37, n23_c, n62571, n25425, n46121, n59283, n25423, n46120, 
        n59284, n25421, n46119, n59286, n25419, n46118, n59287, 
        n25417, n46117, n59288, n62559, n62562, n62553, n62556, 
        n62547, n62550, n62541, n62529, n22, n2_adj_5328, n2_adj_5329, 
        n2_adj_5330, n2_adj_5331, n20, n24145, n26_adj_5332, n2_adj_5333, 
        n2_adj_5334, n2_adj_5335, n2_adj_5336, n2_adj_5337, n2_adj_5338, 
        n2_adj_5339, n2_adj_5340, n2_adj_5341, n25415, n46116, n59289, 
        n2_adj_5342, n52473, n23676, n2_adj_5343, n2_adj_5344, n2_adj_5345, 
        n2_adj_5346, n2_adj_5347, n2_adj_5348, n2_adj_5349, n2_adj_5350, 
        n62454, n59383, n62523, n25413, n46115, n59290, n62442, 
        n61187, n62517, n2_adj_5351, n2_adj_5352, n2_adj_5353, n2_adj_5354, 
        n2_adj_5355, n2_adj_5356, n2_adj_5357, n2_adj_5358, n2_adj_5359, 
        n2_adj_5360, n2_adj_5361, n2_adj_5362, n2_adj_5363, n2_adj_5364, 
        n2_adj_5365, n2_adj_5366, n2_adj_5367, n2_adj_5368, n2_adj_5369, 
        n2_adj_5370, n2_adj_5371, n2_adj_5372, n2_adj_5373, n2_adj_5374, 
        n2_adj_5375, n2_adj_5376, n2_adj_5377, n2_adj_5378, n2_adj_5379, 
        n2_adj_5380, n2_adj_5381, n2_adj_5382, n2_adj_5383, n2_adj_5384, 
        n2_adj_5385, n2_adj_5386, n2_adj_5387, n25411, n46114, n59291, 
        n2_adj_5388, n2_adj_5389, n2_adj_5390, n2_adj_5391, n2_adj_5392, 
        n2_adj_5393, n2_adj_5394, n2_adj_5395, n2_adj_5396, n2_adj_5397, 
        n2_adj_5398, n2_adj_5399, n2_adj_5400, n55133, n47424, n54509, 
        n47264, n47882, n12_c, n22497, n23500, n54710, n52988, 
        n2_adj_5401, n2_adj_5402, n2_adj_5403, n2_adj_5404, n2_adj_5405, 
        n54639, n53049, n6_adj_5406, n2_adj_5407, n2_adj_5408, n2_adj_5409, 
        n52668, n22606, n12_adj_5410, n52883, n54729, n52695, n53014, 
        n55049, n52813, Kp_23__N_1595, n53029, n10_adj_5411, n2_adj_5412, 
        n2_adj_5413, n54169, n52828, n48593, n48509, n4_adj_5414, 
        n52752, n47491, n47458, n54113, n53134, n2_adj_5415, n52868, 
        n52954, n53146, n52875, n16_c, n53170, n23115, n17, n52857, 
        n23821, n18, n14_adj_5416, n2_adj_5417, n52532, n52785, 
        n48458, n15_adj_5418, n52678, n23797, n23318, n6_adj_5419, 
        n23052, n52548, n6_adj_5420, n23294, n23107, n23639, n52969, 
        n12_adj_5421, n3_c, n52343, n47558, n54272, n48503, Kp_23__N_1247, 
        n10_adj_5422, n23313, n52735, n53072, n54381, n52819, n52942, 
        n29_c, n52617, n21, n34, n32_c, n52816, n52801, n52845, 
        n33, n53164, n31, n6_adj_5424;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(99[12:25])
    
    wire n23199, n53058, n52804, n52788, n24073, n3_adj_5425, n52344, 
        n3_adj_5426, n52345, n52725, n3_adj_5427, n52346, n25409, 
        n46113, n59293, n3_adj_5428, n52342, n3_adj_5429, n52339, 
        n3_adj_5430, n52337, n3_adj_5431, n52347, n3_adj_5432, n52348, 
        n3_adj_5433, n52349, n10_adj_5434, n3_adj_5435, n52350, n14_adj_5436, 
        n26797, n3_adj_5437, n52336, n3_adj_5438, n52340, n23135, 
        n52749, n25407, n46112, n59294, n12_adj_5439, n3_adj_5440, 
        n52341, n25405, n46111, n59298, n52972, n52692, n54985, 
        n23283, n53064, n3_adj_5441, n52338, n3_adj_5442, n52351, 
        n1_adj_5443, n1_adj_5444, n1_adj_5445, n2_adj_5446, n2_adj_5447, 
        n2_adj_5448, n1_adj_5449, n2_adj_5450, n1_adj_5451, n1_adj_5452, 
        n1_adj_5453, n2_adj_5454, n2_adj_5455, n2_adj_5456, n2_adj_5457, 
        n2_adj_5458, n2_adj_5459, n2_adj_5460, n2_adj_5461, n1_adj_5462, 
        n26205, n5_adj_5463, n26204, n2_adj_5464, n52834, n6_adj_5465, 
        n24257, n26200, n14_adj_5466, n10_adj_5467, n1_adj_5468, n25403, 
        n46110, n59299, n62511, n62514, n62505, n62508, n25401, 
        n46109, n59300, n25395, n2_adj_5469, n2_adj_5470, n2_adj_5471, 
        n2_adj_5472, n2_adj_5473, n2_adj_5474, n2_adj_5475, n2_adj_5476, 
        n2_adj_5477, n2_adj_5478, n2_adj_5479, n2_adj_5480, n2_adj_5481, 
        n2_adj_5482, n2_adj_5483, n2_adj_5484, n2_adj_5485, n2_adj_5486, 
        n2_adj_5487, n2_adj_5488, n25397, n25399, n26840, n26843, 
        n27428, n27427, n27426, n27425, n27424, n27423, n27422, 
        n27421;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n27420, n27419, n27418, n27417, n27416, n27415, n27414, 
        n27413;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n27412, n27411, n27410, n27409, n27408, n27407, n27406, 
        n27405;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n27404, n27403, n27402, n27401, n27400, n27399, n27398, 
        n26846, n26849, n26852, n26855, n26858, n26861, n26864, 
        n26867, n51689, n51685, n26876, n26879, n26906, n26909, 
        n26912, n47517, n48465, n10_adj_5489, n48650, n52659, n6_adj_5490, 
        n2_adj_5491, n23367, n47444, n46108, n59301, n46107, n59302, 
        n46106, n59303, n2_adj_5492, n2_adj_5493, n51777, n2_adj_5494, 
        n2_adj_5495;
    wire [31:0]n133;
    
    wire n4_adj_5496, n54734, Kp_23__N_950, n26937, n26940, n2_adj_5497, 
        n52577, n52510, n6_adj_5499, n14_adj_5500, n53061, n15_adj_5501, 
        n48450, n23518, n23627, n47579, n6_adj_5502, n52889, n52738, 
        n48127, n48370, n47487, n24165, n23234, n52653, n52982, 
        n52469, n12_adj_5503, n53131, n48439, n6_adj_5504, n47475, 
        n53152, n52662, n15_adj_5505, n8_adj_5506, n52906, n14_adj_5507, 
        n52541, n52900, n52985, n52997, n22_adj_5508, n53155, n24, 
        n20_adj_5510, n52629, n47797, n14_adj_5511, n23607, n13_adj_5512, 
        n6_adj_5513, n52438, n52886, n48578, n2059, n2056, n2062, 
        n54168, n52671, n52702, n24017, n31_adj_5514, n52909, n10_adj_5515, 
        n21154, n52916, n28, n23091, n32_adj_5516, n52903, n53000, 
        n52526, n30, n23670, n31_adj_5517, n52623, n29_adj_5518, 
        n52443, n6_adj_5519, n23750, n23251, n54753, n23763, n23680, 
        n52839, n10_adj_5520, n24061, n53017, n10_adj_5521, n3303, 
        n2110, n22848, n23993, n53020, n23673, n52595, n22929, 
        n5_adj_5522, n6_adj_5523, n52492, n23220, n52871, n23_adj_5524, 
        n25675, n52506, n23238, n10_adj_5525, n23812, n52592, n23269, 
        n6_adj_5526, n52466, Kp_23__N_1037, n53089, n771, n56449, 
        n52635, n23534, n12_adj_5528, n14_adj_5530, n4452, n2125, 
        n7_adj_5531, n10_adj_5532, n6_adj_5533, n53116, n5_adj_5534, 
        n12_adj_5536, n59358, n62478, n61049, n56646, n25461, n56647, 
        n56645, n56843, n12_adj_5537, n56844, n52755, n10_adj_5538, 
        n52846, n56583, n56582, n54791, n7_adj_5539, n56282, n56640, 
        n56641, n52770, n54763, n56594, n56595, n62499, n54087, 
        n56639, n54247, n56367, n59368, n55172, n4_adj_5540, n62700, 
        n62436, n61175, n56603, n56604, n54019, n56823, n56822, 
        n12_adj_5541, n52791, n8_adj_5542, n6_adj_5543, n54630, n10_adj_5544, 
        n54968, n56702, n54614, n56703, n16_adj_5545, n56700, n56699, 
        n56708, n56709, n14_adj_5546, n56670, n56669, n56339, n56711, 
        n13_adj_5547, n56712, n56652, n56651, n56726, n56727, n52948, 
        n15_adj_5548, n14_adj_5549, n54671, n10_adj_5550, n14_adj_5551, 
        n55189, n16_adj_5552, n56365, n18_adj_5553, LED_N_3384, n8_adj_5554, 
        n25012, n10_adj_5555, n34_adj_5556, n23_adj_5557, n22_adj_5558, 
        n35699, n38, n36, n37_adj_5559, n35, n54637, n2122, n52458, 
        n25721, n8_adj_5561, n4_adj_5562, n24203, n1655, n1510, 
        n53052, n52862, n52894, n23577, n52913, n52484, n52475, 
        n52567, n53083, n52587, n10_adj_5563, n52604, n23964, n53043, 
        n53175, n24120, n47422, n54100, n10_adj_5564, n52851, n17_adj_5565, 
        n23005, n1312, n52951, n6_adj_5566, n23601, n53024, n47581, 
        n23155, n48240, n52705, n52520, n10_adj_5567, n52892, n4_adj_5568, 
        n21050, n10_adj_5569, n23568, n52776, n48527, n2054, n48568, 
        n53036, n23185, n52627, n52991, n54349, n52601, n47527, 
        n47720, n52807, n11_adj_5570, n52598, n52860, n54449, n21097, 
        n54473, n53046, n48247, n52632, n52478, n52716, n23713, 
        n48629, n48474, n52764, n48523, n10_adj_5571, n2394, n52552, 
        n10_adj_5572, n1720, n6_adj_5573, n1168, n23869, n10_adj_5574, 
        n24097, n52523, n53040, n48601, n24628, n23_adj_5575, n30909, 
        n6_adj_5576, n25336, n56631, n56632, n56630, n62412, n52529, 
        n23041, n44537, n52489, n23012, n23_adj_5578, n7_adj_5579, 
        n7_adj_5580, n56635, n56633, n62162, n7_adj_5581, n30913, 
        n52674, n47944, n48452, n33540, n14_adj_5582, n4_adj_5583, 
        n8_adj_5584, n48611, n48499, n62493, n52712, n48587, n53078, 
        n48469, n62496, n48494, n48603, n52957, n52683, n6_adj_5585, 
        n52665, n48441, n53143, n2342, n54351, n53023, n53104, 
        n12_adj_5586, n53167, n52761, n47428, n52825, n14_adj_5587, 
        n53149, n6_adj_5588, n14_adj_5589, n53107, n15_adj_5590, n8_adj_5591, 
        n48471, n53003, n62487, n52810, n22527, n21093, n52686, 
        n53011, n10_adj_5594, n23699, n7_adj_5595, n48525, n52403, 
        n47856, n2217, n52932, n52854, n13_adj_5596, n52808, n47968, 
        n16_adj_5597, n52709, n17_adj_5598, n53101, n48463, n23967, 
        n23455, n10_adj_5599, n52721, n52935, n62481, n52758, n16_adj_5600, 
        n17_adj_5601, n54016, n52864, n62166, n24_adj_5602, n23754, 
        n26_adj_5603, n52794, n25_adj_5604, n27_c, n6_adj_5605, n53026, 
        n1699, n52481, n53075, n52773, n1835, n10_adj_5606, n47641, 
        n52452, n1673, n18_adj_5607, n52614, n19, n22437, n10_adj_5608, 
        n52779, n23437, n14_adj_5609, n52822, n14_adj_5610, n52555, 
        n6_adj_5611, n55042, n54735, n28_adj_5612, n26_adj_5613, n27_adj_5614, 
        n53008, n25_adj_5615, n2329, n55052, n8_adj_5616, n48308, 
        n6_adj_5617, n47456, n53032, n6_adj_5618, n52966, n16_adj_5619, 
        n17_adj_5620, n23613, n10_adj_5621, n47502, n53158, n52963, 
        n59351, n23263, n56634, n52897, n12_adj_5622, n23758, n24002, 
        n26_adj_5623, n52647, n24_adj_5624, n25_adj_5625, n54139, 
        n23434, n12_adj_5626, n54459, n12_adj_5627, n47414, n52500, 
        n53119, n10_adj_5630, n53110, n10_adj_5631, n1191, n62475, 
        n23410, n53128, n52975, n52919, n12_adj_5633, n52446, n28_adj_5634, 
        n38_adj_5635, n36_adj_5636, n42, n40, n41, n39, n10_adj_5637, 
        n12_adj_5638, n52746, n12_adj_5639, n62457, n62451, n62445, 
        n54683, n2113, n2060, n22768, n20118, n24375, n4_adj_5641, 
        n24379, n62439, n10_adj_5642, n14_adj_5643, n22932, n20_adj_5644, 
        n22787, n19_adj_5645, n56471, n22884, n18_adj_5646, n22867, 
        n20_adj_5647, n15_adj_5648, n16_adj_5649, n17_adj_5650, n10_adj_5651, 
        n14_adj_5652, n15_adj_5653, n16_adj_5654, n17_adj_5655, n6_adj_5656, 
        n62433, n62697, n62691, n62409;
    wire [2:0]r_SM_Main_2__N_3512;
    
    wire n53934;
    
    SB_LUT4 i44591_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59174));   // verilog/coms.v(158[12:15])
    defparam i44591_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(\byte_transmit_counter[4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[1] ), 
            .O(n4_adj_5254));
    defparam i1_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47739 (.I0(\byte_transmit_counter[3] ), 
            .I1(n61019), .I2(n59363), .I3(\byte_transmit_counter[4] ), 
            .O(n62679));
    defparam byte_transmit_counter_3__bdd_4_lut_47739.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n26947));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n26950));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i44590_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59173));   // verilog/coms.v(158[12:15])
    defparam i44590_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2), .S(n52280));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5255), .S(n52279));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5256), .S(n52310));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5257), .S(n52278));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i44587_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59172));   // verilog/coms.v(158[12:15])
    defparam i44587_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24826_4_lut (.I0(\byte_transmit_counter[3] ), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_5254), .I3(n4_c), .O(n38421));
    defparam i24826_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i24291_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3521[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37879));
    defparam i24291_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n26953));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i44586_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59171));   // verilog/coms.v(158[12:15])
    defparam i44586_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44766_2_lut (.I0(\data_out_frame[3][3] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n59217));
    defparam i44766_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n26));   // verilog/coms.v(105[12:33])
    defparam i46_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44585_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59170));   // verilog/coms.v(158[12:15])
    defparam i44585_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5258));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44582_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59169));   // verilog/coms.v(158[12:15])
    defparam i44582_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5259), .S(n52309));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5260), .S(n52308));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5259));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44808_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59168));   // verilog/coms.v(158[12:15])
    defparam i44808_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44859_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59167));   // verilog/coms.v(158[12:15])
    defparam i44859_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11968_1_lut (.I0(n3543), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25674));   // verilog/coms.v(148[4] 304[11])
    defparam i11968_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5261), .S(n52307));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5262), .S(n52306));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n26957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5263), .S(n26691));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5264), .S(n52154));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5265), .S(n52305));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n26960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5266), .S(n52304));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5267), .S(n52318));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5268), .S(n52303));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5269), .S(n52158));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13]_c [3]), .C(clk16MHz), 
           .D(n26965));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13][4] ), .C(clk16MHz), 
           .D(n26969));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13][5] ), .C(clk16MHz), 
           .D(n26972));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27218));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13][6] ), .C(clk16MHz), 
           .D(n26979));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13][7] ), .C(clk16MHz), 
           .D(n26982));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27213));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n26987));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n62679_bdd_4_lut (.I0(n62679), .I1(n62490), .I2(n7), .I3(\byte_transmit_counter[4] ), 
            .O(tx_data[6]));
    defparam n62679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47729 (.I0(\byte_transmit_counter[3] ), 
            .I1(n61017), .I2(n59337), .I3(\byte_transmit_counter[4] ), 
            .O(n62673));
    defparam byte_transmit_counter_3__bdd_4_lut_47729.LUT_INIT = 16'he4aa;
    SB_LUT4 n62673_bdd_4_lut (.I0(n62673), .I1(n62484), .I2(n7_adj_5270), 
            .I3(\byte_transmit_counter[4] ), .O(tx_data[7]));
    defparam n62673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n26990));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n26993));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
           .D(n26996));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n26999));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n27005));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27203));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27200));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n27011));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_775_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5257));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45078_2_lut (.I0(n62574), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59363));
    defparam i45078_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5256));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5271));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5272));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5273));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5274));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5275));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5276));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5277));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5278));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5279));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5280));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5281));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5282));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5283));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5284));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1129 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[10] [2]), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5255));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1129.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47719 (.I0(\byte_transmit_counter[3] ), 
            .I1(n60999), .I2(n59336), .I3(\byte_transmit_counter[4] ), 
            .O(n62661));
    defparam byte_transmit_counter_3__bdd_4_lut_47719.LUT_INIT = 16'he4aa;
    SB_LUT4 n62661_bdd_4_lut (.I0(n62661), .I1(n14), .I2(n7_adj_5285), 
            .I3(\byte_transmit_counter[4] ), .O(tx_data[1]));
    defparam n62661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n27024));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47734 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n62655));
    defparam byte_transmit_counter_0__bdd_4_lut_47734.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5286), .S(n52156));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n62655_bdd_4_lut (.I0(n62655), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n62658));
    defparam n62655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46119_3_lut (.I0(n62544), .I1(n62460), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n61019));
    defparam i46119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47709 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n62649));
    defparam byte_transmit_counter_0__bdd_4_lut_47709.LUT_INIT = 16'he4aa;
    SB_LUT4 n62649_bdd_4_lut (.I0(n62649), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n62652));
    defparam n62649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n4_adj_5287), .I2(n13_c), .I3(\byte_transmit_counter[2] ), 
            .O(n62643));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n27029));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n62643_bdd_4_lut (.I0(n62643), .I1(n59216), .I2(n59215), .I3(\byte_transmit_counter[2] ), 
            .O(n56617));
    defparam n62643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1724), .C(clk16MHz), 
            .D(n2173), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n27032));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n27035));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27192));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n25059), 
            .D(n4757[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27189));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n27063));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n27066));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n27069));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5284), .S(n52277));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5283), .S(n52276));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5282), .S(n52275));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5281), .S(n52274));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5280), .S(n52273));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5279), .S(n52272));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5278), .S(n52271));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5277), .S(n52270));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5276), .S(n52269));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5275), .S(n52268));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5274), .S(n52267));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5273), .S(n52266));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5272), .S(n52265));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5271), .S(n52264));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n27072));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n27075));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n35706));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'hbbbb;
    SB_DFFE data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27171));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n27101));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27167));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27164));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1082_9_lut (.I0(n52326), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n45647), .O(n52332)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1082_8_lut (.I0(n52326), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n45646), .O(n52333)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1082_8 (.CI(n45646), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n45647));
    SB_LUT4 add_1082_7_lut (.I0(n52326), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n45645), .O(n52334)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1082_7 (.CI(n45645), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n45646));
    SB_LUT4 add_1082_6_lut (.I0(n52326), .I1(\byte_transmit_counter[4] ), 
            .I2(GND_net), .I3(n45644), .O(n52331)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1082_6 (.CI(n45644), .I0(\byte_transmit_counter[4] ), .I1(GND_net), 
            .CO(n45645));
    SB_LUT4 add_1082_5_lut (.I0(n52326), .I1(\byte_transmit_counter[3] ), 
            .I2(GND_net), .I3(n45643), .O(n52330)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n27105));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1082_5 (.CI(n45643), .I0(\byte_transmit_counter[3] ), .I1(GND_net), 
            .CO(n45644));
    SB_LUT4 add_1082_4_lut (.I0(n52326), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n45642), .O(n52329)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_4_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27160));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27157));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1082_4 (.CI(n45642), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n45643));
    SB_LUT4 add_1082_3_lut (.I0(n52326), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n45641), .O(n52328)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1082_3 (.CI(n45641), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n45642));
    SB_LUT4 add_1082_2_lut (.I0(n52326), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3392), .I3(GND_net), .O(n52327)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1082_2_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27154));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n23706));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n51701));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i21438_3_lut_4_lut (.I0(\Kp[5] ), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26921));
    defparam i21438_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_1082_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3392), .CO(n45641));
    SB_DFFE data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27148));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n27130));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[1]), .I3(ID[5]), .O(n8_c));
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1131 (.I0(ID[7]), .I1(\data_in_frame[0] [2]), .I2(\data_in_frame[0][7] ), 
            .I3(ID[2]), .O(n7_adj_5288));
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'h7bde;
    SB_DFFE data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27144));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n27133));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut (.I0(ID[6]), .I1(ID[3]), .I2(\data_in_frame[0] [6]), 
            .I3(\data_in_frame[0] [3]), .O(n9_c));
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_DFFE data_in_frame_0___i134 (.Q(\data_in_frame[16]_c [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27142));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5289), .S(n52263));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(n9_c), .I1(n7_adj_5288), .I2(n8_c), .I3(GND_net), 
            .O(n1_adj_5290));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1132 (.I0(\data_in_frame[0] [0]), .I1(ID[4]), .I2(ID[0]), 
            .I3(\data_in_frame[0] [4]), .O(n9_adj_5291));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1132.LUT_INIT = 16'h7bde;
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16][4] ), .C(clk16MHz), 
           .D(n27136));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1133 (.I0(n9_adj_5291), .I1(n1_adj_5290), .I2(GND_net), 
            .I3(GND_net), .O(n25));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52472));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n27129), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n27128), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n27127), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n27126), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n26731));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n26734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n26737));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n26740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n27260));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n27263));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n27266));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n51825));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n51823));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n27275));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0][7] ), .C(clk16MHz), 
           .D(n51817));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
           .D(n27281));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
           .D(n27284));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
           .D(n27287));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
           .D(n27291));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n27294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n27297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27772));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n27125), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n27124), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n27123), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n27122), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n27121), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n27120), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n26743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n27300));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n27303));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n51681));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n51677));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n27312));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n27317));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n51673));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n27321));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2]_c [6]), .C(clk16MHz), 
           .D(n51693));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n26746));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n26749));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2][7] ), .C(clk16MHz), 
           .D(n27327));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
           .D(n27331));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n27757));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n51805));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6][1] ), .C(clk16MHz), 
           .D(n26758));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3][1] ), .C(clk16MHz), 
           .D(n51669));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
           .D(n51667));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n51663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3][4] ), .C(clk16MHz), 
           .D(n51659));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n27119), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n27118), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n27117), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n27116), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n27115), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n27114), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n27113), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n27112), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n27111), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n27110), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n51691));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
           .D(n51695));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3][7] ), .C(clk16MHz), 
           .D(n51655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n27365));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n27370));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n27375));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n27379));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n27387));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n27391));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18]_c [6]), .C(clk16MHz), 
           .D(n27394));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18][7] ), .C(clk16MHz), 
           .D(n27430));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n27433));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n51579));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n27439));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27734));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27731));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52689));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n27109), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n27108), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27728));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27725));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27722));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27719));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27716));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27713));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27710));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n27104), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27707));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27704));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27701));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27698));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27695));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27692));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n27100));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n27099));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n27098));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n27097));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n27096));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27689));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27686));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27683));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27680));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27677));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n27095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n27094));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n27093));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n27092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n27091));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n51803));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27671));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27668));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27665));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27662));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27659));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i20953_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n20140), .I3(GND_net), .O(n27098));
    defparam i20953_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n27090));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n27089));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n27088));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1136 (.I0(\data_in_frame[0][7] ), .I1(n52689), 
            .I2(n52472), .I3(n52463), .O(Kp_23__N_724));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n27087));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n27086));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n27085));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n27084));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n27083));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n27082));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n27081));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n27080));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27656));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27653));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27650));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27647));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27644));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n27079));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n27078));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n51577));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n51575));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6][2] ), .C(clk16MHz), 
           .D(n26761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6][3] ), .C(clk16MHz), 
           .D(n26764));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27637));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n27636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n27635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n27634));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n27633));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n27632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n27062), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1137 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n23149));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n27061), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n27060), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n27056));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n27055), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n27054), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n27053), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n27052), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n27631));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n27630));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n27629));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n27628));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n27627));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n27051), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n27050), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n27049), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n27048), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n27047), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n27046), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n27045), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n27044), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n27043), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n27042), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n27041), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n27040), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n27039), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n27038), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n27626));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n27625));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n27624));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n27623));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n27622));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n27621));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n27620));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n27619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n27028), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n27027), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n27618));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n27617));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n27616));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n27615));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n27614), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n27613), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n27612), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n27611), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n27610), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n27609), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n27608), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n27023), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n27022), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n27021), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n27020), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n27019), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n27018), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n27607), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n27606), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n27605), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n27604), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n27603), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n27602), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n27601), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n27600), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n27599), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n27598), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n27017), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n27016), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n27597), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n27596), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n27595), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n27594), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n27593), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27590));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6][4] ), .C(clk16MHz), 
           .D(n51791));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n27015), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
           .D(n51797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27569));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n27014), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n27010), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_33_lut  (.I0(n59167), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n46136), .O(n25455)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_32_lut  (.I0(n59168), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n46135), .O(n25453)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_32  (.CI(n46135), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n46136));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_31_lut  (.I0(n59169), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n46134), .O(n25451)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_31  (.CI(n46134), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n46135));
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6][6] ), .C(clk16MHz), 
           .D(n26776));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52463));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5258), .S(n52302));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_724), 
            .I2(GND_net), .I3(GND_net), .O(n52611));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n26986), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n26985), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_30_lut  (.I0(n59170), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n46133), .O(n25449)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_1044_i23_3_lut_4_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i23_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52561));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6][7] ), .C(clk16MHz), 
           .D(n26779));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47699 (.I0(\byte_transmit_counter[1] ), 
            .I1(n26), .I2(n5), .I3(\byte_transmit_counter[2] ), .O(n62631));
    defparam byte_transmit_counter_1__bdd_4_lut_47699.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n26783));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n51567));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n26788));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n26791));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n26794));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n51549));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27551));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n26978), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n62631_bdd_4_lut (.I0(n62631), .I1(n59217), .I2(n1), .I3(\byte_transmit_counter[2] ), 
            .O(n56626));
    defparam n62631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_30  (.CI(n46133), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n46134));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47704 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n62625));
    defparam byte_transmit_counter_0__bdd_4_lut_47704.LUT_INIT = 16'he4aa;
    SB_LUT4 n62625_bdd_4_lut (.I0(n62625), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n62628));
    defparam n62625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47684 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n62619));
    defparam byte_transmit_counter_0__bdd_4_lut_47684.LUT_INIT = 16'he4aa;
    SB_LUT4 n62619_bdd_4_lut (.I0(n62619), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n62622));
    defparam n62619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_29_lut  (.I0(n59171), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n46132), .O(n25447)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47679 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n62613));
    defparam byte_transmit_counter_0__bdd_4_lut_47679.LUT_INIT = 16'he4aa;
    SB_LUT4 n62613_bdd_4_lut (.I0(n62613), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n62616));
    defparam n62613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47674 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n62607));
    defparam byte_transmit_counter_0__bdd_4_lut_47674.LUT_INIT = 16'he4aa;
    SB_LUT4 n62607_bdd_4_lut (.I0(n62607), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n62610));
    defparam n62607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_29  (.CI(n46132), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n46133));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_28_lut  (.I0(n59172), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n46131), .O(n25445)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n26977), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n25059), 
            .D(n4757[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_28  (.CI(n46131), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n46132));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_27_lut  (.I0(n59173), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n46130), .O(n25443)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n26976), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_27  (.CI(n46130), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n46131));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_26_lut  (.I0(n59174), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n46129), .O(n25441)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_26  (.CI(n46129), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n46130));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_25_lut  (.I0(n59183), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n46128), .O(n25439)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 equal_1925_i10_2_lut (.I0(\data_in_frame[0][7] ), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // verilog/coms.v(169[9:87])
    defparam equal_1925_i10_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5292), .S(n26705));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5293), .S(n52317));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5294), .S(n52316));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5295), .S(n52315));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5296), .S(n52314));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5297), .S(n52313));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5298), .S(n52312));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5299), .S(n52311));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5300), .S(n52157));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n26975), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n26968), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n26956), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5301), .S(n52218));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5302), .S(n52301));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n26946), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n26945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n26944), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1044_i22_3_lut_4_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i22_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n26930), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n26929), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n26925), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n26924), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n26921), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n26920), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n26919));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n26918));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n26917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n26916), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n26915), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5303), .S(n52262));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i24178_3_lut (.I0(encoder0_position_scaled[13]), .I1(\motor_state_23__N_67[13] ), 
            .I2(n15), .I3(GND_net), .O(n9));
    defparam i24178_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1044_i21_3_lut_4_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i21_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_25  (.CI(n46128), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n46129));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_24_lut  (.I0(n59187), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n46127), .O(n25437)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5305), .S(n52261));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5306), .S(n52260));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5307), .S(n52259));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5308), .S(n52258));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5309), .S(n52257));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5310), .S(n52256));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5311), .S(n52255));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5312), .S(n52254));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5313), .S(n52160));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5314), .S(n52253));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5315), .S(n52252));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5316), .S(n52251));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5317), .S(n52250));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5318), .S(n52249));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5319), .S(n52248));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5320), .S(n26347));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5321), .S(n52247));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5322), .S(n52246));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1141 (.I0(\data_in_frame[0][7] ), .I1(\data_in_frame[2] [0]), 
            .I2(n52561), .I3(n52611), .O(n6_c));
    defparam i2_4_lut_adj_1141.LUT_INIT = 16'h4812;
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5323), .S(n52217));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5324), .S(n52245));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5325), .S(n52244));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5326), .S(n52243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5327), .S(n52242));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n26798));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n27549), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n26801));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n26804));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1044_i20_3_lut_4_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i20_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n26807));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n26810));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n26813));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_24  (.CI(n46127), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n46128));
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n26816));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8]_c [3]), .C(clk16MHz), 
           .D(n26819));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8][4] ), .C(clk16MHz), 
           .D(n26822));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8][5] ), .C(clk16MHz), 
           .D(n26825));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8][6] ), .C(clk16MHz), 
           .D(n26828));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8][7] ), .C(clk16MHz), 
           .D(n26831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n51565));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n26834));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n26837));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1142 (.I0(\FRAME_MATCHER.i[1] ), .I1(n52409), .I2(\FRAME_MATCHER.i[0] ), 
            .I3(GND_net), .O(n25685));
    defparam i2_3_lut_adj_1142.LUT_INIT = 16'hefef;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n25059), 
            .D(n4757[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n25059), 
            .D(n4757[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n25059), 
            .D(n4757[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n25059), 
            .D(n4757[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n25059), 
            .D(n4757[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n25059), 
            .D(n4757[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n25059), 
            .D(n4757[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n25059), 
            .D(n4757[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n25059), 
            .D(n4757[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n25059), 
            .D(n4757[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n25059), 
            .D(n4757[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n25059), 
            .D(n4757[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n25059), 
            .D(n4757[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n25059), 
            .D(n4757[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n25059), 
            .D(n4757[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n25059), 
            .D(n4757[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n25059), 
            .D(n4757[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n25059), 
            .D(n4757[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n25059), 
            .D(n4757[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n25059), 
            .D(n4757[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n25059), 
            .D(n4757[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n25059), 
            .D(n4757[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1044_i19_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i19_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1044_i18_3_lut_4_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i18_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i21604_3_lut_4_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[16]));
    defparam i21604_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_23_lut  (.I0(n59188), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n46126), .O(n25435)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_23  (.CI(n46126), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n46127));
    SB_LUT4 i3_4_lut_adj_1143 (.I0(n23149), .I1(n6_c), .I2(Kp_23__N_724), 
            .I3(\data_in_frame[2] [1]), .O(n55166));
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h0440;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_22_lut  (.I0(n59189), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n46125), .O(n25433)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_1044_i16_3_lut_4_lut (.I0(\data_in_frame[18][7] ), .I1(\data_in_frame[2][7] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i16_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFFR \FRAME_MATCHER.i_1933__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n25384), .R(reset));   // verilog/coms.v(158[12:15])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_22  (.CI(n46125), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n46126));
    SB_LUT4 i21272_3_lut_4_lut (.I0(\data_in_frame[18]_c [6]), .I1(\data_in_frame[2]_c [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[14]));
    defparam i21272_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2483 ), 
            .C(clk16MHz), .D(n62844), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_21_lut  (.I0(n59280), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n46124), .O(n25431)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_21  (.CI(n46124), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n46125));
    SB_LUT4 mux_1044_i14_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i14_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_20_lut  (.I0(n59281), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n46123), .O(n25429)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_20  (.CI(n46123), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n46124));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47659 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n62583));
    defparam byte_transmit_counter_0__bdd_4_lut_47659.LUT_INIT = 16'he4aa;
    SB_LUT4 n62583_bdd_4_lut (.I0(n62583), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n62586));
    defparam n62583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47650 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n62577));
    defparam byte_transmit_counter_0__bdd_4_lut_47650.LUT_INIT = 16'he4aa;
    SB_LUT4 n62577_bdd_4_lut (.I0(n62577), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n62580));
    defparam n62577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1044_i13_3_lut_4_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i13_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_19_lut  (.I0(n59282), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n46122), .O(n25427)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_19  (.CI(n46122), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n46123));
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2484 ), 
            .C(clk16MHz), .D(n24380), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2485 ), 
            .C(clk16MHz), .D(n2153), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2154), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2487 ), 
            .C(clk16MHz), .D(n18397), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2488 ), 
            .C(clk16MHz), .D(n51443), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2489 ), 
            .C(clk16MHz), .D(n2165), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2490 ), 
            .C(clk16MHz), .D(n24602), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i14007_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n27713));
    defparam i14007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(n25), .O(n23_c));
    defparam i9_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i14010_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n27716));
    defparam i14010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1044_i12_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i12_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47645 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n62571));
    defparam byte_transmit_counter_0__bdd_4_lut_47645.LUT_INIT = 16'he4aa;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_18_lut  (.I0(n59283), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n46121), .O(n25425)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_18  (.CI(n46121), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n46122));
    SB_LUT4 mux_1044_i11_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i11_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 n62571_bdd_4_lut (.I0(n62571), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n62574));
    defparam n62571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14013_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n27719));
    defparam i14013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1044_i10_3_lut_4_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i10_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_17_lut  (.I0(n59284), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n46120), .O(n25423)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_17  (.CI(n46120), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n46121));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_16_lut  (.I0(n59286), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n46119), .O(n25421)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_16  (.CI(n46119), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n46120));
    SB_LUT4 mux_1044_i9_3_lut_4_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i9_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_15_lut  (.I0(n59287), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n46118), .O(n25419)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_15  (.CI(n46118), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n46119));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_14_lut  (.I0(n59288), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n46117), .O(n25417)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47635 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n62559));
    defparam byte_transmit_counter_0__bdd_4_lut_47635.LUT_INIT = 16'he4aa;
    SB_LUT4 n62559_bdd_4_lut (.I0(n62559), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n62562));
    defparam n62559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47630 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n62553));
    defparam byte_transmit_counter_0__bdd_4_lut_47630.LUT_INIT = 16'he4aa;
    SB_LUT4 n62553_bdd_4_lut (.I0(n62553), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n62556));
    defparam n62553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47625 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n62547));
    defparam byte_transmit_counter_0__bdd_4_lut_47625.LUT_INIT = 16'he4aa;
    SB_LUT4 n62547_bdd_4_lut (.I0(n62547), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n62550));
    defparam n62547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47620 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n62541));
    defparam byte_transmit_counter_0__bdd_4_lut_47620.LUT_INIT = 16'he4aa;
    SB_LUT4 n62541_bdd_4_lut (.I0(n62541), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n62544));
    defparam n62541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1044_i8_3_lut_4_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3][7] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[7]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i8_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47615 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n62529));
    defparam byte_transmit_counter_0__bdd_4_lut_47615.LUT_INIT = 16'he4aa;
    SB_LUT4 n62529_bdd_4_lut (.I0(n62529), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n62532));
    defparam n62529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_14  (.CI(n46117), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n46118));
    SB_LUT4 i8_4_lut (.I0(n10_c), .I1(\data_in_frame[1] [2]), .I2(\data_in_frame[1] [5]), 
            .I3(n23706), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h0040;
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5328), .S(n52241));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5329), .S(n52240));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5330), .S(n52239));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5331), .S(n52223));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut (.I0(n23_c), .I1(n55166), .I2(n20), .I3(n24145), 
            .O(n26_adj_5332));
    defparam i12_4_lut.LUT_INIT = 16'h0080;
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5333), .S(n52238));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5334), .S(n52237));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5335), .S(n52236));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5336), .S(n52235));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5337), .S(n52234));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5338), .S(n52233));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5339), .S(n52232));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5340), .S(n52231));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n27935), .D(n2_adj_5341), .S(n26327));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14016_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n27722));
    defparam i14016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_13_lut  (.I0(n59289), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n46116), .O(n25415)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5342), .S(n52230));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13_4_lut (.I0(n52473), .I1(n26_adj_5332), .I2(n22), .I3(n23676), 
            .O(\FRAME_MATCHER.state_31__N_2588 [3]));
    defparam i13_4_lut.LUT_INIT = 16'h0040;
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5343), .S(n52229));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_13  (.CI(n46116), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n46117));
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5344), .S(n52228));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5345), .S(n52227));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5346), .S(n52226));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5347), .S(n52225));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5348), .S(n52155));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5349), .S(n26319));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5350), .S(n52220));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47714 (.I0(\byte_transmit_counter[3] ), 
            .I1(n62454), .I2(n59383), .I3(\byte_transmit_counter[4] ), 
            .O(n62523));
    defparam byte_transmit_counter_3__bdd_4_lut_47714.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1044_i7_3_lut_4_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i7_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1044_i6_3_lut_4_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i6_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_12_lut  (.I0(n59290), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n46115), .O(n25413)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 n62523_bdd_4_lut (.I0(n62523), .I1(n62442), .I2(n56626), .I3(\byte_transmit_counter[4] ), 
            .O(tx_data[3]));
    defparam n62523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_12  (.CI(n46115), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n46116));
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47600 (.I0(\byte_transmit_counter[3] ), 
            .I1(n61187), .I2(n59364), .I3(\byte_transmit_counter[4] ), 
            .O(n62517));
    defparam byte_transmit_counter_3__bdd_4_lut_47600.LUT_INIT = 16'he4aa;
    SB_LUT4 n62517_bdd_4_lut (.I0(n62517), .I1(n62466), .I2(n56617), .I3(\byte_transmit_counter[4] ), 
            .O(tx_data[4]));
    defparam n62517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_775_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n27945), .D(n2_adj_5351), .S(n26317));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5352), .S(n52221));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5353), .S(n52222));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5354), .S(n52224));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5355), .S(n52159));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5356), .S(n52219));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5357), .S(n52161));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5358), .S(n52162));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5359), .S(n52163));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5360), .S(n52164));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5361), .S(n52165));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5362), .S(n52166));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5363), .S(n52167));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5364), .S(n52168));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5365), .S(n52169));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n27960), .D(n2_adj_5366), .S(n26302));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5367), .S(n52170));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n27962), .D(n2_adj_5368), .S(n26300));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5369), .S(n52171));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5370), .S(n52172));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5371), .S(n52173));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5372), .S(n52174));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5373), .S(n52175));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n27968), .D(n2_adj_5374), .S(n26294));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5375), .S(n52176));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n27970), .D(n2_adj_5376), .S(n26292));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5377), .S(n52177));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5378), .S(n52178));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5379), .S(n52179));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5380), .S(n52180));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5381), .S(n52181));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5382), .S(n52182));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5383), .S(n52183));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n27978), .D(n2_adj_5384), .S(n26284));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n27979), .D(n2_adj_5385), .S(n26283));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5386), .S(n52184));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n27981), .D(n2_adj_5387), .S(n26281));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_11_lut  (.I0(n59291), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n46114), .O(n25411)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5388), .S(n52185));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5389), .S(n52186));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5390), .S(n52187));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n27985), .D(n2_adj_5391), .S(n26277));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n27986), .D(n2_adj_5392), .S(n26276));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13688_3_lut (.I0(\data_in_frame[18]_c [6]), .I1(rx_data[6]), 
            .I2(n54720), .I3(GND_net), .O(n27394));   // verilog/coms.v(130[12] 305[6])
    defparam i13688_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n27987), .D(n2_adj_5393), .S(n26275));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5394), .S(n52188));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5395), .S(n52189));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5396), .S(n52190));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5397), .S(n52191));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5398), .S(n52192));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5399), .S(n52193));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5400), .S(n52194));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1144 (.I0(\data_in_frame[18] [0]), .I1(n55133), 
            .I2(n47424), .I3(GND_net), .O(n54509));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut (.I0(n47264), .I1(n54509), .I2(n55133), .I3(n47882), 
            .O(n12_c));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1044_i5_3_lut_4_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3][4] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i5_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i6_4_lut (.I0(n22497), .I1(n12_c), .I2(n23500), .I3(n54710), 
            .O(n52988));
    defparam i6_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5401), .S(n52195));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5402), .S(n52196));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5403), .S(n52197));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1044_i4_3_lut_4_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3][3] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i4_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5404), .S(n52198));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5405), .S(n52199));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1044_i3_3_lut_4_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3][2] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i3_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[17] [5]), .I1(n54639), .I2(n53049), 
            .I3(n6_adj_5406), .O(n47424));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5407), .S(n52200));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5408), .S(n52201));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5409), .S(n52202));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1145 (.I0(\data_in_frame[18]_c [6]), .I1(n52668), 
            .I2(\data_in_frame[21] [0]), .I3(n22606), .O(n12_adj_5410));
    defparam i5_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1146 (.I0(\data_in_frame[18] [4]), .I1(n12_adj_5410), 
            .I2(n52883), .I3(\data_in_frame[18][7] ), .O(n54729));
    defparam i6_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(n54729), .I1(n52695), .I2(GND_net), 
            .I3(GND_net), .O(n53014));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(n55049), .I1(n52813), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1595));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1149 (.I0(\data_in_frame[20] [2]), .I1(n53029), 
            .I2(\data_in_frame[13][4] ), .I3(\data_in_frame[15] [6]), .O(n10_adj_5411));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5412), .S(n52203));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5413), .S(n52204));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[19] [4]), .I1(n54169), .I2(n52828), 
            .I3(GND_net), .O(n48593));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[16] [6]), .I1(n48509), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5414));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1151 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[17] [1]), 
            .I2(n52752), .I3(n4_adj_5414), .O(n52813));
    defparam i2_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(n47491), .I1(n52813), .I2(GND_net), 
            .I3(GND_net), .O(n47458));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1153 (.I0(\data_in_frame[19] [6]), .I1(n54113), 
            .I2(\data_in_frame[20] [1]), .I3(GND_net), .O(n53134));
    defparam i2_3_lut_adj_1153.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5415), .S(n52205));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14019_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n27725));
    defparam i14019_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53049));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1044_i2_3_lut_4_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3][1] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i2_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n52868), .I1(n52954), .I2(n53146), 
            .I3(n52875), .O(n16_c));
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n53049), .I1(n53170), .I2(n23115), .I3(\data_in_frame[16][4] ), 
            .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1156 (.I0(n52857), .I1(n23821), .I2(n17), .I3(n18), 
            .O(n14_adj_5416));
    defparam i5_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5417), .S(n52206));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1157 (.I0(n52532), .I1(\data_in_frame[17] [1]), 
            .I2(n52785), .I3(n48458), .O(n15_adj_5418));
    defparam i6_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1158 (.I0(n15_adj_5418), .I1(\data_in_frame[15] [4]), 
            .I2(n14_adj_5416), .I3(n52678), .O(n55133));
    defparam i8_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(n23797), .I1(n23318), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5419));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[14] [0]), 
            .I2(n23052), .I3(n6_adj_5419), .O(n52548));
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[15] [6]), .I1(n52548), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5420));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(\data_in_frame[13][5] ), .I1(\data_in_frame[13][6] ), 
            .I2(n23294), .I3(n6_adj_5420), .O(n52954));
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1163 (.I0(\data_in_frame[11] [2]), .I1(n23107), 
            .I2(\data_in_frame[8][6] ), .I3(n23639), .O(n53029));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1164 (.I0(n52954), .I1(n52969), .I2(\data_in_frame[16] [1]), 
            .I3(\data_in_frame[16] [0]), .O(n12_adj_5421));
    defparam i5_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i14022_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n27728));
    defparam i14022_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2978), .D(n3_c), .S(n52343));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1165 (.I0(n47558), .I1(n12_adj_5421), .I2(n53029), 
            .I3(\data_in_frame[13] [1]), .O(n54272));
    defparam i6_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1166 (.I0(\data_in_frame[16] [2]), .I1(n52548), 
            .I2(n48503), .I3(Kp_23__N_1247), .O(n10_adj_5422));
    defparam i4_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1167 (.I0(\data_in_frame[14] [2]), .I1(n10_adj_5422), 
            .I2(n23313), .I3(GND_net), .O(n52883));
    defparam i5_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(\data_in_frame[16] [3]), .I1(n52883), 
            .I2(n54272), .I3(GND_net), .O(n47882));
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(n47882), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[18] [4]), .O(n52735));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_in_frame[16] [3]), .I1(n22606), 
            .I2(GND_net), .I3(GND_net), .O(n52532));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1171 (.I0(n53072), .I1(n54381), .I2(\data_in_frame[18] [5]), 
            .I3(n52819), .O(n52942));
    defparam i3_4_lut_adj_1171.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut (.I0(n52735), .I1(n53072), .I2(\data_in_frame[21] [7]), 
            .I3(\data_in_frame[21] [6]), .O(n29_c));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[21] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52617));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut (.I0(n29_c), .I1(n21), .I2(n55133), .I3(\data_in_frame[19] [7]), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1173 (.I0(n53134), .I1(n55049), .I2(n47458), 
            .I3(\data_in_frame[21] [4]), .O(n32_c));
    defparam i13_4_lut_adj_1173.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut (.I0(n52816), .I1(n52801), .I2(n52617), .I3(n52845), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1174 (.I0(n48593), .I1(n53164), .I2(\data_in_frame[21] [1]), 
            .I3(\data_in_frame[17] [7]), .O(n31));
    defparam i12_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33), .I2(n32_c), .I3(n34), .O(n52695));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14025_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n27731));
    defparam i14025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[12] [7]), .I1(n4), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5424));
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1176 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10]_c [5]), 
            .I2(n23199), .I3(n6_adj_5424), .O(n53058));
    defparam i4_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1177 (.I0(\data_in_frame[17] [2]), .I1(n52804), 
            .I2(n53058), .I3(n52788), .O(n53146));
    defparam i1_4_lut_adj_1177.LUT_INIT = 16'h9669;
    SB_LUT4 i14028_3_lut_4_lut (.I0(n37), .I1(n52430), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n27734));
    defparam i14028_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(n23313), .I1(n24073), .I2(GND_net), 
            .I3(GND_net), .O(n52804));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5425), .S(n52344));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26][2] ), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5426), .S(n52345));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[13][5] ), .I1(n23313), 
            .I2(GND_net), .I3(GND_net), .O(n52725));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_11  (.CI(n46114), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n46115));
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5427), .S(n52346));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_10_lut  (.I0(n59293), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n46113), .O(n25409)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5428), .S(n52342));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5429), .S(n52339));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5430), .S(n52337));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5431), .S(n52347));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5432), .S(n52348));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5433), .S(n52349));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[10][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5434));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27][2] ), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5435), .S(n52350));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1180 (.I0(n23199), .I1(n23375), .I2(Kp_23__N_645), 
            .I3(n52455), .O(n14_adj_5436));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n26797), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5437), .S(n52336));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5438), .S(n52340));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_10  (.CI(n46113), .I0(n25674), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n46114));
    SB_LUT4 i7_4_lut_adj_1181 (.I0(\data_in_frame[8][6] ), .I1(n14_adj_5436), 
            .I2(n10_adj_5434), .I3(n23135), .O(n52749));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_9_lut  (.I0(n59294), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n46112), .O(n25407)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i5_4_lut_adj_1182 (.I0(n52749), .I1(n52788), .I2(\data_in_frame[17] [3]), 
            .I3(n52725), .O(n12_adj_5439));
    defparam i5_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5440), .S(n52341));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_9  (.CI(n46112), .I0(n25674), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n46113));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_8_lut  (.I0(n59298), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n46111), .O(n25405)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i6_4_lut_adj_1183 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_5439), 
            .I2(n52972), .I3(n52692), .O(n54169));
    defparam i6_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1184 (.I0(\data_in_frame[17] [4]), .I1(n52749), 
            .I2(n54985), .I3(\data_in_frame[15] [3]), .O(n54113));
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1185 (.I0(n52656), .I1(\data_in_frame[12] [6]), 
            .I2(n23283), .I3(GND_net), .O(n53064));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n51701));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5441), .S(n52338));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1186 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n52785));
    defparam i2_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n26787), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13448_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n27154));
    defparam i13448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2978), .D(n3_adj_5442), .S(n52351));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n26786), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), 
            .C(clk16MHz), .E(n2978), .D(n1_adj_5443), .S(n52328));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2978), .D(n1_adj_5444), .S(n52329));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[3] [6]), .I1(n25709), .I2(n25766), 
            .I3(rx_data[6]), .O(n51695));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut.LUT_INIT = 16'h3a0a;
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(\byte_transmit_counter[3] ), 
            .C(clk16MHz), .E(n2978), .D(n1_adj_5445), .S(n52330));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5446), .S(n52207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5447), .S(n52208));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5448), .S(n52209));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(\byte_transmit_counter[4] ), 
            .C(clk16MHz), .E(n2978), .D(n1_adj_5449), .S(n52331));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5450), .S(n52210));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n2978), .D(n1_adj_5451), .S(n52332));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n2978), .D(n1_adj_5452), .S(n52333));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n2978), .D(n1_adj_5453), .S(n52334));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5454), .S(n52211));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5455), .S(n52212));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n26782), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n28044), .D(n2_adj_5456), .S(n26215));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5457), .S(n52213));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n28046), .D(n2_adj_5458), .S(n26213));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut_adj_1187 (.I0(\data_in_frame[3] [5]), .I1(n25709), 
            .I2(n25766), .I3(rx_data[5]), .O(n51691));
    defparam i12_4_lut_adj_1187.LUT_INIT = 16'h3a0a;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5459), .S(n52214));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5460), .S(n52215));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n28052), .D(n2_adj_5461), .S(n26207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3521[0]), .C(clk16MHz), 
            .E(n2978), .D(n1_adj_5462), .S(n26205));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2978), .D(n5_adj_5463), 
            .S(n26204));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5464), .S(n52216));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1188 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [5]), 
            .I2(n52834), .I3(n6_adj_5465), .O(n48509));
    defparam i4_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2978), .D(n24257), 
            .S(n26200));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1189 (.I0(n53064), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[14] [6]), .O(n14_adj_5466));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1190 (.I0(n53146), .I1(n14_adj_5466), .I2(n10_adj_5467), 
            .I3(n23375), .O(n52828));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1191 (.I0(\data_in_frame[19] [3]), .I1(n52828), 
            .I2(n48509), .I3(\data_in_frame[17] [1]), .O(n47491));
    defparam i2_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1192 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[19] [5]), 
            .I2(n54113), .I3(n54169), .O(n52816));
    defparam i3_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n2978), .D(n1_adj_5468), .S(n52327));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n26769), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13451_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n27157));
    defparam i13451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n26768), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_8  (.CI(n46111), .I0(n25674), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n46112));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_7_lut  (.I0(n59299), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n46110), .O(n25403)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_7  (.CI(n46110), .I0(n25674), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n46111));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47605 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n62511));
    defparam byte_transmit_counter_0__bdd_4_lut_47605.LUT_INIT = 16'he4aa;
    SB_LUT4 n62511_bdd_4_lut (.I0(n62511), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n62514));
    defparam n62511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47590 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n62505));
    defparam byte_transmit_counter_0__bdd_4_lut_47590.LUT_INIT = 16'he4aa;
    SB_LUT4 n62505_bdd_4_lut (.I0(n62505), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n62508));
    defparam n62505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_6_lut  (.I0(n59300), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n46109), .O(n25401)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_6  (.CI(n46109), .I0(n25674), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n46110));
    SB_DFFR \FRAME_MATCHER.i_1933__i1  (.Q(\FRAME_MATCHER.i[1] ), .C(clk16MHz), 
            .D(n25395), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i13454_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n27160));
    defparam i13454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5469), .S(n52300));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5470), .S(n52299));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5471), .S(n52298));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5472), .S(n52297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5473), .S(n52296));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5474), .S(n52295));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n28093), .D(n2_adj_5475), .S(n26402));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5476), .S(n52294));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n28095), .D(n2_adj_5477), .S(n26400));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n28096), .D(n2_adj_5478), .S(n26399));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5479), .S(n52293));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5480), .S(n52292));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5481), .S(n52291));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5482), .S(n52290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5483), .S(n52289));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5484), .S(n52288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5485), .S(n52287));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5486), .S(n26391));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n28105), .D(n2_adj_5487), .S(n26390));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5488), .S(n52286));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1933__i2  (.Q(\FRAME_MATCHER.i[2] ), .C(clk16MHz), 
            .D(n25397), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n25399), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n25401), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n25403), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n25405), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n25407), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n25409), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n25411), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n25413), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n25415), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n25417), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n25419), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n25421), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n25423), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n25425), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n25427), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n25429), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n25431), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n25433), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n25435), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n25437), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n25439), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n25441), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n25443), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n25445), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n25447), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n25449), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n25451), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n25453), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1933__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n25455), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n26840));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n26843));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n27428));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n27427));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n27426));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n27425));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n27424));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n27423));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n27422));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n27421));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n27420));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n27419));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n27418));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n27417));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n27416));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n27415));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n27414));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n27413));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n27412));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n27411));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n27410));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n27409));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n27408));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n27407));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n27406));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n27405));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n27404));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n27403));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n27402));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n27401));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n27400));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n27399));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n27398));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n26846));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n26849));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n26852));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n26855));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10][0] ), .C(clk16MHz), 
           .D(n26858));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10][1] ), .C(clk16MHz), 
           .D(n26861));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10][2] ), .C(clk16MHz), 
           .D(n26864));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10][3] ), .C(clk16MHz), 
           .D(n26867));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10][4] ), .C(clk16MHz), 
           .D(n51689));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10]_c [5]), .C(clk16MHz), 
           .D(n51685));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n26876));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10][7] ), .C(clk16MHz), 
           .D(n26879));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n51563));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n51585));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n51561));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n51559));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n51557));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n51555));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n51553));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n51551));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n26906));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n26909));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n26912));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1193 (.I0(\data_in_frame[13][7] ), .I1(n47517), 
            .I2(\data_in_frame[17] [7]), .I3(n48465), .O(n10_adj_5489));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1194 (.I0(\data_in_frame[15] [5]), .I1(n10_adj_5489), 
            .I2(n52678), .I3(GND_net), .O(n22497));
    defparam i5_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1195 (.I0(n48650), .I1(\data_in_frame[20] [3]), 
            .I2(n52659), .I3(\data_in_frame[20] [4]), .O(n52845));
    defparam i3_4_lut_adj_1195.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5490));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5491), .S(n52285));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1197 (.I0(n23367), .I1(n47444), .I2(\data_in_frame[12] [4]), 
            .I3(n6_adj_5490), .O(n53170));
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_5_lut  (.I0(n59301), .I1(n25674), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n46108), .O(n25399)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(n54381), .I1(n53170), .I2(\data_in_frame[16] [7]), 
            .I3(GND_net), .O(n52752));
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h6969;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_5  (.CI(n46108), .I0(n25674), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n46109));
    SB_LUT4 i13458_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n27164));
    defparam i13458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_4_lut  (.I0(n59302), .I1(n25674), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n46107), .O(n25397)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_4  (.CI(n46107), .I0(n25674), .I1(\FRAME_MATCHER.i[2] ), 
            .CO(n46108));
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_3_lut  (.I0(n59303), .I1(n25674), 
            .I2(\FRAME_MATCHER.i[1] ), .I3(n46106), .O(n25395)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5492), .S(n52284));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5493), .S(n52283));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n51777));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5494), .S(n52282));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_3  (.CI(n46106), .I0(n25674), .I1(\FRAME_MATCHER.i[1] ), 
            .CO(n46107));
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n28111), .D(n2_adj_5495), .S(n26384));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1933_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1933_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(n52819), .I1(\data_in_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5496));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1200 (.I0(n52752), .I1(n54734), .I2(\data_in_frame[18][7] ), 
            .I3(n4_adj_5496), .O(n55049));
    defparam i2_4_lut_adj_1200.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23135));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(n22568), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n52875));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1933_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n46106));
    SB_LUT4 i1_2_lut_adj_1203 (.I0(Kp_23__N_950), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52455));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1204 (.I0(\data_in_frame[10]_c [5]), .I1(n4), .I2(\data_in_frame[12] [4]), 
            .I3(GND_net), .O(n52656));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(n23824), .I1(n53055), .I2(GND_net), 
            .I3(GND_net), .O(n47444));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_12__7__I_0_4035_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_645));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_12__7__I_0_4035_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n26937));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[13][6] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1247));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n26940));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2978), .D(n2_adj_5497), .S(n52281));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13461_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n27167));
    defparam i13461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1206 (.I0(n23375), .I1(n23824), .I2(\data_in_frame[12] [5]), 
            .I3(GND_net), .O(n23367));
    defparam i2_3_lut_adj_1206.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1207 (.I0(\data_in_frame[13][5] ), .I1(n52972), 
            .I2(n52577), .I3(n52510), .O(n24073));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_in_frame[13] [0]), .I1(n23367), 
            .I2(GND_net), .I3(GND_net), .O(n23821));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i13465_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n27171));
    defparam i13465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13483_3_lut_4_lut (.I0(n25685), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n27189));
    defparam i13483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n52577));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1210 (.I0(rx_data[6]), .I1(n10), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5499));
    defparam i2_2_lut_adj_1210.LUT_INIT = 16'h2222;
    SB_LUT4 i14_4_lut_adj_1211 (.I0(\data_in_frame[2]_c [6]), .I1(n38306), 
            .I2(n25768), .I3(n6_adj_5499), .O(n51693));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1211.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[13]_c [3]), .I1(n47517), 
            .I2(GND_net), .I3(GND_net), .O(n52969));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1213 (.I0(\data_in_frame[13][7] ), .I1(n52969), 
            .I2(n52577), .I3(n23294), .O(n47558));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1214 (.I0(n47452), .I1(n23107), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n14_adj_5500));
    defparam i5_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1215 (.I0(n53061), .I1(\data_in_frame[14] [1]), 
            .I2(\data_in_frame[13][7] ), .I3(n52831), .O(n15_adj_5501));
    defparam i6_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1216 (.I0(n15_adj_5501), .I1(n48450), .I2(n14_adj_5500), 
            .I3(\data_in_frame[9] [2]), .O(n23518));
    defparam i8_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52868));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1218 (.I0(\data_in_frame[11] [5]), .I1(n23627), 
            .I2(n47579), .I3(n6_adj_5502), .O(n48465));
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1219 (.I0(n48465), .I1(n52868), .I2(n23518), 
            .I3(n47558), .O(n54710));
    defparam i3_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1220 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[4] [5]), 
            .I2(n52889), .I3(n52738), .O(n53061));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n48127), .I1(n53061), .I2(GND_net), 
            .I3(GND_net), .O(n48370));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1222 (.I0(n47487), .I1(n24165), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n52848));
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1223 (.I0(n23234), .I1(n52848), .I2(\data_in_frame[12] [3]), 
            .I3(\data_in_frame[10][1] ), .O(n52834));
    defparam i3_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1224 (.I0(n52653), .I1(n52982), .I2(\data_in_frame[10][3] ), 
            .I3(n52469), .O(n12_adj_5503));   // verilog/coms.v(79[16:43])
    defparam i5_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1225 (.I0(\data_in_frame[5] [6]), .I1(n12_adj_5503), 
            .I2(n53131), .I3(\data_in_frame[6][1] ), .O(n23824));   // verilog/coms.v(79[16:43])
    defparam i6_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1226 (.I0(\data_in_frame[14] [5]), .I1(n23824), 
            .I2(n52834), .I3(\data_in_frame[12] [4]), .O(n54734));
    defparam i3_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(n48439), .I1(n48370), .I2(n23338), 
            .I3(\data_in_frame[10][2] ), .O(n53055));
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_in_frame[12] [2]), .I1(n53055), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5504));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1229 (.I0(\data_in_frame[14] [4]), .I1(n47989), 
            .I2(\data_in_frame[12] [3]), .I3(n6_adj_5504), .O(n54381));
    defparam i4_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_in_frame[16] [6]), .I1(n54734), 
            .I2(GND_net), .I3(GND_net), .O(n52857));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1231 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n47475), .I3(GND_net), .O(n47579));
    defparam i2_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53131));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1233 (.I0(n53152), .I1(n48127), .I2(n52662), 
            .I3(n53131), .O(n15_adj_5505));
    defparam i6_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i13983_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n27689));
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1234 (.I0(n15_adj_5505), .I1(n52906), .I2(n14_adj_5507), 
            .I3(\data_in_frame[8] [0]), .O(n47452));
    defparam i8_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1235 (.I0(n52541), .I1(n52900), .I2(n52985), 
            .I3(n52997), .O(n22_adj_5508));
    defparam i9_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1236 (.I0(n53155), .I1(n22_adj_5508), .I2(n16), 
            .I3(\data_in_frame[12] [0]), .O(n24));
    defparam i11_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i13986_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n27692));
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1237 (.I0(n23283), .I1(n24), .I2(n20_adj_5510), 
            .I3(n23149), .O(n48503));
    defparam i12_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[10][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n53140));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1239 (.I0(n53140), .I1(n23234), .I2(n52629), 
            .I3(n47797), .O(n14_adj_5511));
    defparam i6_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1240 (.I0(n23607), .I1(n52997), .I2(n24165), 
            .I3(\data_in_frame[11] [7]), .O(n13_adj_5512));
    defparam i5_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1241 (.I0(n13_adj_5512), .I1(\data_in_frame[14] [3]), 
            .I2(n14_adj_5511), .I3(GND_net), .O(n6_adj_5513));
    defparam i2_3_lut_adj_1241.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_in_frame[18]_c [6]), .I1(n55049), 
            .I2(GND_net), .I3(GND_net), .O(n52438));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1243 (.I0(\data_in_frame[18][7] ), .I1(n52886), 
            .I2(n52438), .I3(n23500), .O(n48578));
    defparam i3_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[18] [3]), .I1(n54710), 
            .I2(GND_net), .I3(GND_net), .O(n48650));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_4_lut (.I0(n2059), .I1(n2056), .I2(n2062), .I3(\FRAME_MATCHER.i_31__N_2483 ), 
            .O(n54168));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52671));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_in_frame[13]_c [3]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52510));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(n52702), .I1(n24017), .I2(n31_adj_5514), 
            .I3(n52909), .O(n10_adj_5515));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1248 (.I0(n21154), .I1(n52916), .I2(\data_in_frame[4] [3]), 
            .I3(\data_in_frame[4] [1]), .O(n28));   // verilog/coms.v(76[16:42])
    defparam i10_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(\data_in_frame[4] [7]), .I1(n28), .I2(n23091), 
            .I3(GND_net), .O(n32_adj_5516));   // verilog/coms.v(76[16:42])
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1249 (.I0(\data_in_frame[3][7] ), .I1(n52903), 
            .I2(n53000), .I3(n52526), .O(n30));   // verilog/coms.v(76[16:42])
    defparam i12_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1250 (.I0(Kp_23__N_724), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[3] [6]), .I3(n23670), .O(n31_adj_5517));   // verilog/coms.v(76[16:42])
    defparam i13_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i13989_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n27695));
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1251 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[5] [2]), 
            .I2(n52623), .I3(\data_in_frame[4] [2]), .O(n29_adj_5518));   // verilog/coms.v(76[16:42])
    defparam i11_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i13992_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n27698));
    defparam i13992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut (.I0(n29_adj_5518), .I1(n31_adj_5517), .I2(n30), 
            .I3(n32_adj_5516), .O(n48127));   // verilog/coms.v(76[16:42])
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[4] [5]), .I1(n48127), 
            .I2(GND_net), .I3(GND_net), .O(n52443));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_in_frame[5] [5]), .I1(n21154), 
            .I2(GND_net), .I3(GND_net), .O(n52738));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i13995_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n27701));
    defparam i13995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13998_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n27704));
    defparam i13998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[6][3] ), .I1(\data_in_frame[6][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5514));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1255 (.I0(\data_in_frame[6][1] ), .I1(\data_in_frame[6][2] ), 
            .I2(n31_adj_5514), .I3(\data_in_frame[6] [0]), .O(n52541));
    defparam i3_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i14001_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n27707));
    defparam i14001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14004_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52430), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n27710));
    defparam i14004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[5] [6]), .I1(n52889), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5519));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1257 (.I0(n23750), .I1(n23251), .I2(n52443), 
            .I3(n6_adj_5519), .O(n54753));
    defparam i4_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[8] [1]), .I1(n54753), 
            .I2(GND_net), .I3(GND_net), .O(n52878));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h9999;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(n52463), .I2(n52611), 
            .I3(\data_in_frame[1] [7]), .O(n20));   // verilog/coms.v(169[9:87])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h0990;
    SB_LUT4 i3_4_lut_adj_1259 (.I0(\data_in_frame[8] [0]), .I1(n52469), 
            .I2(\data_in_frame[3] [5]), .I3(n23763), .O(n23234));
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1260 (.I0(n23680), .I1(n52839), .I2(\data_in_frame[5] [1]), 
            .I3(n23149), .O(n10_adj_5520));
    defparam i4_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1261 (.I0(\data_in_frame[5] [0]), .I1(n52903), 
            .I2(\data_in_frame[7] [2]), .I3(GND_net), .O(n23797));
    defparam i2_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[2] [0]), .I1(n23706), 
            .I2(GND_net), .I3(GND_net), .O(n24017));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1263 (.I0(\data_in_frame[6] [5]), .I1(n53000), 
            .I2(n52662), .I3(\data_in_frame[6][4] ), .O(Kp_23__N_950));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n23607));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n23052));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(n23639), .I1(n23797), .I2(GND_net), 
            .I3(GND_net), .O(n24061));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1267 (.I0(n47487), .I1(n53017), .I2(n24061), 
            .I3(n23283), .O(n10_adj_5521));
    defparam i4_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i419_2_lut_3_lut (.I0(n2059), .I1(n2056), .I2(n3303), .I3(GND_net), 
            .O(n2110));   // verilog/coms.v(142[4] 144[7])
    defparam i419_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2487 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3521[0]), .I3(n38421), .O(n22848));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52702));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[2] [5]), .I1(n52463), 
            .I2(n24145), .I3(\data_in_frame[4] [7]), .O(n23993));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1270 (.I0(n23676), .I1(\data_in_frame[4] [4]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n53020));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1271 (.I0(\data_in_frame[6][6] ), .I1(\data_in_frame[1] [7]), 
            .I2(n53020), .I3(n52702), .O(n53155));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(\data_in_frame[4] [4]), .I1(n23149), 
            .I2(n23706), .I3(GND_net), .O(n23673));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n23673), .I1(n53155), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(n52595));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1274 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n22929), .I3(\FRAME_MATCHER.i[1] ), .O(n5_adj_5522));   // verilog/coms.v(158[12:15])
    defparam i1_3_lut_4_lut_adj_1274.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_in_frame[5] [1]), .I1(n52916), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5523));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(\data_in_frame[7] [3]), .I1(n23993), 
            .I2(n52492), .I3(n6_adj_5523), .O(n47475));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_in_frame[4] [5]), .I1(n52595), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_969));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1278 (.I0(\data_in_frame[0] [6]), .I1(n23220), 
            .I2(\data_in_frame[3][0] ), .I3(GND_net), .O(n23680));
    defparam i2_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1279 (.I0(\data_in_frame[5] [4]), .I1(n52871), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n23091));
    defparam i2_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5524));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 i13959_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n27665));
    defparam i13959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(n23_adj_5524), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[1] [6]), .O(n52506));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n23238));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[2][7] ), .I1(n23220), 
            .I2(GND_net), .I3(GND_net), .O(n52839));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1284 (.I0(n23091), .I1(\data_in_frame[7] [6]), 
            .I2(n23251), .I3(GND_net), .O(n23338));
    defparam i2_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_LUT4 i13962_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n27668));
    defparam i13962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1285 (.I0(n52492), .I1(n24145), .I2(\data_in_frame[5] [3]), 
            .I3(n52871), .O(n10_adj_5525));
    defparam i4_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1286 (.I0(n23680), .I1(n10_adj_5525), .I2(\data_in_frame[7] [4]), 
            .I3(GND_net), .O(n23318));
    defparam i5_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(n23318), .I1(n23338), .I2(GND_net), 
            .I3(GND_net), .O(n23812));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i13965_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n27671));
    defparam i13965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 data_in_frame_8__7__I_0_4031_2_lut (.I0(\data_in_frame[8][7] ), 
            .I1(\data_in_frame[8][6] ), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_675));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_8__7__I_0_4031_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52526));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_4_lut_adj_1289 (.I0(n25675), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n51803));
    defparam i11_4_lut_4_lut_adj_1289.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_2_lut (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n23763));   // verilog/coms.v(99[12:25])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n52653));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52623));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i13974_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n27680));
    defparam i13974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1292 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[3][7] ), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n52982));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1293 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[6][1] ), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n52592));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1294 (.I0(n52592), .I1(n52982), .I2(n23750), 
            .I3(GND_net), .O(n23269));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1295 (.I0(\data_in_frame[1] [5]), .I1(n23251), 
            .I2(\data_in_frame[1] [4]), .I3(n6_adj_5526), .O(n24165));
    defparam i4_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1296 (.I0(\data_in_frame[8] [2]), .I1(n24165), 
            .I2(n23269), .I3(GND_net), .O(n3));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1297 (.I0(n23269), .I1(n52906), .I2(n52466), 
            .I3(\data_in_frame[1] [6]), .O(n4));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1298 (.I0(n4), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1037));   // verilog/coms.v(77[16:43])
    defparam i2_2_lut_adj_1298.LUT_INIT = 16'h6666;
    SB_LUT4 i13977_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n27683));
    defparam i13977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(n48439), .I1(n53089), .I2(n48450), 
            .I3(Kp_23__N_1037), .O(n53017));
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2484 ), 
            .I2(n22848), .I3(\FRAME_MATCHER.i_31__N_2483 ), .O(n56449));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i3_4_lut_adj_1300 (.I0(n23670), .I1(n23993), .I2(\data_in_frame[7] [1]), 
            .I3(\data_in_frame[6][7] ), .O(n52635));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(PWMLimit[5]), .I1(n375), .I2(GND_net), .I3(GND_net), 
            .O(n11));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[4] [5]), .I1(n52635), 
            .I2(GND_net), .I3(GND_net), .O(n23627));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1302 (.I0(n23534), .I1(\data_in_frame[3][1] ), 
            .I2(\data_in_frame[7] [5]), .I3(\data_in_frame[3][3] ), .O(n12_adj_5528));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1303 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_5528), 
            .I2(n52506), .I3(\data_in_frame[5] [3]), .O(n47487));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1304 (.I0(n23283), .I1(\data_in_frame[11] [1]), 
            .I2(n23199), .I3(GND_net), .O(n53137));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 i8_2_lut (.I0(deadband[5]), .I1(n375), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_8));
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1305 (.I0(n53137), .I1(n47487), .I2(n52985), 
            .I3(n23627), .O(n14_adj_5530));
    defparam i6_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i434_4_lut_4_lut (.I0(n2056), .I1(n2062), .I2(n4452), .I3(n2059), 
            .O(n2125));   // verilog/coms.v(139[4] 141[7])
    defparam i434_4_lut_4_lut.LUT_INIT = 16'h0d05;
    SB_LUT4 i7_4_lut_adj_1306 (.I0(n7_adj_5531), .I1(n14_adj_5530), .I2(n10_adj_5532), 
            .I3(Kp_23__N_950), .O(n54985));
    defparam i7_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_in_frame[13]_c [3]), .I1(\data_in_frame[13][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n52692));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_in_frame[8][7] ), .I1(n52635), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5533));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1309 (.I0(\data_in_frame[11] [3]), .I1(n23607), 
            .I2(n52595), .I3(n6_adj_5533), .O(n23294));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_in_frame[3][7] ), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52909));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n53116));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2484 ), 
            .I2(\FRAME_MATCHER.i_31__N_2483 ), .I3(GND_net), .O(n5_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 i3_4_lut_adj_1312 (.I0(\data_in_frame[1] [4]), .I1(n53116), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[2] [0]), .O(n52466));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1313 (.I0(\data_in_frame[10][7] ), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[11] [2]), .O(n52925));
    defparam i3_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1314 (.I0(n13), .I1(n52900), .I2(n23676), .I3(n23673), 
            .O(n23639));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i13980_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n27686));
    defparam i13980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1315 (.I0(\data_in_frame[15] [5]), .I1(n23294), 
            .I2(n52692), .I3(n54985), .O(n52801));
    defparam i1_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1316 (.I0(n23639), .I1(n52925), .I2(n23283), 
            .I3(\data_in_frame[11] [0]), .O(n12_adj_5536));
    defparam i5_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1317 (.I0(\data_in_frame[9] [1]), .I1(n12_adj_5536), 
            .I2(\data_in_frame[15] [4]), .I3(n52510), .O(n54639));
    defparam i6_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(n54639), .I1(n52801), .I2(GND_net), 
            .I3(GND_net), .O(n23115));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h9999;
    SB_LUT4 i13971_3_lut_4_lut (.I0(n25675), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n27677));
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i45169_2_lut (.I0(n62616), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59358));
    defparam i45169_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46149_3_lut (.I0(n62550), .I1(n62478), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n61049));
    defparam i46149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41746_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56646));
    defparam i41746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41747_4_lut (.I0(n56646), .I1(n25461), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][0] ), .O(n56647));
    defparam i41747_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i41745_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56645));
    defparam i41745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41943_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56843));
    defparam i41943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1319 (.I0(\data_in_frame[20] [5]), .I1(n52671), 
            .I2(n48650), .I3(n48578), .O(n12_adj_5537));
    defparam i5_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i41944_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56844));
    defparam i41944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1320 (.I0(n48458), .I1(\data_in_frame[22] [1]), 
            .I2(\data_in_frame[21] [7]), .I3(n52755), .O(n10_adj_5538));
    defparam i4_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\data_in_frame[22] [5]), .I1(n52845), 
            .I2(GND_net), .I3(GND_net), .O(n52846));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i41683_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56583));
    defparam i41683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41682_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56582));
    defparam i41682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1322 (.I0(\data_in_frame[21] [6]), .I1(n52816), 
            .I2(n47491), .I3(\data_in_frame[23] [7]), .O(n54791));
    defparam i3_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1323 (.I0(\data_in_frame[19] [7]), .I1(n52846), 
            .I2(n10_adj_5538), .I3(\data_in_frame[19] [5]), .O(n7_adj_5539));
    defparam i1_4_lut_adj_1323.LUT_INIT = 16'h2112;
    SB_LUT4 i11755_2_lut (.I0(\byte_transmit_counter[1] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n25461));   // verilog/coms.v(109[34:55])
    defparam i11755_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i41394_4_lut (.I0(n1_adj_5290), .I1(n52695), .I2(n52942), 
            .I3(\data_in_frame[23] [1]), .O(n56282));
    defparam i41394_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i41740_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56640));
    defparam i41740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41741_4_lut (.I0(n56640), .I1(n25461), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][5] ), .O(n56641));
    defparam i41741_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i3_4_lut_adj_1324 (.I0(\data_in_frame[23] [5]), .I1(n52770), 
            .I2(Kp_23__N_1595), .I3(\data_in_frame[21] [3]), .O(n54763));
    defparam i3_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47689 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56594), .I2(n56595), .I3(\byte_transmit_counter[2] ), 
            .O(n62499));
    defparam byte_transmit_counter_1__bdd_4_lut_47689.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1325 (.I0(\data_in_frame[23] [3]), .I1(n52942), 
            .I2(\data_in_frame[21] [2]), .I3(\data_in_frame[21] [1]), .O(n54087));
    defparam i3_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i41739_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56639));
    defparam i41739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1326 (.I0(\data_in_frame[22] [7]), .I1(n12_adj_5537), 
            .I2(n53014), .I3(n47264), .O(n54247));
    defparam i6_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i41477_4_lut (.I0(n48578), .I1(n54763), .I2(n53014), .I3(\data_in_frame[23] [0]), 
            .O(n56367));
    defparam i41477_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i45299_2_lut (.I0(n62580), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59368));
    defparam i45299_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_1327 (.I0(n56282), .I1(n7_adj_5539), .I2(n9_adj_5291), 
            .I3(n54791), .O(n55172));
    defparam i5_4_lut_adj_1327.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1328 (.I0(n47491), .I1(n48593), .I2(n52770), 
            .I3(\data_in_frame[23] [6]), .O(n4_adj_5540));
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'h9669;
    SB_LUT4 i46275_3_lut (.I0(n62700), .I1(n62436), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n61175));
    defparam i46275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41703_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56603));
    defparam i41703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41704_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56604));
    defparam i41704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1329 (.I0(\data_in_frame[23] [4]), .I1(n52617), 
            .I2(Kp_23__N_1595), .I3(n48578), .O(n54019));
    defparam i3_4_lut_adj_1329.LUT_INIT = 16'h9669;
    SB_LUT4 i41923_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56823));
    defparam i41923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41922_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56822));
    defparam i41922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1330 (.I0(n55172), .I1(n56367), .I2(n54247), 
            .I3(n54087), .O(n12_adj_5541));
    defparam i2_4_lut_adj_1330.LUT_INIT = 16'h0020;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[18] [2]), 
            .I2(n52791), .I3(GND_net), .O(n8_adj_5542));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1331 (.I0(\data_in_frame[22] [0]), .I1(n48593), 
            .I2(\data_in_frame[19] [6]), .I3(n6_adj_5543), .O(n54630));
    defparam i4_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1332 (.I0(\data_in_frame[20] [1]), .I1(n52659), 
            .I2(n52791), .I3(\data_in_frame[22] [3]), .O(n10_adj_5544));
    defparam i4_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(\data_in_frame[22] [2]), .I1(n53134), 
            .I2(n52988), .I3(n52755), .O(n54968));
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i41802_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56702));
    defparam i41802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1334 (.I0(\data_in_frame[22] [6]), .I1(n52735), 
            .I2(\data_in_frame[20] [4]), .I3(GND_net), .O(n54614));
    defparam i2_3_lut_adj_1334.LUT_INIT = 16'h9696;
    SB_LUT4 i41803_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56703));
    defparam i41803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1335 (.I0(\data_in_frame[21] [5]), .I1(n12_adj_5541), 
            .I2(n54019), .I3(n4_adj_5540), .O(n16_adj_5545));
    defparam i6_4_lut_adj_1335.LUT_INIT = 16'h4080;
    SB_LUT4 i41800_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56700));
    defparam i41800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41799_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56699));
    defparam i41799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41808_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56708));
    defparam i41808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41809_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56709));
    defparam i41809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1336 (.I0(n54630), .I1(n54272), .I2(n8_adj_5542), 
            .I3(\data_in_frame[22] [4]), .O(n14_adj_5546));
    defparam i4_4_lut_adj_1336.LUT_INIT = 16'h2882;
    SB_LUT4 i41770_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56670));
    defparam i41770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41769_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56669));
    defparam i41769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41449_4_lut (.I0(\data_in_frame[19] [7]), .I1(n54968), .I2(n10_adj_5544), 
            .I3(n52988), .O(n56339));
    defparam i41449_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i41811_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56711));
    defparam i41811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1337 (.I0(n54614), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [2]), .I3(n54729), .O(n13_adj_5547));
    defparam i3_4_lut_adj_1337.LUT_INIT = 16'h8228;
    SB_LUT4 i41812_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56712));
    defparam i41812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41752_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56652));
    defparam i41752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41751_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56651));
    defparam i41751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41826_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56726));
    defparam i41826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41827_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56727));
    defparam i41827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41695_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56595));
    defparam i41695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1338 (.I0(n13_adj_5547), .I1(n56339), .I2(n14_adj_5546), 
            .I3(n16_adj_5545), .O(n30905));
    defparam i9_4_lut_adj_1338.LUT_INIT = 16'h2000;
    SB_LUT4 i41694_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56594));
    defparam i41694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1339 (.I0(n53116), .I1(\data_in_frame[8] [1]), 
            .I2(n52443), .I3(n52948), .O(n15_adj_5548));
    defparam i6_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1340 (.I0(n15_adj_5548), .I1(n52592), .I2(n14_adj_5549), 
            .I3(n31_adj_5514), .O(n54671));
    defparam i8_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1341 (.I0(n7_adj_5531), .I1(n54753), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n10_adj_5550));
    defparam i2_3_lut_adj_1341.LUT_INIT = 16'h4141;
    SB_LUT4 i6_4_lut_adj_1342 (.I0(n48370), .I1(n23627), .I2(n23797), 
            .I3(n54671), .O(n14_adj_5551));
    defparam i6_4_lut_adj_1342.LUT_INIT = 16'h0002;
    SB_LUT4 i7_4_lut_adj_1343 (.I0(n3), .I1(n14_adj_5551), .I2(n10_adj_5550), 
            .I3(n47487), .O(n55189));
    defparam i7_4_lut_adj_1343.LUT_INIT = 16'h0040;
    SB_LUT4 i6_4_lut_adj_1344 (.I0(n23338), .I1(n23318), .I2(n4), .I3(n55189), 
            .O(n16_adj_5552));
    defparam i6_4_lut_adj_1344.LUT_INIT = 16'h0800;
    SB_LUT4 i41475_3_lut (.I0(n23283), .I1(Kp_23__N_950), .I2(\data_in_frame[8][6] ), 
            .I3(GND_net), .O(n56365));
    defparam i41475_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i8_3_lut (.I0(n23639), .I1(n16_adj_5552), .I2(n23199), .I3(GND_net), 
            .O(n18_adj_5553));
    defparam i8_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i9_4_lut_adj_1345 (.I0(n25), .I1(n18_adj_5553), .I2(n56365), 
            .I3(n47475), .O(LED_N_3384));
    defparam i9_4_lut_adj_1345.LUT_INIT = 16'h0400;
    SB_LUT4 i13125_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[7]), 
            .I3(\data_in_frame[8][7] ), .O(n26831));
    defparam i13125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(Kp_23__N_1724), .I1(n30905), .I2(GND_net), 
            .I3(GND_net), .O(n25012));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h8888;
    SB_LUT4 i17211_4_lut (.I0(\FRAME_MATCHER.i_31__N_2489 ), .I1(Kp_23__N_1724), 
            .I2(LED_N_3384), .I3(n30905), .O(n25059));   // verilog/coms.v(18[27:29])
    defparam i17211_4_lut.LUT_INIT = 16'he420;
    SB_LUT4 i13122_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[6]), 
            .I3(\data_in_frame[8][6] ), .O(n26828));
    defparam i13122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13119_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[5]), 
            .I3(\data_in_frame[8][5] ), .O(n26825));
    defparam i13119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13116_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[4]), 
            .I3(\data_in_frame[8][4] ), .O(n26822));
    defparam i13116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13113_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[3]), 
            .I3(\data_in_frame[8]_c [3]), .O(n26819));
    defparam i13113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13110_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n26816));
    defparam i13110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13107_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n26813));
    defparam i13107_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1347 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [12]), .O(n10_adj_5555));
    defparam i4_4_lut_adj_1347.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [29]), .O(n34_adj_5556));
    defparam i13_4_lut_adj_1348.LUT_INIT = 16'hfffe;
    SB_LUT4 i13104_3_lut_4_lut (.I0(n8_adj_5554), .I1(n52424), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n26810));
    defparam i13104_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1349 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(n10_adj_5555), .I3(\FRAME_MATCHER.i [27]), .O(n23_adj_5557));
    defparam i2_4_lut_adj_1349.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1350 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5558));
    defparam i1_2_lut_adj_1350.LUT_INIT = 16'heeee;
    SB_LUT4 i13149_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n26855));
    defparam i13149_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut_adj_1351 (.I0(n23_adj_5557), .I1(n34_adj_5556), .I2(\FRAME_MATCHER.i [22]), 
            .I3(\FRAME_MATCHER.i [26]), .O(n38));
    defparam i17_4_lut_adj_1351.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1352 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(\FRAME_MATCHER.i [6]), .I3(\FRAME_MATCHER.i [5]), .O(n36));
    defparam i15_4_lut_adj_1352.LUT_INIT = 16'hfffe;
    SB_LUT4 i13146_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n26852));
    defparam i13146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13143_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n26849));
    defparam i13143_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n22_adj_5558), .O(n37_adj_5559));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1353 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [21]), .O(n35));
    defparam i14_4_lut_adj_1353.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37_adj_5559), .I2(n36), .I3(n38), 
            .O(n22929));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24457_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22929), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i24457_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i471_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2490 ), .I2(GND_net), 
            .I3(GND_net), .O(n2173));   // verilog/coms.v(148[4] 304[11])
    defparam i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13140_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n26846));
    defparam i13140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13137_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n26843));
    defparam i13137_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13134_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n26840));
    defparam i13134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13131_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n26837));
    defparam i13131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13128_3_lut_4_lut (.I0(n35699), .I1(n52424), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n26834));
    defparam i13128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_4_lut (.I0(n2056), .I1(n4452), .I2(n56449), .I3(\FRAME_MATCHER.i_31__N_2490 ), 
            .O(n54637));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i431_2_lut_3_lut (.I0(n2056), .I1(n4452), .I2(n2059), .I3(GND_net), 
            .O(n2122));   // verilog/coms.v(145[4] 147[7])
    defparam i431_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i44565_2_lut (.I0(\data_out_frame[0][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n59215));
    defparam i44565_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44809_2_lut (.I0(\data_out_frame[3][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n59216));
    defparam i44809_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2]_c [6]), 
            .I2(n52458), .I3(n10_adj_5520), .O(n52903));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(n10), .I1(n38302), .I2(GND_net), .I3(GND_net), 
            .O(n52412));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'hbbbb;
    SB_LUT4 i17_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n13_c));   // verilog/coms.v(105[12:33])
    defparam i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n4_adj_5287));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2]_c [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n24145));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i12033_3_lut_4_lut (.I0(n10_adj_9), .I1(n38302), .I2(reset), 
            .I3(n8_adj_5554), .O(n25739));
    defparam i12033_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[6][4] ), .O(n51791));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1356 (.I0(n25721), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n51797));
    defparam i1_4_lut_4_lut_4_lut_adj_1356.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n10_adj_9), .I1(n38302), .I2(n35706), 
            .I3(\FRAME_MATCHER.i[0] ), .O(n25675));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[25] [7]), .I3(GND_net), .O(n8_adj_5561));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1358 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[9] [2]), .O(n23958));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5554));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n35699));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'hefef;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[12] [3]), .I1(n1513), .I2(\data_out_frame[17] [0]), 
            .I3(n4_adj_5562), .O(n24203));   // verilog/coms.v(77[16:43])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n52564), .I3(GND_net), .O(n1655));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(n53052), .I3(GND_net), .O(n52862));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n4_adj_5562));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1364 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[10] [4]), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5286));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1364.LUT_INIT = 16'ha088;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n23958), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[10][7] ), .O(n10_adj_5532));   // verilog/coms.v(88[17:63])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n52894));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(\FRAME_MATCHER.i[2] ), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(GND_net), .O(n35696));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[8] [4]), .O(n23577));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n52913));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1369 (.I0(\data_out_frame[6] [2]), .I1(n52484), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[5] [7]), .O(n52475));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1370 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[9] [6]), .O(n52567));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n53098));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1372 (.I0(n25705), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n51825));
    defparam i1_4_lut_4_lut_4_lut_adj_1372.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5494));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1373 (.I0(n25705), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n51823));
    defparam i1_4_lut_4_lut_4_lut_adj_1373.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1374 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[6] [0]), .O(n53083));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44849_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59303));   // verilog/coms.v(158[12:15])
    defparam i44849_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44848_2_lut (.I0(\FRAME_MATCHER.i[2] ), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59302));   // verilog/coms.v(158[12:15])
    defparam i44848_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44847_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59301));   // verilog/coms.v(158[12:15])
    defparam i44847_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1375 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [2]), .I3(\data_out_frame[16] [3]), 
            .O(n52587));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1376 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[13] [3]), 
            .I2(n10_adj_5563), .I3(n52842), .O(n52604));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n23964));
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n53043));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [3]), .I3(GND_net), .O(n53175));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(\data_out_frame[15] [6]), .I1(n47380), 
            .I2(n24120), .I3(GND_net), .O(n47422));
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut (.I0(n54100), .I1(n52862), .I2(\data_out_frame[19] [0]), 
            .I3(GND_net), .O(n10_adj_5564));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i6_3_lut_4_lut_adj_1381 (.I0(\data_out_frame[12] [0]), .I1(n52851), 
            .I2(\data_out_frame[6] [1]), .I3(\data_out_frame[10] [3]), .O(n17_adj_5565));
    defparam i6_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1382 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(n23427), .I3(n23005), .O(n1312));
    defparam i2_3_lut_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n52951));
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n6_adj_5566));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1385 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[11] [5]), 
            .I2(n52851), .I3(n53035), .O(n23601));
    defparam i1_2_lut_4_lut_adj_1385.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1386 (.I0(n53024), .I1(\data_out_frame[16] [1]), 
            .I2(n47581), .I3(n23155), .O(n48240));
    defparam i2_3_lut_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[16] [3]), .I1(n54100), 
            .I2(n52705), .I3(GND_net), .O(n53024));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1388 (.I0(n52520), .I1(n10_adj_5567), .I2(n52892), 
            .I3(\data_out_frame[23] [2]), .O(n4_adj_5568));
    defparam i1_2_lut_4_lut_adj_1388.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1389 (.I0(n25707), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[10][4] ), .O(n51689));
    defparam i1_4_lut_4_lut_4_lut_adj_1389.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1390 (.I0(n25707), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[10]_c [5]), .O(n51685));
    defparam i1_4_lut_4_lut_4_lut_adj_1390.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1391 (.I0(\data_out_frame[20] [0]), .I1(n21050), 
            .I2(n10_adj_5569), .I3(n23568), .O(n52776));
    defparam i5_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1392 (.I0(\data_out_frame[20] [3]), .I1(n48527), 
            .I2(\data_out_frame[20] [2]), .I3(n2054), .O(n48568));
    defparam i1_2_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\data_out_frame[11] [5]), .I1(n52851), 
            .I2(n53035), .I3(GND_net), .O(n53036));
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1394 (.I0(\data_out_frame[22] [4]), .I1(n23185), 
            .I2(n52627), .I3(n52991), .O(n54349));
    defparam i2_3_lut_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1395 (.I0(\data_out_frame[11] [5]), .I1(n52851), 
            .I2(n24120), .I3(n52601), .O(n47527));
    defparam i2_3_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut (.I0(n47720), .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[19] [6]), 
            .I3(n52807), .O(n11_adj_5570));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1396 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n52598));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1396.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1397 (.I0(\data_out_frame[20] [3]), .I1(n48527), 
            .I2(\data_out_frame[22] [5]), .I3(n52860), .O(n23185));
    defparam i2_3_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1398 (.I0(n48527), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [1]), .I3(n54449), .O(n21097));
    defparam i2_3_lut_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1399 (.I0(\data_out_frame[20] [4]), .I1(n54473), 
            .I2(n48240), .I3(\data_out_frame[20] [5]), .O(n53046));
    defparam i2_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1400 (.I0(\data_out_frame[24] [3]), .I1(n52776), 
            .I2(n53046), .I3(n48247), .O(n52632));
    defparam i1_2_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(\data_out_frame[24] [5]), .I1(n48527), 
            .I2(n52478), .I3(n54449), .O(n52716));
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1402 (.I0(n23713), .I1(\data_out_frame[23] [3]), 
            .I2(n48629), .I3(n48474), .O(n52764));
    defparam i1_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1403 (.I0(\data_out_frame[23] [0]), .I1(n48523), 
            .I2(n10_adj_5571), .I3(n2394), .O(n52552));
    defparam i5_3_lut_4_lut_adj_1403.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [5]), .I3(n48523), .O(n10_adj_5572));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21411_3_lut_4_lut (.I0(\Kp[6] ), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n26797));
    defparam i21411_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1404 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(\data_out_frame[18] [1]), .I3(\data_out_frame[18] [0]), 
            .O(n6_adj_5573));
    defparam i1_2_lut_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [0]), 
            .O(n52343));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1405 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [1]), 
            .O(n52344));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1405.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1406 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26][2] ), 
            .O(n52345));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1406.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1407 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [3]), 
            .O(n52346));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1407.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1408 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [4]), 
            .O(n52342));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1408.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1409 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [5]), 
            .O(n52339));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1409.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1410 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [6]), 
            .O(n52337));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1410.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1411 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[26] [7]), 
            .O(n52347));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1411.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5488));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1412 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [0]), 
            .O(n52348));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1412.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1413 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[9] [1]), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1413.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1414 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [1]), 
            .O(n52349));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1414.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\data_out_frame[4] [7]), .I1(n1168), 
            .I2(n23531), .I3(GND_net), .O(n22594));
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5486));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1416 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27][2] ), 
            .O(n52350));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1416.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_70_i2_4_lut (.I0(\data_out_frame[8] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1417 (.I0(\data_out_frame[4] [7]), .I1(n1168), 
            .I2(n23869), .I3(n10_adj_5574), .O(n24120));
    defparam i5_3_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1418 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [3]), 
            .O(n52336));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1418.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1419 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [4]), 
            .O(n52340));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1419.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1420 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [5]), 
            .O(n52341));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1420.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5481));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1421 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [6]), 
            .O(n52338));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1421.LUT_INIT = 16'h5100;
    SB_LUT4 select_775_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5480));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1422 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(\data_out_frame[27] [7]), 
            .O(n52351));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1422.LUT_INIT = 16'h5100;
    SB_LUT4 i17_3_lut_4_lut (.I0(\data_out_frame[5] [0]), .I1(n1168), .I2(\data_out_frame[6] [7]), 
            .I3(\data_out_frame[4] [5]), .O(n23531));   // verilog/coms.v(88[17:70])
    defparam i17_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5478));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21634_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n27630));   // verilog/coms.v(130[12] 305[6])
    defparam i21634_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1423 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[4] [6]), .O(n23688));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i13318_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n27024));
    defparam i13318_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13305_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n27011));
    defparam i13305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13299_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n27005));
    defparam i13299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1424 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[7] [5]), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1424.LUT_INIT = 16'ha088;
    SB_LUT4 i13293_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n26999));
    defparam i13293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1425 (.I0(n24097), .I1(n52523), .I2(\data_out_frame[19] [3]), 
            .I3(n53040), .O(n48601));
    defparam i1_2_lut_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12499_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n26205));   // verilog/coms.v(130[12] 305[6])
    defparam i12499_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13290_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n26996));
    defparam i13290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12498_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2489 ), 
            .I2(n24628), .I3(n23_adj_5575), .O(n26204));   // verilog/coms.v(130[12] 305[6])
    defparam i12498_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 select_775_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_4_lut_adj_1426 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2487 ), 
            .I2(\FRAME_MATCHER.i_31__N_2490 ), .I3(n30909), .O(n6_adj_5576));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_LUT4 select_775_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13287_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n26993));
    defparam i13287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12494_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2484 ), 
            .I2(GND_net), .I3(GND_net), .O(n26200));   // verilog/coms.v(130[12] 305[6])
    defparam i12494_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_775_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11632_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n25336));   // verilog/coms.v(109[34:55])
    defparam i11632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13923_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [1]), 
            .I3(current_limit[1]), .O(n27629));   // verilog/coms.v(130[12] 305[6])
    defparam i13923_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13284_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n26990));
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i41731_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56631));
    defparam i41731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41732_4_lut (.I0(n56631), .I1(n25336), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n56632));
    defparam i41732_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i13281_3_lut_4_lut (.I0(n8_adj_5506), .I1(n52424), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n26987));
    defparam i13281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i41730_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56630));
    defparam i41730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44846_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59300));   // verilog/coms.v(158[12:15])
    defparam i44846_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24985146_i1_3_lut (.I0(n62652), .I1(n62412), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14));
    defparam i24985146_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n37));
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h8080;
    SB_LUT4 i44845_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59299));   // verilog/coms.v(158[12:15])
    defparam i44845_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5506));
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_4_lut_adj_1429 (.I0(\data_out_frame[6] [6]), .I1(n1130), 
            .I2(\data_out_frame[11] [1]), .I3(n52529), .O(n23041));
    defparam i2_3_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(\data_out_frame[6] [6]), .I1(n1130), 
            .I2(n23945), .I3(n23531), .O(n44537));
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n52489));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[4] [2]), .O(n32));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(\data_out_frame[6] [1]), .I1(n23012), 
            .I2(\data_out_frame[11] [0]), .I3(n52475), .O(n53161));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_4_lut (.I0(\data_out_frame[6] [1]), .I1(n23012), .I2(n52951), 
            .I3(\data_out_frame[8] [1]), .O(n23_adj_5578));   // verilog/coms.v(76[16:42])
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13922_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [2]), 
            .I3(current_limit[2]), .O(n27628));   // verilog/coms.v(130[12] 305[6])
    defparam i13922_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n52705), .I3(n4_adj_5562), .O(n52892));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n56647), .I3(n56645), 
            .O(n7_adj_5579));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n56641), .I3(n56639), 
            .O(n7_adj_5580));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13918_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [6]), 
            .I3(current_limit[6]), .O(n27624));   // verilog/coms.v(130[12] 305[6])
    defparam i13918_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n56632), .I3(n56630), 
            .O(n7_adj_5285));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n56674), .I3(n56672), 
            .O(n7));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13929_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n27635));   // verilog/coms.v(130[12] 305[6])
    defparam i13929_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1435 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(n6_adj_5576), .I3(\FRAME_MATCHER.i_31__N_2488 ), .O(n24257));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1435.LUT_INIT = 16'haaa8;
    SB_LUT4 i12_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), .I1(\byte_transmit_counter[1] ), 
            .I2(n56635), .I3(n56633), .O(n52053));   // verilog/coms.v(109[34:55])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_775_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(LED_c), .I1(LED_N_3384), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5575));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_3_lut_adj_1437 (.I0(\data_out_frame[16] [0]), .I1(n52604), 
            .I2(n62162), .I3(GND_net), .O(n7_adj_5581));
    defparam i2_2_lut_3_lut_adj_1437.LUT_INIT = 16'h6969;
    SB_LUT4 i17207_4_lut (.I0(Kp_23__N_1724), .I1(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2485 ), .I3(LED_c), .O(n30913));   // verilog/coms.v(118[11:12])
    defparam i17207_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i1_2_lut_adj_1438 (.I0(n30913), .I1(n25012), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5463));
    defparam i1_2_lut_adj_1438.LUT_INIT = 16'heeee;
    SB_LUT4 select_1625_Select_0_i1_2_lut (.I0(tx_transmit_N_3392), .I1(\FRAME_MATCHER.i_31__N_2487 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_1625_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_775_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(\data_out_frame[16] [0]), .I1(n52604), 
            .I2(n52674), .I3(GND_net), .O(n47944));
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5289));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1440 (.I0(n24097), .I1(n52523), .I2(n48452), 
            .I3(GND_net), .O(n52807));
    defparam i1_2_lut_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1441 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[4] [3]), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1441.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20442_3_lut (.I0(n25739), .I1(rx_data[5]), .I2(\data_in_frame[16]_c [5]), 
            .I3(GND_net), .O(n27142));   // verilog/coms.v(94[13:20])
    defparam i20442_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 select_775_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(n8_adj_5554), .I1(n10), .I2(n38302), 
            .I3(GND_net), .O(n25705));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'hefef;
    SB_LUT4 select_775_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_1044_i1_3_lut_4_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3][0] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i1_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i5_3_lut_4_lut_adj_1443 (.I0(n23149), .I1(n23676), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[3] [5]), .O(n14_adj_5549));
    defparam i5_3_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i19866_3_lut (.I0(n151), .I1(n203), .I2(n181), .I3(GND_net), 
            .O(n33540));
    defparam i19866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_775_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(n54639), .I1(n52801), .I2(\data_in_frame[17] [6]), 
            .I3(\data_in_frame[20] [0]), .O(n52755));
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h9669;
    SB_LUT4 i19867_3_lut (.I0(n33540), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[3] ));
    defparam i19867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13909_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [7]), 
            .I3(current_limit[15]), .O(n27615));   // verilog/coms.v(130[12] 305[6])
    defparam i13909_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n62499_bdd_4_lut (.I0(n62499), .I1(n56727), .I2(n56726), .I3(\byte_transmit_counter[2] ), 
            .O(n14_adj_5582));
    defparam n62499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(\data_in_frame[8][4] ), .I1(\data_in_frame[3][7] ), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[6][3] ), .O(n53152));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_223_i3_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n52764), .I3(\data_out_frame[25] [6]), 
            .O(n3_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i23744_3_lut (.I0(\current[11] ), .I1(\data[11] ), .I2(n25021), 
            .I3(GND_net), .O(n27452));
    defparam i23744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13913_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [3]), 
            .I3(current_limit[11]), .O(n27619));   // verilog/coms.v(130[12] 305[6])
    defparam i13913_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13915_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [1]), 
            .I3(current_limit[9]), .O(n27621));   // verilog/coms.v(130[12] 305[6])
    defparam i13915_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13692_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n27398));   // verilog/coms.v(130[12] 305[6])
    defparam i13692_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_222_i3_4_lut (.I0(n4_adj_5583), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5584), .I3(n4_adj_5568), .O(n3_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_222_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13709_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n27415));   // verilog/coms.v(130[12] 305[6])
    defparam i13709_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13715_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n27421));   // verilog/coms.v(130[12] 305[6])
    defparam i13715_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13714_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n27420));   // verilog/coms.v(130[12] 305[6])
    defparam i13714_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(n23234), .I1(\data_in_frame[8] [1]), 
            .I2(n54753), .I3(GND_net), .O(n48439));
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h6969;
    SB_LUT4 i13713_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n27419));   // verilog/coms.v(130[12] 305[6])
    defparam i13713_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1447 (.I0(\data_in_frame[8][7] ), .I1(\data_in_frame[8][6] ), 
            .I2(n23318), .I3(n23338), .O(n53089));
    defparam i1_2_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1448 (.I0(\data_in_frame[4] [5]), .I1(n52595), 
            .I2(n47475), .I3(GND_net), .O(n48450));
    defparam i1_2_lut_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i44842_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59298));   // verilog/coms.v(158[12:15])
    defparam i44842_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13712_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n27418));   // verilog/coms.v(130[12] 305[6])
    defparam i13712_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13711_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n27417));   // verilog/coms.v(130[12] 305[6])
    defparam i13711_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[5] [6]), .O(n6_adj_5526));
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i13239_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n26945));   // verilog/coms.v(130[12] 305[6])
    defparam i13239_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(GND_net), .O(n23750));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_221_i3_4_lut (.I0(n48611), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n48499), .I3(\data_out_frame[25] [4]), .O(n3_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i13722_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n27428));   // verilog/coms.v(130[12] 305[6])
    defparam i13722_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13910_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [6]), 
            .I3(current_limit[14]), .O(n27616));   // verilog/coms.v(130[12] 305[6])
    defparam i13910_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47580 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56651), .I2(n56652), .I3(\byte_transmit_counter[2] ), 
            .O(n62493));
    defparam byte_transmit_counter_1__bdd_4_lut_47580.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3][4] ), .I3(GND_net), .O(n23251));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(n52712), .I3(GND_net), .O(n47720));
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i13721_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n27427));   // verilog/coms.v(130[12] 305[6])
    defparam i13721_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13720_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n27426));   // verilog/coms.v(130[12] 305[6])
    defparam i13720_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13719_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n27425));   // verilog/coms.v(130[12] 305[6])
    defparam i13719_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1453 (.I0(\data_out_frame[16] [2]), .I1(n48587), 
            .I2(n53024), .I3(\data_out_frame[18] [4]), .O(n52520));
    defparam i1_3_lut_4_lut_adj_1453.LUT_INIT = 16'h9669;
    SB_LUT4 i13718_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n27424));   // verilog/coms.v(130[12] 305[6])
    defparam i13718_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1454 (.I0(\data_out_frame[16] [2]), .I1(n48587), 
            .I2(\data_out_frame[18] [3]), .I3(n53078), .O(n54473));
    defparam i2_3_lut_4_lut_adj_1454.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1455 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2][7] ), .I3(n23220), .O(n52492));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i44834_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59294));   // verilog/coms.v(158[12:15])
    defparam i44834_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n48469), .I2(n52716), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5430));
    defparam select_775_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h9600;
    SB_LUT4 i2_3_lut_4_lut_adj_1456 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3][2] ), .I3(\data_in_frame[1] [1]), .O(n52871));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 n62493_bdd_4_lut (.I0(n62493), .I1(n56712), .I2(n56711), .I3(\byte_transmit_counter[2] ), 
            .O(n62496));
    defparam n62493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2][7] ), 
            .I2(n23220), .I3(GND_net), .O(n23534));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_213_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n48469), .I2(n52632), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5429));
    defparam select_775_Select_213_i3_3_lut_4_lut.LUT_INIT = 16'h6900;
    SB_LUT4 i3_3_lut_4_lut_adj_1458 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n48494), .I3(\data_out_frame[23] [4]), .O(n8_adj_5584));
    defparam i3_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(\data_out_frame[25] [3]), .I1(n48603), 
            .I2(GND_net), .I3(GND_net), .O(n48611));
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i13717_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n27423));   // verilog/coms.v(130[12] 305[6])
    defparam i13717_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_220_i3_4_lut (.I0(n2394), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[25] [2]), .I3(n48611), .O(n3_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_220_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13917_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [7]), 
            .I3(current_limit[7]), .O(n27623));   // verilog/coms.v(130[12] 305[6])
    defparam i13917_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13716_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n27422));   // verilog/coms.v(130[12] 305[6])
    defparam i13716_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_219_i3_3_lut (.I0(n52552), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n52957), .I3(GND_net), .O(n3_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_219_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n52683), .I3(GND_net), .O(n6_adj_5585));
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i13708_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n27414));   // verilog/coms.v(130[12] 305[6])
    defparam i13708_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n52665), .I3(n48441), .O(n3_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(\data_out_frame[20] [6]), .I1(n48587), 
            .I2(GND_net), .I3(GND_net), .O(n53143));
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1462 (.I0(n2342), .I1(\data_out_frame[16] [6]), 
            .I2(n52892), .I3(\data_out_frame[18] [4]), .O(n54351));
    defparam i3_4_lut_adj_1462.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1463 (.I0(n53023), .I1(n53104), .I2(n54351), 
            .I3(n52860), .O(n12_adj_5586));
    defparam i5_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1464 (.I0(n53167), .I1(n12_adj_5586), .I2(\data_out_frame[16] [1]), 
            .I3(n53143), .O(n48523));
    defparam i6_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1465 (.I0(n53143), .I1(n52761), .I2(n47428), 
            .I3(n52825), .O(n14_adj_5587));
    defparam i6_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1466 (.I0(n53149), .I1(n14_adj_5587), .I2(n10_adj_5572), 
            .I3(\data_out_frame[16] [3]), .O(n2394));
    defparam i7_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1467 (.I0(\data_out_frame[23] [0]), .I1(n48523), 
            .I2(GND_net), .I3(GND_net), .O(n48441));
    defparam i1_2_lut_adj_1467.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1468 (.I0(\data_out_frame[22] [6]), .I1(n23185), 
            .I2(\data_out_frame[24] [7]), .I3(n53046), .O(n10_adj_5571));
    defparam i4_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n52506), .I3(\data_in_frame[1] [0]), .O(n23220));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(n48629), .I1(n48474), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5583));
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1471 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5588));
    defparam i1_2_lut_adj_1471.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1472 (.I0(\data_out_frame[16] [4]), .I1(n47581), 
            .I2(\data_out_frame[22] [7]), .I3(n6_adj_5588), .O(n52761));
    defparam i4_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1473 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(n52761), .I3(GND_net), .O(n14_adj_5589));
    defparam i5_3_lut_adj_1473.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1474 (.I0(n53107), .I1(\data_out_frame[23] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(n52892), .O(n15_adj_5590));
    defparam i6_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1475 (.I0(n15_adj_5590), .I1(n52598), .I2(n14_adj_5589), 
            .I3(n48587), .O(n48603));
    defparam i8_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i20443_3_lut_4_lut (.I0(deadband[5]), .I1(\data_in_frame[16]_c [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27125));
    defparam i20443_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i3_3_lut_adj_1476 (.I0(n48499), .I1(n48603), .I2(n52764), 
            .I3(GND_net), .O(n8_adj_5591));
    defparam i3_3_lut_adj_1476.LUT_INIT = 16'h6969;
    SB_LUT4 select_775_Select_217_i3_4_lut (.I0(n48471), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5591), .I3(n52552), .O(n3_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_adj_1477 (.I0(n54349), .I1(\data_out_frame[24] [6]), 
            .I2(\data_out_frame[25] [0]), .I3(GND_net), .O(n52665));
    defparam i2_3_lut_adj_1477.LUT_INIT = 16'h6969;
    SB_LUT4 i13707_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n27413));   // verilog/coms.v(130[12] 305[6])
    defparam i13707_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_216_i3_3_lut (.I0(n52665), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n53003), .I3(GND_net), .O(n3_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52957));
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i13706_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n27412));   // verilog/coms.v(130[12] 305[6])
    defparam i13706_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13920_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [4]), 
            .I3(current_limit[4]), .O(n27626));   // verilog/coms.v(130[12] 305[6])
    defparam i13920_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1479 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [3]), 
            .I2(n52957), .I3(n6_adj_5585), .O(n48471));
    defparam i4_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(n23713), .I1(n48471), .I2(GND_net), 
            .I3(GND_net), .O(n53003));
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_215_i3_4_lut (.I0(n52716), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n53003), .I3(\data_out_frame[25] [0]), .O(n3_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i21608_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n26918));   // verilog/coms.v(130[12] 305[6])
    defparam i21608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47575 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56669), .I2(n56670), .I3(\byte_transmit_counter[2] ), 
            .O(n62487));
    defparam byte_transmit_counter_1__bdd_4_lut_47575.LUT_INIT = 16'he4aa;
    SB_LUT4 i13911_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [5]), 
            .I3(current_limit[13]), .O(n27617));   // verilog/coms.v(130[12] 305[6])
    defparam i13911_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13705_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n27411));   // verilog/coms.v(130[12] 305[6])
    defparam i13705_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13916_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [0]), 
            .I3(current_limit[8]), .O(n27622));   // verilog/coms.v(130[12] 305[6])
    defparam i13916_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13704_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n27410));   // verilog/coms.v(130[12] 305[6])
    defparam i13704_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i45370_2_lut (.I0(n62628), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59336));
    defparam i45370_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13703_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n27409));   // verilog/coms.v(130[12] 305[6])
    defparam i13703_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13702_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n27408));   // verilog/coms.v(130[12] 305[6])
    defparam i13702_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_212_i3_3_lut (.I0(n52632), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n52810), .I3(GND_net), .O(n3_adj_5428));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_212_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i44926_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59293));   // verilog/coms.v(158[12:15])
    defparam i44926_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46099_3_lut (.I0(n62562), .I1(n62514), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n60999));
    defparam i46099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(\data_out_frame[24] [2]), .I1(n22527), 
            .I2(GND_net), .I3(GND_net), .O(n52810));
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 select_775_Select_211_i3_4_lut (.I0(n21093), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n52810), .I3(\data_out_frame[24] [1]), .O(n3_adj_5427));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i23343_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_10), .I3(n15_adj_11), .O(\motor_state_23__N_67[17] ));
    defparam i23343_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13701_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n27407));   // verilog/coms.v(130[12] 305[6])
    defparam i13701_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1482 (.I0(n52686), .I1(n21093), .I2(\data_out_frame[24] [0]), 
            .I3(n53011), .O(n10_adj_5594));
    defparam i4_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_210_i3_4_lut (.I0(n23699), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5594), .I3(\data_out_frame[21] [6]), .O(n3_adj_5426));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_2_lut_adj_1483 (.I0(n23713), .I1(\data_out_frame[24] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5595));
    defparam i2_2_lut_adj_1483.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1484 (.I0(n7_adj_5595), .I1(n23185), .I2(\data_out_frame[25] [7]), 
            .I3(n48525), .O(n52683));
    defparam i4_4_lut_adj_1484.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\data_out_frame[20] [4]), .I1(n54473), 
            .I2(GND_net), .I3(GND_net), .O(n52860));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h9999;
    SB_LUT4 select_777_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1486 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2487 ), 
            .I2(\FRAME_MATCHER.i_31__N_2490 ), .I3(GND_net), .O(n52403));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1486.LUT_INIT = 16'hfefe;
    SB_LUT4 select_777_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(byte_transmit_counter[5]), 
            .I3(GND_net), .O(n1_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_adj_1487 (.I0(\data_out_frame[19] [5]), .I1(n48452), 
            .I2(n47856), .I3(GND_net), .O(n23699));
    defparam i2_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1488 (.I0(n2217), .I1(n52932), .I2(n52520), .I3(n23699), 
            .O(n48247));
    defparam i3_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i13930_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n27636));   // verilog/coms.v(130[12] 305[6])
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_777_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(byte_transmit_counter[6]), 
            .I3(GND_net), .O(n1_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_777_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(byte_transmit_counter[7]), 
            .I3(GND_net), .O(n1_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_777_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(\byte_transmit_counter[4] ), 
            .I3(GND_net), .O(n1_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_777_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(\byte_transmit_counter[3] ), 
            .I3(GND_net), .O(n1_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_777_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n1_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 n62487_bdd_4_lut (.I0(n62487), .I1(n56709), .I2(n56708), .I3(\byte_transmit_counter[2] ), 
            .O(n62490));
    defparam n62487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i23395_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n27632));   // verilog/coms.v(130[12] 305[6])
    defparam i23395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_777_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2487 ), .I2(\byte_transmit_counter[1] ), 
            .I3(GND_net), .O(n1_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52478));
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'h6666;
    SB_LUT4 i13921_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [3]), 
            .I3(current_limit[3]), .O(n27627));   // verilog/coms.v(130[12] 305[6])
    defparam i13921_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13919_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [5]), 
            .I3(current_limit[5]), .O(n27625));   // verilog/coms.v(130[12] 305[6])
    defparam i13919_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1490 (.I0(n52598), .I1(\data_out_frame[20] [2]), 
            .I2(\data_out_frame[20] [4]), .I3(n52478), .O(n2217));
    defparam i3_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1491 (.I0(\data_out_frame[23] [7]), .I1(n52854), 
            .I2(\data_out_frame[19] [5]), .I3(\data_out_frame[21] [7]), 
            .O(n13_adj_5596));
    defparam i5_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1492 (.I0(n13_adj_5596), .I1(n11_adj_5570), .I2(\data_out_frame[21] [5]), 
            .I3(n52808), .O(n21093));
    defparam i7_4_lut_adj_1492.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1493 (.I0(n2054), .I1(n52808), .I2(n48247), .I3(n47968), 
            .O(n16_adj_5597));
    defparam i6_4_lut_adj_1493.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1494 (.I0(n52709), .I1(n48527), .I2(\data_out_frame[22] [1]), 
            .I3(n2217), .O(n17_adj_5598));
    defparam i7_4_lut_adj_1494.LUT_INIT = 16'h9669;
    SB_LUT4 i13928_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n27634));   // verilog/coms.v(130[12] 305[6])
    defparam i13928_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_4_lut_adj_1495 (.I0(n17_adj_5598), .I1(n21050), .I2(n16_adj_5597), 
            .I3(n54473), .O(n22527));
    defparam i9_4_lut_adj_1495.LUT_INIT = 16'h9669;
    SB_LUT4 i13925_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n27631));   // verilog/coms.v(130[12] 305[6])
    defparam i13925_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1496 (.I0(\data_out_frame[22] [3]), .I1(n53101), 
            .I2(n52991), .I3(\data_out_frame[20] [0]), .O(n48469));
    defparam i3_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i13700_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n27406));   // verilog/coms.v(130[12] 305[6])
    defparam i13700_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1497 (.I0(n48463), .I1(n47422), .I2(n23967), 
            .I3(n6_adj_5573), .O(n2054));
    defparam i4_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_out_frame[20] [2]), .I1(n2054), 
            .I2(GND_net), .I3(GND_net), .O(n52991));
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1499 (.I0(\data_out_frame[18] [5]), .I1(n53024), 
            .I2(n52862), .I3(n23455), .O(n10_adj_5599));
    defparam i4_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1500 (.I0(n24097), .I1(n10_adj_5599), .I2(\data_out_frame[17] [0]), 
            .I3(GND_net), .O(n53104));
    defparam i5_3_lut_adj_1500.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1501 (.I0(n52721), .I1(n52935), .I2(GND_net), 
            .I3(GND_net), .O(n53107));
    defparam i1_2_lut_adj_1501.LUT_INIT = 16'h6666;
    SB_LUT4 i13914_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [2]), 
            .I3(current_limit[10]), .O(n27620));   // verilog/coms.v(130[12] 305[6])
    defparam i13914_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13927_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n27633));   // verilog/coms.v(130[12] 305[6])
    defparam i13927_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47570 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56699), .I2(n56700), .I3(\byte_transmit_counter[2] ), 
            .O(n62481));
    defparam byte_transmit_counter_1__bdd_4_lut_47570.LUT_INIT = 16'he4aa;
    SB_LUT4 i13912_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[20] [4]), 
            .I3(current_limit[12]), .O(n27618));   // verilog/coms.v(130[12] 305[6])
    defparam i13912_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52758));
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n23967));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1504 (.I0(n23967), .I1(\data_out_frame[17] [3]), 
            .I2(n24203), .I3(\data_out_frame[17] [1]), .O(n16_adj_5600));   // verilog/coms.v(79[16:43])
    defparam i6_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1505 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[16] [5]), 
            .I2(n52604), .I3(\data_out_frame[17] [2]), .O(n17_adj_5601));   // verilog/coms.v(79[16:43])
    defparam i7_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1506 (.I0(n17_adj_5601), .I1(\data_out_frame[17] [4]), 
            .I2(n16_adj_5600), .I3(n62162), .O(n54016));   // verilog/coms.v(79[16:43])
    defparam i9_4_lut_adj_1506.LUT_INIT = 16'h9669;
    SB_LUT4 i47266_4_lut (.I0(n54016), .I1(\data_out_frame[18] [5]), .I2(n52864), 
            .I3(\data_out_frame[14] [4]), .O(n62166));
    defparam i47266_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1507 (.I0(n52587), .I1(n52758), .I2(n62166), 
            .I3(\data_out_frame[14] [5]), .O(n24_adj_5602));
    defparam i9_4_lut_adj_1507.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1508 (.I0(n52564), .I1(n47944), .I2(n23754), 
            .I3(\data_out_frame[19] [3]), .O(n26_adj_5603));
    defparam i11_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i13213_3_lut_4_lut (.I0(n2978), .I1(n25012), .I2(\data_in_frame[21] [0]), 
            .I3(current_limit[0]), .O(n26919));   // verilog/coms.v(130[12] 305[6])
    defparam i13213_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut_adj_1509 (.I0(n23155), .I1(n52794), .I2(n2076), 
            .I3(n52712), .O(n25_adj_5604));
    defparam i10_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1510 (.I0(\data_out_frame[19] [4]), .I1(n24_adj_5602), 
            .I2(n53052), .I3(n47720), .O(n27_c));
    defparam i12_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1511 (.I0(n27_c), .I1(n53107), .I2(n25_adj_5604), 
            .I3(n26_adj_5603), .O(n6_adj_5605));
    defparam i1_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1512 (.I0(n23964), .I1(\data_out_frame[19] [5]), 
            .I2(n53104), .I3(n6_adj_5605), .O(n21050));
    defparam i4_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(\data_out_frame[20] [0]), .I1(n21050), 
            .I2(GND_net), .I3(GND_net), .O(n52932));
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_out_frame[19] [6]), .I1(n53026), 
            .I2(GND_net), .I3(GND_net), .O(n52794));
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1515 (.I0(\data_out_frame[17] [6]), .I1(n52794), 
            .I2(n47856), .I3(\data_out_frame[22] [2]), .O(n53101));
    defparam i3_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53149));
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1517 (.I0(\data_in_frame[2] [0]), .I1(n23706), 
            .I2(n53020), .I3(GND_net), .O(n53000));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1517.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1518 (.I0(\data_out_frame[21] [7]), .I1(n53101), 
            .I2(\data_out_frame[22] [1]), .I3(n48568), .O(n10_adj_5569));
    defparam i4_4_lut_adj_1518.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1519 (.I0(n1699), .I1(n53035), .I2(n52601), .I3(n54100), 
            .O(n48587));
    defparam i3_4_lut_adj_1519.LUT_INIT = 16'h9669;
    SB_LUT4 i13699_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n27405));   // verilog/coms.v(130[12] 305[6])
    defparam i13699_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1520 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23568));
    defparam i1_2_lut_adj_1520.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52935));
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i13698_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n27404));   // verilog/coms.v(130[12] 305[6])
    defparam i13698_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1522 (.I0(\data_out_frame[21] [0]), .I1(n52935), 
            .I2(n23568), .I3(\data_out_frame[16] [4]), .O(n10_adj_5567));
    defparam i4_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1523 (.I0(n52520), .I1(n10_adj_5567), .I2(n52892), 
            .I3(GND_net), .O(n47428));
    defparam i5_3_lut_adj_1523.LUT_INIT = 16'h6969;
    SB_LUT4 i13173_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[10][7] ), .O(n26879));
    defparam i13173_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13170_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n26876));
    defparam i13170_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n62481_bdd_4_lut (.I0(n62481), .I1(n56703), .I2(n56702), .I3(\byte_transmit_counter[2] ), 
            .O(n62484));
    defparam n62481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13161_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[10][3] ), .O(n26867));
    defparam i13161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13158_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[10][2] ), .O(n26864));
    defparam i13158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1524 (.I0(n48629), .I1(\data_out_frame[23] [3]), 
            .I2(n4_adj_5568), .I3(GND_net), .O(n48499));
    defparam i1_3_lut_adj_1524.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(n54100), .I1(n52705), .I2(GND_net), 
            .I3(GND_net), .O(n53023));
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h9999;
    SB_LUT4 i13697_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n27403));   // verilog/coms.v(130[12] 305[6])
    defparam i13697_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13696_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n27402));   // verilog/coms.v(130[12] 305[6])
    defparam i13696_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23155));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1527 (.I0(n23041), .I1(n52481), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n47856));
    defparam i2_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i13155_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[10][1] ), .O(n26861));
    defparam i13155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13152_3_lut_4_lut (.I0(n25707), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[10][0] ), .O(n26858));
    defparam i13152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1528 (.I0(n47720), .I1(\data_out_frame[22] [0]), 
            .I2(\data_out_frame[19] [6]), .I3(GND_net), .O(n53075));
    defparam i2_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1529 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52864));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1529.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1530 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n47527), .I3(GND_net), .O(n47581));
    defparam i2_3_lut_adj_1530.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[16] [1]), .I1(n47581), 
            .I2(GND_net), .I3(GND_net), .O(n52773));
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1532 (.I0(n1835), .I1(n52864), .I2(n23601), .I3(n47380), 
            .O(n53078));
    defparam i3_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1533 (.I0(n52674), .I1(n23601), .I2(n47944), 
            .I3(n24120), .O(n10_adj_5606));
    defparam i4_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1534 (.I0(\data_out_frame[15] [7]), .I1(n10_adj_5606), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n48463));
    defparam i5_3_lut_adj_1534.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1535 (.I0(n48463), .I1(n53078), .I2(n52773), 
            .I3(\data_out_frame[18] [1]), .O(n48527));
    defparam i3_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1536 (.I0(n47641), .I1(n48494), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n23713));
    defparam i2_3_lut_adj_1536.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\data_out_frame[20] [3]), .I1(n48527), 
            .I2(GND_net), .I3(GND_net), .O(n52627));
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1538 (.I0(\data_out_frame[23] [7]), .I1(\data_out_frame[24] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53011));
    defparam i1_2_lut_adj_1538.LUT_INIT = 16'h6666;
    SB_LUT4 i13695_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n27401));   // verilog/coms.v(130[12] 305[6])
    defparam i13695_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1539 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [3]), 
            .I2(n52452), .I3(n6_adj_5566), .O(n1673));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1540 (.I0(\data_out_frame[11] [0]), .I1(n52475), 
            .I2(n52979), .I3(n1673), .O(n18_adj_5607));
    defparam i7_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1541 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[4] [6]), .O(n52458));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1542 (.I0(n53083), .I1(n52614), .I2(n52928), 
            .I3(\data_out_frame[8] [2]), .O(n19));
    defparam i8_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i13694_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n27400));   // verilog/coms.v(130[12] 305[6])
    defparam i13694_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_4_lut_adj_1543 (.I0(n19), .I1(n22437), .I2(n17_adj_5565), 
            .I3(n18_adj_5607), .O(n10_adj_5608));
    defparam i2_4_lut_adj_1543.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1544 (.I0(n52779), .I1(n1510), .I2(n23437), .I3(\data_out_frame[13] [7]), 
            .O(n14_adj_5609));
    defparam i6_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1545 (.I0(n1513), .I1(n14_adj_5609), .I2(n10_adj_5608), 
            .I3(n1673), .O(n54100));
    defparam i7_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1546 (.I0(n54100), .I1(n52862), .I2(GND_net), 
            .I3(GND_net), .O(n52825));
    defparam i1_2_lut_adj_1546.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1547 (.I0(n53043), .I1(\data_out_frame[18] [6]), 
            .I2(n52822), .I3(\data_out_frame[20] [7]), .O(n14_adj_5610));
    defparam i6_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1548 (.I0(\data_out_frame[21] [1]), .I1(n14_adj_5610), 
            .I2(n10_adj_5564), .I3(\data_out_frame[16] [7]), .O(n48474));
    defparam i7_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i1554_2_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2342));   // verilog/coms.v(81[16:27])
    defparam i1554_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1549 (.I0(n23041), .I1(n23594), .I2(\data_out_frame[15] [3]), 
            .I3(\data_out_frame[17] [5]), .O(n52712));
    defparam i3_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1550 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6][7] ), 
            .I2(\data_in_frame[6][6] ), .I3(GND_net), .O(n52948));
    defparam i1_2_lut_3_lut_adj_1550.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1551 (.I0(\data_out_frame[19] [7]), .I1(n47380), 
            .I2(n52555), .I3(n23041), .O(n53026));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(\data_out_frame[18] [0]), .I1(n53026), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5611));
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1553 (.I0(\data_out_frame[17] [7]), .I1(n47422), 
            .I2(n52712), .I3(n6_adj_5611), .O(n47968));
    defparam i4_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1554 (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[22] [4]), 
            .I2(n47968), .I3(GND_net), .O(n54449));
    defparam i2_3_lut_adj_1554.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1555 (.I0(\data_out_frame[21] [6]), .I1(n53075), 
            .I2(n47856), .I3(n48240), .O(n52709));
    defparam i3_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1556 (.I0(n2342), .I1(\data_out_frame[20] [1]), 
            .I2(n48474), .I3(\data_out_frame[20] [6]), .O(n55042));
    defparam i3_4_lut_adj_1556.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1557 (.I0(n48601), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[24] [3]), .I3(n52709), .O(n54735));
    defparam i3_4_lut_adj_1557.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1558 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[23] [1]), 
            .I2(\data_out_frame[24] [7]), .I3(n48499), .O(n28_adj_5612));
    defparam i12_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i13693_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n27399));   // verilog/coms.v(130[12] 305[6])
    defparam i13693_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1559 (.I0(n53011), .I1(n52627), .I2(n23713), 
            .I3(n55042), .O(n26_adj_5613));
    defparam i10_4_lut_adj_1559.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1560 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(n54449), .I3(\data_out_frame[24] [6]), .O(n27_adj_5614));
    defparam i11_4_lut_adj_1560.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1561 (.I0(n54735), .I1(n52776), .I2(n53149), 
            .I3(n53008), .O(n25_adj_5615));
    defparam i9_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1562 (.I0(n25_adj_5615), .I1(n27_adj_5614), .I2(n26_adj_5613), 
            .I3(n28_adj_5612), .O(n48525));
    defparam i15_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1563 (.I0(n52776), .I1(n53046), .I2(n48247), 
            .I3(GND_net), .O(n2329));
    defparam i2_3_lut_adj_1563.LUT_INIT = 16'h9696;
    SB_LUT4 i13710_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n27416));   // verilog/coms.v(130[12] 305[6])
    defparam i13710_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1564 (.I0(n48469), .I1(n54349), .I2(n22527), 
            .I3(n21093), .O(n55052));
    defparam i3_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1565 (.I0(n52683), .I1(n55052), .I2(n21097), 
            .I3(GND_net), .O(n8_adj_5616));
    defparam i3_3_lut_adj_1565.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_209_i3_4_lut (.I0(n2329), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5616), .I3(n48525), .O(n3_adj_5425));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_209_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_2_lut_3_lut_adj_1566 (.I0(\data_in_frame[8][7] ), .I1(\data_in_frame[4] [5]), 
            .I2(n52595), .I3(GND_net), .O(n7_adj_5531));
    defparam i2_2_lut_3_lut_adj_1566.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1567 (.I0(\data_out_frame[19] [3]), .I1(n53040), 
            .I2(GND_net), .I3(GND_net), .O(n52854));
    defparam i1_2_lut_adj_1567.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53008));
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1569 (.I0(\data_in_frame[2] [5]), .I1(n52463), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[7] [0]), .O(n52900));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1569.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1570 (.I0(\data_in_frame[16] [6]), .I1(n54734), 
            .I2(\data_in_frame[19] [0]), .I3(n54381), .O(n52886));
    defparam i2_3_lut_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1571 (.I0(n47797), .I1(\data_in_frame[9] [7]), 
            .I2(Kp_23__N_675), .I3(n23812), .O(n14_adj_5507));
    defparam i5_3_lut_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1572 (.I0(n48308), .I1(n23594), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5617));
    defparam i1_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1573 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_5617), .O(n48452));
    defparam i4_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1574 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [4]), .I3(n47475), .O(n52997));
    defparam i1_2_lut_4_lut_adj_1574.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1575 (.I0(n47456), .I1(n53032), .I2(\data_out_frame[17] [2]), 
            .I3(GND_net), .O(n52523));
    defparam i2_3_lut_adj_1575.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(\data_out_frame[19] [3]), .I1(n52523), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5618));
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1577 (.I0(\data_out_frame[21] [4]), .I1(n23964), 
            .I2(n24203), .I3(n6_adj_5618), .O(n47641));
    defparam i4_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1578 (.I0(\data_in_frame[13] [0]), .I1(n23367), 
            .I2(n24073), .I3(GND_net), .O(n6_adj_5502));
    defparam i1_2_lut_3_lut_adj_1578.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1579 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[12] [6]), 
            .I2(n52966), .I3(\data_out_frame[8] [4]), .O(n16_adj_5619));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1580 (.I0(\data_out_frame[4] [1]), .I1(n52484), 
            .I2(n53122), .I3(\data_out_frame[5] [5]), .O(n17_adj_5620));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1581 (.I0(n17_adj_5620), .I1(\data_out_frame[5] [6]), 
            .I2(n16_adj_5619), .I3(\data_out_frame[10] [3]), .O(n48308));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n23613));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1583 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[11] [7]), 
            .I2(n23639), .I3(n23797), .O(n52831));
    defparam i2_3_lut_4_lut_adj_1583.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1584 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[14] [5]), 
            .I2(n48308), .I3(\data_out_frame[15] [0]), .O(n10_adj_5621));
    defparam i4_4_lut_adj_1584.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1585 (.I0(n1655), .I1(n10_adj_5621), .I2(\data_out_frame[16] [7]), 
            .I3(GND_net), .O(n53040));
    defparam i5_3_lut_adj_1585.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1586 (.I0(n47502), .I1(n7_adj_5581), .I2(n2076), 
            .I3(GND_net), .O(n52822));
    defparam i2_3_lut_adj_1586.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1587 (.I0(n22568), .I1(\data_in_frame[13][7] ), 
            .I2(\data_in_frame[13][6] ), .I3(GND_net), .O(n52972));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1587.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1588 (.I0(n53098), .I1(n53158), .I2(\data_out_frame[11] [7]), 
            .I3(GND_net), .O(n22437));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1588.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1589 (.I0(n22437), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[12] [1]), .I3(GND_net), .O(n53052));
    defparam i2_3_lut_adj_1589.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_3_lut (.I0(reset), .I1(\FRAME_MATCHER.i[0] ), .I2(n38302), 
            .I3(GND_net), .O(n68));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_adj_1590 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52614));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1590.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1591 (.I0(n52614), .I1(n47380), .I2(\data_out_frame[15] [5]), 
            .I3(n52963), .O(n10_adj_5563));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1591.LUT_INIT = 16'h6996;
    SB_LUT4 i44551_2_lut (.I0(\data_out_frame[0][2] ), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n59351));
    defparam i44551_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13369_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n27075));
    defparam i13369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(\data_out_frame[16] [5]), .I1(n52587), 
            .I2(GND_net), .I3(GND_net), .O(n23263));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1593 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23754));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1593.LUT_INIT = 16'h6666;
    SB_LUT4 i13366_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n27072));
    defparam i13366_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i41734_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56634));
    defparam i41734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1594 (.I0(n8_adj_5506), .I1(n10), .I2(n38302), 
            .I3(GND_net), .O(n25721));
    defparam i1_2_lut_3_lut_adj_1594.LUT_INIT = 16'hefef;
    SB_LUT4 i3_4_lut_adj_1595 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(n23754), .I3(n23263), .O(n52674));
    defparam i3_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i13363_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n27069));
    defparam i13363_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1596 (.I0(n23367), .I1(n22568), .I2(\data_in_frame[15] [7]), 
            .I3(n23135), .O(n47517));
    defparam i2_3_lut_4_lut_adj_1596.LUT_INIT = 16'h6996;
    SB_LUT4 i41735_4_lut (.I0(n56634), .I1(n59351), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n56635));
    defparam i41735_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i47262_3_lut (.I0(n47502), .I1(n52862), .I2(n47944), .I3(GND_net), 
            .O(n62162));
    defparam i47262_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i41733_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n56633));
    defparam i41733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13360_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n27066));
    defparam i13360_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13357_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n27063));
    defparam i13357_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13329_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n27035));
    defparam i13329_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_4_lut_adj_1597 (.I0(\data_in_frame[16]_c [5]), .I1(n13_adj_5512), 
            .I2(\data_in_frame[14] [3]), .I3(n14_adj_5511), .O(n52819));
    defparam i2_2_lut_4_lut_adj_1597.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1598 (.I0(\data_in_frame[15] [5]), .I1(n10_adj_5489), 
            .I2(n52678), .I3(\data_in_frame[18] [1]), .O(n52659));
    defparam i1_2_lut_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1599 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n52555));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1599.LUT_INIT = 16'h6666;
    SB_LUT4 i13326_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n27032));
    defparam i13326_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13323_3_lut_4_lut (.I0(n37), .I1(n52424), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n27029));
    defparam i13323_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1600 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n52897));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1600.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1601 (.I0(\data_out_frame[8] [4]), .I1(n53083), 
            .I2(n52489), .I3(n52894), .O(n12_adj_5622));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1601.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1602 (.I0(\data_out_frame[4] [2]), .I1(n12_adj_5622), 
            .I2(\data_out_frame[13] [0]), .I3(n52897), .O(n47456));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1602.LUT_INIT = 16'h6996;
    SB_LUT4 i45231_2_lut (.I0(n62598), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59386));
    defparam i45231_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1603 (.I0(n47456), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n52481));
    defparam i2_3_lut_adj_1603.LUT_INIT = 16'h9696;
    SB_LUT4 i11651_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n25356));   // verilog/coms.v(109[34:55])
    defparam i11651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1604 (.I0(\data_out_frame[9] [1]), .I1(n23758), 
            .I2(GND_net), .I3(GND_net), .O(n52963));
    defparam i1_2_lut_adj_1604.LUT_INIT = 16'h6666;
    SB_LUT4 i13863_3_lut_4_lut (.I0(n25705), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n27569));
    defparam i13863_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1605 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n24002));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1605.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1606 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[7] [1]), .O(n26_adj_5623));   // verilog/coms.v(75[16:27])
    defparam i11_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1607 (.I0(n52484), .I1(n52647), .I2(\data_out_frame[8] [3]), 
            .I3(\data_out_frame[4] [5]), .O(n24_adj_5624));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut_adj_1607.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1608 (.I0(n44537), .I1(n52922), .I2(n23577), 
            .I3(n52641), .O(n25_adj_5625));   // verilog/coms.v(75[16:27])
    defparam i10_4_lut_adj_1608.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n56668), .I1(n56666), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[0] ), 
            .O(n7_adj_5270));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i14_4_lut_adj_1609 (.I0(n23_adj_5578), .I1(n25_adj_5625), .I2(n24_adj_5624), 
            .I3(n26_adj_5623), .O(n54139));   // verilog/coms.v(75[16:27])
    defparam i14_4_lut_adj_1609.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1610 (.I0(n52567), .I1(n52963), .I2(n23434), 
            .I3(n54139), .O(n12_adj_5626));
    defparam i5_4_lut_adj_1610.LUT_INIT = 16'h6996;
    SB_LUT4 i13569_3_lut_4_lut (.I0(n25705), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n27275));
    defparam i13569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1611 (.I0(\data_out_frame[7] [5]), .I1(n12_adj_5626), 
            .I2(n53069), .I3(\data_out_frame[9] [5]), .O(n54459));
    defparam i6_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1612 (.I0(n24002), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[11] [6]), .I3(n54459), .O(n12_adj_5627));
    defparam i5_4_lut_adj_1612.LUT_INIT = 16'h9669;
    SB_LUT4 i44742_2_lut (.I0(n62610), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59337));
    defparam i44742_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1613 (.I0(n23758), .I1(n12_adj_5627), .I2(\data_out_frame[11] [7]), 
            .I3(\data_out_frame[11] [4]), .O(n52979));
    defparam i6_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46117_3_lut (.I0(n62556), .I1(n62508), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n61017));
    defparam i46117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(\data_out_frame[14] [1]), .I1(n52513), 
            .I2(n12), .I3(n8), .O(n52779));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1615 (.I0(n47380), .I1(n24120), .I2(GND_net), 
            .I3(GND_net), .O(n47414));
    defparam i1_2_lut_adj_1615.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1616 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52484));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1616.LUT_INIT = 16'h6666;
    SB_LUT4 i13560_3_lut_4_lut (.I0(n25705), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n27266));
    defparam i13560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13557_3_lut_4_lut (.I0(n25705), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n27263));
    defparam i13557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13554_3_lut_4_lut (.I0(n25705), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n27260));
    defparam i13554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13597_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n27303));
    defparam i13597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11641_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n25346));   // verilog/coms.v(109[34:55])
    defparam i11641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1617 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52500));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1617.LUT_INIT = 16'h6666;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1618 (.I0(\data_out_frame[6] [3]), .I1(n52489), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n23758));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1618.LUT_INIT = 16'h9696;
    SB_LUT4 i13594_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n27300));
    defparam i13594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1619 (.I0(\data_in_frame[15] [0]), .I1(n23824), 
            .I2(n53055), .I3(GND_net), .O(n10_adj_5467));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_3_lut_adj_1619.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1620 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[14] [7]), .I3(n53064), .O(n6_adj_5465));
    defparam i1_2_lut_4_lut_adj_1620.LUT_INIT = 16'h6996;
    SB_LUT4 i13591_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n27297));
    defparam i13591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1621 (.I0(n23758), .I1(n32), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n52939));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53119));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1623 (.I0(n23313), .I1(n24073), .I2(\data_in_frame[14] [7]), 
            .I3(n23821), .O(n52788));
    defparam i2_3_lut_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1624 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[11] [0]), .I3(\data_out_frame[10] [6]), 
            .O(n10_adj_5630));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1624.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1625 (.I0(n23577), .I1(n10_adj_5630), .I2(n23012), 
            .I3(GND_net), .O(n52529));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_adj_1625.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1626 (.I0(n53110), .I1(n52529), .I2(n23688), 
            .I3(n53119), .O(n10_adj_5631));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1627 (.I0(n52939), .I1(n10_adj_5631), .I2(n44537), 
            .I3(GND_net), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_adj_1627.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1628 (.I0(\data_in_frame[20] [0]), .I1(\data_in_frame[18] [5]), 
            .I2(\data_in_frame[20] [6]), .I3(n52886), .O(n21));
    defparam i2_2_lut_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1629 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [6]), 
            .I2(n52886), .I3(GND_net), .O(n52668));
    defparam i1_2_lut_3_lut_adj_1629.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1630 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23434));
    defparam i1_2_lut_adj_1630.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1631 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[18]_c [6]), 
            .I2(n55049), .I3(n52532), .O(n53072));
    defparam i2_3_lut_4_lut_adj_1631.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1632 (.I0(n23869), .I1(n22594), .I2(n23434), 
            .I3(n1312), .O(n52851));
    defparam i3_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1633 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n52647));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1633.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1634 (.I0(\data_out_frame[5] [5]), .I1(n52647), 
            .I2(n1191), .I3(n23005), .O(n1168));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1634.LUT_INIT = 16'h6996;
    SB_LUT4 i13588_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n27294));
    defparam i13588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1635 (.I0(\data_in_frame[13][5] ), .I1(n23313), 
            .I2(n10_adj_5411), .I3(\data_in_frame[18] [0]), .O(n53164));   // verilog/coms.v(78[16:43])
    defparam i5_3_lut_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1636 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n23945));
    defparam i2_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1637 (.I0(n23945), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n53110));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1637.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1638 (.I0(n23688), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n52741));
    defparam i2_3_lut_adj_1638.LUT_INIT = 16'h9696;
    SB_LUT4 i13585_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n27291));
    defparam i13585_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13581_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n27287));
    defparam i13581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(\data_out_frame[7] [1]), .I1(n23427), 
            .I2(GND_net), .I3(GND_net), .O(n23869));
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1640 (.I0(\data_in_frame[21] [4]), .I1(n47491), 
            .I2(n52813), .I3(GND_net), .O(n52770));
    defparam i1_2_lut_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1641 (.I0(n52741), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[13] [5]), .I3(n53110), .O(n10_adj_5574));
    defparam i4_4_lut_adj_1641.LUT_INIT = 16'h6996;
    SB_LUT4 i13578_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n27284));
    defparam i13578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47585 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n62475));
    defparam byte_transmit_counter_0__bdd_4_lut_47585.LUT_INIT = 16'he4aa;
    SB_LUT4 i13575_3_lut_4_lut (.I0(n35699), .I1(n52434), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n27281));
    defparam i13575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1642 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_9));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_adj_1642.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1643 (.I0(n23500), .I1(\data_in_frame[16] [3]), 
            .I2(n22606), .I3(GND_net), .O(n47264));
    defparam i1_2_lut_3_lut_adj_1643.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1644 (.I0(n23410), .I1(n53128), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n52601));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1644.LUT_INIT = 16'h9696;
    SB_LUT4 i13234_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n26940));
    defparam i13234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1645 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n52662));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1645.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1646 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(n52466), .I3(n53152), .O(n23283));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1647 (.I0(reset), .I1(n52409), .I2(\FRAME_MATCHER.i[1] ), 
            .I3(\FRAME_MATCHER.i[0] ), .O(n54720));
    defparam i3_4_lut_adj_1647.LUT_INIT = 16'hffef;
    SB_LUT4 i13231_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n26937));
    defparam i13231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1648 (.I0(\data_in_frame[9] [3]), .I1(n24061), 
            .I2(n47797), .I3(n53017), .O(n52985));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1649 (.I0(\data_in_frame[9] [3]), .I1(n24061), 
            .I2(\data_in_frame[11] [4]), .I3(\data_in_frame[9] [2]), .O(n23313));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1650 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n23005));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1650.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n203), .I1(n151), .I2(n204), 
            .I3(GND_net), .O(n6));
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i45312_3_lut_4_lut (.I0(n203), .I1(n151), .I2(n204), .I3(n152), 
            .O(n60212));
    defparam i45312_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i2_3_lut_adj_1651 (.I0(n1312), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n53128));
    defparam i2_3_lut_adj_1651.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1652 (.I0(\data_in_frame[0][7] ), .I1(n23238), 
            .I2(n23251), .I3(\data_in_frame[3][3] ), .O(n21154));
    defparam i2_3_lut_4_lut_adj_1652.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1653 (.I0(\data_in_frame[0][7] ), .I1(n23238), 
            .I2(n52506), .I3(\data_in_frame[3][1] ), .O(n52916));
    defparam i2_3_lut_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1654 (.I0(\data_out_frame[9] [5]), .I1(n52951), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [3]), .O(n23410));   // verilog/coms.v(76[16:34])
    defparam i3_4_lut_adj_1654.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(\data_in_frame[2][7] ), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n52473));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1656 (.I0(n23410), .I1(\data_out_frame[10] [0]), 
            .I2(n52975), .I3(GND_net), .O(n53158));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1656.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1657 (.I0(\data_out_frame[12] [1]), .I1(n53158), 
            .I2(n52567), .I3(n52919), .O(n12_adj_5633));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1658 (.I0(\data_out_frame[12] [0]), .I1(n12_adj_5633), 
            .I2(\data_out_frame[14] [2]), .I3(n53128), .O(n52705));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1659 (.I0(n52705), .I1(n4_adj_5562), .I2(GND_net), 
            .I3(GND_net), .O(n52446));
    defparam i2_2_lut_adj_1659.LUT_INIT = 16'h6666;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1660 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53032));
    defparam i1_2_lut_adj_1660.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut_adj_1661 (.I0(\data_out_frame[6] [0]), .I1(n1720), 
            .I2(GND_net), .I3(GND_net), .O(n28_adj_5634));   // verilog/coms.v(75[16:27])
    defparam i5_2_lut_adj_1661.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_1662 (.I0(n24120), .I1(n53113), .I2(n53161), 
            .I3(n52913), .O(n38_adj_5635));   // verilog/coms.v(75[16:27])
    defparam i15_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1663 (.I0(\data_out_frame[14] [6]), .I1(n47414), 
            .I2(n52779), .I3(n1835), .O(n36_adj_5636));   // verilog/coms.v(75[16:27])
    defparam i13_4_lut_adj_1663.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n53032), .I1(n38_adj_5635), .I2(n28_adj_5634), 
            .I3(n52513), .O(n42));   // verilog/coms.v(75[16:27])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1664 (.I0(n1699), .I1(\data_out_frame[14] [3]), 
            .I2(n47527), .I3(n52446), .O(n40));   // verilog/coms.v(75[16:27])
    defparam i17_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1665 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[8][5] ), .I3(n10_adj_5515), .O(n23199));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1666 (.I0(\data_out_frame[5] [5]), .I1(n36_adj_5636), 
            .I2(n52481), .I3(n53122), .O(n41));   // verilog/coms.v(75[16:27])
    defparam i18_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1667 (.I0(n52555), .I1(\data_out_frame[6] [1]), 
            .I2(n52500), .I3(n53036), .O(n39));   // verilog/coms.v(75[16:27])
    defparam i16_4_lut_adj_1667.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n47502));   // verilog/coms.v(75[16:27])
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1668 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[8]_c [3]), .O(n52906));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_4_lut_adj_1669 (.I0(n25699), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n51777));
    defparam i11_4_lut_4_lut_adj_1669.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1670 (.I0(n7_adj_5581), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[19] [1]), .I3(n47502), .O(n53167));
    defparam i4_4_lut_adj_1670.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1671 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52966));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1671.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1672 (.I0(n23958), .I1(n23052), .I2(\data_in_frame[9] [3]), 
            .I3(n52629), .O(n47797));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1672.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1673 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53125));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1673.LUT_INIT = 16'h6666;
    SB_LUT4 i13206_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n26912));
    defparam i13206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1674 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n23812), .I3(\data_in_frame[10][0] ), .O(n47989));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 n62475_bdd_4_lut (.I0(n62475), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n62478));
    defparam n62475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1675 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n23012));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1675.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1676 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52975));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1676.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_950), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n23107));
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1678 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n52452));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1678.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1679 (.I0(n52975), .I1(n23012), .I2(\data_out_frame[8] [1]), 
            .I3(n53125), .O(n10_adj_5637));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1680 (.I0(n52894), .I1(n10_adj_5637), .I2(\data_out_frame[8] [0]), 
            .I3(GND_net), .O(n23437));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1680.LUT_INIT = 16'h9696;
    SB_LUT4 i13203_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n26909));
    defparam i13203_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1681 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n52496));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1681.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1682 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52919));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1682.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1683 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[5] [6]), .I3(n52496), .O(n12_adj_5638));   // verilog/coms.v(77[16:27])
    defparam i5_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1684 (.I0(\data_out_frame[7] [5]), .I1(n12_adj_5638), 
            .I2(n52919), .I3(\data_out_frame[10] [0]), .O(n1510));   // verilog/coms.v(77[16:27])
    defparam i6_4_lut_adj_1684.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1685 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_950), 
            .I2(n23627), .I3(n10_adj_5521), .O(n52629));
    defparam i5_3_lut_4_lut_adj_1685.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1686 (.I0(n23437), .I1(n52452), .I2(\data_out_frame[14] [6]), 
            .I3(GND_net), .O(n24097));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1686.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1687 (.I0(n23149), .I1(n23676), .I2(n52541), 
            .I3(n52948), .O(n52889));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1688 (.I0(n53167), .I1(n53175), .I2(\data_out_frame[16] [4]), 
            .I3(GND_net), .O(n52746));
    defparam i2_3_lut_adj_1688.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1689 (.I0(\data_out_frame[19] [0]), .I1(n52892), 
            .I2(n52822), .I3(n23263), .O(n52721));
    defparam i3_4_lut_adj_1689.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1690 (.I0(n23149), .I1(n23676), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n23670));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1690.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1691 (.I0(n24203), .I1(n52746), .I2(n24097), 
            .I3(\data_out_frame[16] [6]), .O(n23455));
    defparam i3_4_lut_adj_1691.LUT_INIT = 16'h6996;
    SB_LUT4 i13200_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n26906));
    defparam i13200_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1692 (.I0(n23455), .I1(n52721), .I2(\data_out_frame[21] [2]), 
            .I3(GND_net), .O(n48629));
    defparam i2_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1693 (.I0(\data_out_frame[21] [3]), .I1(n53040), 
            .I2(n52746), .I3(n23613), .O(n48494));
    defparam i3_4_lut_adj_1693.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1694 (.I0(n47641), .I1(n52808), .I2(\data_out_frame[23] [6]), 
            .I3(GND_net), .O(n52686));
    defparam i2_3_lut_adj_1694.LUT_INIT = 16'h6969;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[7] [7]), .I1(n52738), .I2(n23318), 
            .I3(\data_in_frame[9] [7]), .O(n20_adj_5510));   // verilog/coms.v(78[16:27])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1695 (.I0(\data_in_frame[7] [7]), .I1(n52738), 
            .I2(\data_in_frame[5] [7]), .I3(n23_adj_5524), .O(n52469));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i13244_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n26950));
    defparam i13244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13241_3_lut_4_lut (.I0(n25699), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n26947));
    defparam i13241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1696 (.I0(n48601), .I1(n52686), .I2(\data_out_frame[25] [6]), 
            .I3(n48494), .O(n12_adj_5639));
    defparam i5_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_208_i3_4_lut (.I0(n48629), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5639), .I3(n8_adj_5561), .O(n3_c));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[25] [6]), 
            .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[25] [5]), 
            .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[25] [4]), 
            .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[24] [6]), 
            .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_3_lut_adj_1702 (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2489 ), 
            .I2(LED_N_3384), .I3(GND_net), .O(n20140));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut_adj_1702.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1703 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n10_adj_9), .I3(n68), .O(n25734));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut_adj_1703.LUT_INIT = 16'h0200;
    SB_LUT4 select_775_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1704 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n161), .I3(n3543), .O(n38306));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1704.LUT_INIT = 16'h2000;
    SB_LUT4 select_775_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1705 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n10_adj_12), .I3(n68), .O(n25750));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut_adj_1705.LUT_INIT = 16'h0200;
    SB_LUT4 select_775_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1706 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n10), .I3(GND_net), .O(n35727));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1706.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1707 (.I0(\data_in_frame[14] [2]), .I1(n48503), 
            .I2(n23518), .I3(GND_net), .O(n22606));
    defparam i1_2_lut_3_lut_adj_1707.LUT_INIT = 16'h6969;
    SB_LUT4 i3_3_lut_4_lut_adj_1708 (.I0(\data_in_frame[14] [2]), .I1(n48503), 
            .I2(n6_adj_5513), .I3(\data_in_frame[16][4] ), .O(n23500));
    defparam i3_3_lut_4_lut_adj_1708.LUT_INIT = 16'h9669;
    SB_LUT4 select_775_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[23] [5]), 
            .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[23] [3]), 
            .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'ha088;
    SB_LUT4 i13073_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[6][7] ), .O(n26779));
    defparam i13073_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44831_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59291));   // verilog/coms.v(158[12:15])
    defparam i44831_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13070_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[6][6] ), .O(n26776));
    defparam i13070_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13058_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[6][3] ), .O(n26764));
    defparam i13058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1711 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n23676));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1711.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13055_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[6][2] ), .O(n26761));
    defparam i13055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_775_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13052_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[6][1] ), .O(n26758));
    defparam i13052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_3_lut_4_lut (.I0(n25721), .I1(reset), .I2(\data_in_frame[6] [0]), 
            .I3(rx_data[0]), .O(n51805));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 select_775_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(\data_in_frame[13] [1]), .I1(n54985), 
            .I2(n53058), .I3(GND_net), .O(n6_adj_5406));
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[21] [3]), 
            .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'ha088;
    SB_LUT4 i1_3_lut_4_lut_adj_1714 (.I0(\FRAME_MATCHER.i_31__N_2484 ), .I1(\FRAME_MATCHER.i_31__N_2488 ), 
            .I2(n52403), .I3(LED_c), .O(n24628));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1714.LUT_INIT = 16'hfe00;
    SB_LUT4 select_775_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1715 (.I0(\data_in_frame[13] [1]), .I1(n54985), 
            .I2(\data_in_frame[16] [0]), .I3(GND_net), .O(n52678));
    defparam i1_2_lut_3_lut_adj_1715.LUT_INIT = 16'h6969;
    SB_LUT4 i19877_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13]_c [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27060));
    defparam i19877_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_775_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_3_lut_4_lut_adj_1716 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[15] [2]), .I3(n16_c), .O(n18));   // verilog/coms.v(73[16:27])
    defparam i8_3_lut_4_lut_adj_1716.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1717 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n53164), .I3(n54639), .O(n52791));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1717.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1718 (.I0(n54113), .I1(n47424), .I2(\data_in_frame[21] [6]), 
            .I3(\data_in_frame[21] [7]), .O(n6_adj_5543));
    defparam i1_3_lut_4_lut_adj_1718.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1719 (.I0(n54113), .I1(n47424), .I2(n54169), 
            .I3(GND_net), .O(n48458));
    defparam i1_2_lut_3_lut_adj_1719.LUT_INIT = 16'h9696;
    SB_LUT4 select_775_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_150_i2_4_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_150_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[18] [5]), 
            .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'ha088;
    SB_LUT4 i24712_2_lut_3_lut (.I0(n3543), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n38302));
    defparam i24712_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_775_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i46287_3_lut (.I0(n62688), .I1(n62430), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n61187));
    defparam i46287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44830_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59290));   // verilog/coms.v(158[12:15])
    defparam i44830_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45329_2_lut (.I0(n62622), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n59383));
    defparam i45329_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1721 (.I0(\FRAME_MATCHER.i_31__N_2484 ), .I1(\FRAME_MATCHER.i_31__N_2488 ), 
            .I2(\FRAME_MATCHER.i_31__N_2490 ), .I3(GND_net), .O(n3543));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1721.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[18] [0]), 
            .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_317_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10));   // verilog/coms.v(157[7:23])
    defparam equal_317_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_309_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_12));   // verilog/coms.v(157[7:23])
    defparam equal_309_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 select_775_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13259_3_lut (.I0(\data_in_frame[13]_c [3]), .I1(rx_data[3]), 
            .I2(n52427), .I3(GND_net), .O(n26965));   // verilog/coms.v(130[12] 305[6])
    defparam i13259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[6] [6]), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5269));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44829_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59289));   // verilog/coms.v(158[12:15])
    defparam i44829_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47560 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n62457));
    defparam byte_transmit_counter_0__bdd_4_lut_47560.LUT_INIT = 16'he4aa;
    SB_LUT4 n62457_bdd_4_lut (.I0(n62457), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n62460));
    defparam n62457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47551 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56822), .I2(n56823), .I3(\byte_transmit_counter[2] ), 
            .O(n62451));
    defparam byte_transmit_counter_1__bdd_4_lut_47551.LUT_INIT = 16'he4aa;
    SB_LUT4 select_775_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n62451_bdd_4_lut (.I0(n62451), .I1(n56604), .I2(n56603), .I3(\byte_transmit_counter[2] ), 
            .O(n62454));
    defparam n62451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_775_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21271_3_lut_4_lut (.I0(\Kp[14] ), .I1(\data_in_frame[2]_c [6]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27027));
    defparam i21271_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_775_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5268));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_47595 (.I0(\byte_transmit_counter[3] ), 
            .I1(n61175), .I2(n59368), .I3(\byte_transmit_counter[4] ), 
            .O(n62445));
    defparam byte_transmit_counter_3__bdd_4_lut_47595.LUT_INIT = 16'he4aa;
    SB_LUT4 n62445_bdd_4_lut (.I0(n62445), .I1(n14_adj_5582), .I2(n7_adj_5580), 
            .I3(\byte_transmit_counter[4] ), .O(tx_data[5]));
    defparam n62445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i44828_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59288));   // verilog/coms.v(158[12:15])
    defparam i44828_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44827_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59287));   // verilog/coms.v(158[12:15])
    defparam i44827_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[6] [4]), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5267));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'ha088;
    SB_LUT4 i44824_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59286));   // verilog/coms.v(158[12:15])
    defparam i44824_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5266));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44822_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59284));   // verilog/coms.v(158[12:15])
    defparam i44822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44819_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59283));   // verilog/coms.v(158[12:15])
    defparam i44819_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5265));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1725 (.I0(n5_adj_5534), .I1(n3303), .I2(n22848), 
            .I3(\FRAME_MATCHER.i_31__N_2488 ), .O(n54683));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1725.LUT_INIT = 16'hfbfa;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(\FRAME_MATCHER.i_31__N_2490 ), .I1(n2056), 
            .I2(n2125), .I3(n54683), .O(n24602));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hb3a0;
    SB_LUT4 i463_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2488 ), .I2(GND_net), 
            .I3(GND_net), .O(n2165));   // verilog/coms.v(148[4] 304[11])
    defparam i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20444_3_lut_4_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10]_c [5]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27610));
    defparam i20444_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(\FRAME_MATCHER.i_31__N_2488 ), .I1(n2059), 
            .I2(n2113), .I3(n54637), .O(n51443));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'hb3a0;
    SB_LUT4 select_775_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5264));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5029_4_lut (.I0(n2060), .I1(\FRAME_MATCHER.state[3] ), .I2(n2062), 
            .I3(n22848), .O(n18397));   // verilog/coms.v(148[4] 304[11])
    defparam i5029_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i452_2_lut (.I0(\FRAME_MATCHER.state_31__N_2588 [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(GND_net), .I3(GND_net), .O(n2154));   // verilog/coms.v(148[4] 304[11])
    defparam i452_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i451_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2484 ), .I2(GND_net), 
            .I3(GND_net), .O(n2153));   // verilog/coms.v(148[4] 304[11])
    defparam i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24456_4_lut (.I0(n8_adj_5554), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22768), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i24456_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1728 (.I0(\FRAME_MATCHER.i [4]), .I1(n22929), .I2(GND_net), 
            .I3(GND_net), .O(n22768));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1728.LUT_INIT = 16'heeee;
    SB_LUT4 i24451_4_lut (.I0(n5_adj_5522), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i24451_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i2_2_lut_adj_1729 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2484 ), 
            .I2(GND_net), .I3(GND_net), .O(n20118));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1729.LUT_INIT = 16'h4444;
    SB_LUT4 i3_2_lut (.I0(n22848), .I1(\FRAME_MATCHER.i_31__N_2483 ), .I2(GND_net), 
            .I3(GND_net), .O(n24375));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n2060), .I1(n2110), .I2(n24375), .I3(\FRAME_MATCHER.i_31__N_2488 ), 
            .O(n4_adj_5641));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'heca0;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n2062), .I1(n2122), .I2(n4_adj_5641), 
            .I3(\FRAME_MATCHER.i_31__N_2490 ), .O(n24379));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'h5450;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n2059), .I1(n24379), .I2(n2056), .I3(n20118), 
            .O(n24380));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'heccc;
    SB_LUT4 i44816_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59282));   // verilog/coms.v(158[12:15])
    defparam i44816_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_47541 (.I0(\byte_transmit_counter[1] ), 
            .I1(n56582), .I2(n56583), .I3(\byte_transmit_counter[2] ), 
            .O(n62439));
    defparam byte_transmit_counter_1__bdd_4_lut_47541.LUT_INIT = 16'he4aa;
    SB_LUT4 i44813_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59281));   // verilog/coms.v(158[12:15])
    defparam i44813_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44511_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59280));   // verilog/coms.v(158[12:15])
    defparam i44511_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_adj_1733 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5642));
    defparam i2_2_lut_adj_1733.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1734 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5643));
    defparam i6_4_lut_adj_1734.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1735 (.I0(\data_in[3] [6]), .I1(n14_adj_5643), 
            .I2(n10_adj_5642), .I3(\data_in[2] [1]), .O(n22932));
    defparam i7_4_lut_adj_1735.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1736 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n22932), .I3(\data_in[0] [1]), .O(n20_adj_5644));
    defparam i8_4_lut_adj_1736.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1737 (.I0(n22787), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5645));
    defparam i7_4_lut_adj_1737.LUT_INIT = 16'hfeff;
    SB_LUT4 i41580_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [5]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n56471));
    defparam i41580_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n56471), .I1(n19_adj_5645), .I2(n20_adj_5644), 
            .I3(GND_net), .O(n2056));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1738 (.I0(\data_in[2] [4]), .I1(n22932), .I2(\data_in[1] [5]), 
            .I3(n22884), .O(n18_adj_5646));
    defparam i7_4_lut_adj_1738.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1739 (.I0(\data_in[0] [6]), .I1(n18_adj_5646), 
            .I2(\data_in[3] [0]), .I3(n22867), .O(n20_adj_5647));
    defparam i9_4_lut_adj_1739.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5648));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1740 (.I0(n15_adj_5648), .I1(n20_adj_5647), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n2059));
    defparam i10_4_lut_adj_1740.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1741 (.I0(Kp_23__N_1724), .I1(\FRAME_MATCHER.i_31__N_2489 ), 
            .I2(GND_net), .I3(GND_net), .O(n30909));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1741.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1742 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5649));
    defparam i6_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1743 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_5650));
    defparam i7_4_lut_adj_1743.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1744 (.I0(n17_adj_5650), .I1(\data_in[1] [6]), 
            .I2(n16_adj_5649), .I3(\data_in[3] [7]), .O(n22867));
    defparam i9_4_lut_adj_1744.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1745 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5651));
    defparam i4_4_lut_adj_1745.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1746 (.I0(\data_in[3] [4]), .I1(n10_adj_5651), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n22884));
    defparam i5_3_lut_adj_1746.LUT_INIT = 16'hdfdf;
    SB_LUT4 i5_3_lut_adj_1747 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5652));
    defparam i5_3_lut_adj_1747.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1748 (.I0(\data_in[0] [6]), .I1(n22884), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5653));
    defparam i6_4_lut_adj_1748.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1749 (.I0(n15_adj_5653), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5652), .I3(\data_in[0] [3]), .O(n22787));
    defparam i8_4_lut_adj_1749.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1750 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n22787), .O(n16_adj_5654));
    defparam i6_4_lut_adj_1750.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1751 (.I0(n22867), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5655));
    defparam i7_4_lut_adj_1751.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1752 (.I0(n17_adj_5655), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5654), .I3(\data_in[3] [3]), .O(n2062));
    defparam i9_4_lut_adj_1752.LUT_INIT = 16'hfbff;
    SB_LUT4 i369_2_lut (.I0(n2059), .I1(n2056), .I2(GND_net), .I3(GND_net), 
            .O(n2060));   // verilog/coms.v(142[4] 144[7])
    defparam i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1753 (.I0(n38421), .I1(n54168), .I2(\FRAME_MATCHER.i_31__N_2487 ), 
            .I3(n37879), .O(n6_adj_5656));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1753.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1754 (.I0(n30909), .I1(n6_adj_5656), .I2(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2485 ), .O(n62844));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1754.LUT_INIT = 16'hefee;
    SB_LUT4 n62439_bdd_4_lut (.I0(n62439), .I1(n56844), .I2(n56843), .I3(\byte_transmit_counter[2] ), 
            .O(n62442));
    defparam n62439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11678_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3543), 
            .I3(\FRAME_MATCHER.i_31__N_2483 ), .O(n25384));   // verilog/coms.v(158[12:15])
    defparam i11678_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47546 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n62433));
    defparam byte_transmit_counter_0__bdd_4_lut_47546.LUT_INIT = 16'he4aa;
    SB_LUT4 n62433_bdd_4_lut (.I0(n62433), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n62436));
    defparam n62433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i44664_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59189));   // verilog/coms.v(158[12:15])
    defparam i44664_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44663_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59188));   // verilog/coms.v(158[12:15])
    defparam i44663_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n62697));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n62691_bdd_4_lut (.I0(n62691), .I1(n62496), .I2(n7_adj_5579), 
            .I3(\byte_transmit_counter[4] ), .O(tx_data[0]));
    defparam n62691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[6] [0]), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5263));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_47514 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n62409));
    defparam byte_transmit_counter_0__bdd_4_lut_47514.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1756 (.I0(reset), .I1(n38302), .I2(n10_adj_9), 
            .I3(GND_net), .O(n52430));
    defparam i1_2_lut_3_lut_adj_1756.LUT_INIT = 16'hfbfb;
    SB_LUT4 n62697_bdd_4_lut (.I0(n62697), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n62700));
    defparam n62697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(\byte_transmit_counter[3] ), 
            .I1(n61049), .I2(n59358), .I3(\byte_transmit_counter[4] ), 
            .O(n62691));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1757 (.I0(reset), .I1(n38302), .I2(n10), 
            .I3(GND_net), .O(n52434));
    defparam i1_2_lut_3_lut_adj_1757.LUT_INIT = 16'hfbfb;
    SB_LUT4 select_775_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5262));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i20770_3_lut_4_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8]_c [3]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27596));
    defparam i20770_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_775_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[14] [7]), 
            .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[14] [6]), 
            .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[14] [4]), 
            .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n62409_bdd_4_lut (.I0(n62409), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n62412));
    defparam n62409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_775_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[13] [5]), 
            .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1762 (.I0(reset), .I1(n38302), .I2(n10_adj_12), 
            .I3(GND_net), .O(n52424));
    defparam i1_2_lut_3_lut_adj_1762.LUT_INIT = 16'hfbfb;
    SB_LUT4 select_775_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[5] [7]), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5261));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5306));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i44662_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59187));   // verilog/coms.v(158[12:15])
    defparam i44662_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_775_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2485 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2487 ), 
            .I2(GND_net), .I3(GND_net), .O(n52326));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21410_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n20140), .I3(GND_net), .O(n26917));
    defparam i21410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13101_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n26807));
    defparam i13101_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13098_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n26804));
    defparam i13098_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i422_4_lut_4_lut (.I0(n2059), .I1(n2062), .I2(n2056), .I3(n3303), 
            .O(n2113));   // verilog/coms.v(139[4] 141[7])
    defparam i422_4_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_4_lut_adj_1764 (.I0(\data_out_frame[19] [4]), .I1(n24097), 
            .I2(n52523), .I3(n48452), .O(n52808));
    defparam i1_2_lut_4_lut_adj_1764.LUT_INIT = 16'h6996;
    SB_LUT4 select_775_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1765 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .I2(\data_out_frame[0][2] ), .I3(GND_net), .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1765.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13095_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n26801));
    defparam i13095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13092_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n26798));
    defparam i13092_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13088_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n26794));
    defparam i13088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5260));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13085_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n26791));
    defparam i13085_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(\FRAME_MATCHER.i_31__N_2485 ), .I1(\data_out_frame[5] [5]), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'ha088;
    SB_LUT4 select_775_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_775_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5296));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5295));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i47426_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3521[0]), 
            .I2(n38421), .I3(GND_net), .O(tx_transmit_N_3392));
    defparam i47426_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 select_775_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5294));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_775_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(\FRAME_MATCHER.state_31__N_2588 [3]), .I3(GND_net), .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13082_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n26788));
    defparam i13082_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_775_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2485 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2588 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_775_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13077_3_lut_4_lut (.I0(n37), .I1(n52434), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n26783));
    defparam i13077_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1044_i24_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n4757[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1044_i24_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i44651_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2483 ), 
            .I2(GND_net), .I3(GND_net), .O(n59183));   // verilog/coms.v(158[12:15])
    defparam i44651_2_lut.LUT_INIT = 16'h2222;
    uart_tx tx (.n62840(n62840), .r_SM_Main({r_SM_Main}), .clk16MHz(clk16MHz), 
            .\r_SM_Main_2__N_3512[1] (r_SM_Main_2__N_3512[1]), .GND_net(GND_net), 
            .r_Clock_Count({r_Clock_Count}), .tx_o(tx_o), .tx_data({tx_data[7:3], 
            \tx_data[2] , tx_data[1:0]}), .VCC_net(VCC_net), .n26943(n26943), 
            .tx_active(tx_active), .n23(n23), .\o_Rx_DV_N_3464[12] (\o_Rx_DV_N_3464[12] ), 
            .n4858(n4858), .\o_Rx_DV_N_3464[24] (\o_Rx_DV_N_3464[24] ), 
            .n27(n27), .n29(n29), .\r_SM_Main_2__N_3521[0] (r_SM_Main_2__N_3521[0]), 
            .n53934(n53934), .n6(n6_adj_13), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .n27247(n27247), .rx_data({rx_data}), 
            .clk16MHz(clk16MHz), .baudrate({baudrate}), .\o_Rx_DV_N_3464[24] (\o_Rx_DV_N_3464[24] ), 
            .n29(n29), .n23(n23), .n55830(n55830), .VCC_net(VCC_net), 
            .n27246(n27246), .n27245(n27245), .n27243(n27243), .n27242(n27242), 
            .\o_Rx_DV_N_3464[8] (\o_Rx_DV_N_3464[8] ), .\o_Rx_DV_N_3464[12] (\o_Rx_DV_N_3464[12] ), 
            .n4855(n4855), .n52352(n52352), .r_SM_Main({Open_27, \r_SM_Main[1]_adj_14 , 
            Open_28}), .n27(n27), .n25039(n25039), .n27241(n27241), 
            .n27240(n27240), .\r_SM_Main[2] (\r_SM_Main[2]_adj_15 ), .n55782(n55782), 
            .r_Clock_Count({r_Clock_Count_adj_24}), .n55798(n55798), .n55750(n55750), 
            .n55766(n55766), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .n22878(n22878), 
            .\o_Rx_DV_N_3464[7] (\o_Rx_DV_N_3464[7] ), .\o_Rx_DV_N_3464[6] (\o_Rx_DV_N_3464[6] ), 
            .\o_Rx_DV_N_3464[5] (\o_Rx_DV_N_3464[5] ), .\o_Rx_DV_N_3464[4] (\o_Rx_DV_N_3464[4] ), 
            .\o_Rx_DV_N_3464[3] (\o_Rx_DV_N_3464[3] ), .\o_Rx_DV_N_3464[2] (\o_Rx_DV_N_3464[2] ), 
            .\o_Rx_DV_N_3464[1] (\o_Rx_DV_N_3464[1] ), .\o_Rx_DV_N_3464[0] (\o_Rx_DV_N_3464[0] ), 
            .n25264(n25264), .n27583(n27583), .n48661(n48661), .rx_data_ready(rx_data_ready), 
            .n27579(n27579), .r_Bit_Index({Open_29, Open_30, \r_Bit_Index[0] }), 
            .n53350(n53350), .n55734(n55734), .n55846(n55846), .n55814(n55814), 
            .n4858(n4858), .\r_SM_Main_2__N_3512[1] (r_SM_Main_2__N_3512[1]), 
            .\r_SM_Main[0]_adj_7 (r_SM_Main[0]), .n53934(n53934)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n62840, r_SM_Main, clk16MHz, \r_SM_Main_2__N_3512[1] , 
            GND_net, r_Clock_Count, tx_o, tx_data, VCC_net, n26943, 
            tx_active, n23, \o_Rx_DV_N_3464[12] , n4858, \o_Rx_DV_N_3464[24] , 
            n27, n29, \r_SM_Main_2__N_3521[0] , n53934, n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input n62840;
    output [2:0]r_SM_Main;
    input clk16MHz;
    input \r_SM_Main_2__N_3512[1] ;
    input GND_net;
    output [8:0]r_Clock_Count;
    output tx_o;
    input [7:0]tx_data;
    input VCC_net;
    input n26943;
    output tx_active;
    input n23;
    input \o_Rx_DV_N_3464[12] ;
    input n4858;
    input \o_Rx_DV_N_3464[24] ;
    input n27;
    input n29;
    input \r_SM_Main_2__N_3521[0] ;
    input n53934;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n53907, n59203, n53390;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n48691;
    wire [8:0]n41;
    
    wire n1, n35561, n3, n20187;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n48693, n46257, n46256;
    wire [2:0]n460;
    
    wire n53939, n52322, n46255, n46254, n46253, n3_adj_5252, n46252, 
        n46251, n62535, n62538, n46250, n32, n55456, n6_c, n9, 
        n53304, n62424, n5, n55564, n55570, n62421;
    
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n62840));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i38343_rep_31_2_lut (.I0(\r_SM_Main_2__N_3512[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n53907));
    defparam i38343_rep_31_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut (.I0(n59203), .I1(n53390), .I2(r_Bit_Index[0]), 
            .I3(n53907), .O(n48691));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_DFFESR r_Clock_Count_1945__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n48693), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n48691));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_1945_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n46257), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1945__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_LUT4 r_Clock_Count_1945_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n46256), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1945__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1945__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n35561));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n53390), 
            .D(n460[1]), .R(n53939));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n53390), 
            .D(n460[2]), .R(n52322));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n26943));   // verilog/uart_tx.v(41[10] 144[8])
    SB_CARRY r_Clock_Count_1945_add_4_9 (.CI(n46256), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n46257));
    SB_LUT4 r_Clock_Count_1945_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n46255), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_8 (.CI(n46255), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n46256));
    SB_LUT4 r_Clock_Count_1945_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n46254), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_7 (.CI(n46254), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n46255));
    SB_LUT4 r_Clock_Count_1945_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n46253), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5252), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n20187), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_CARRY r_Clock_Count_1945_add_4_6 (.CI(n46253), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n46254));
    SB_LUT4 r_Clock_Count_1945_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n46252), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_5 (.CI(n46252), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n46253));
    SB_LUT4 r_Clock_Count_1945_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n46251), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_4 (.CI(n46251), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n46252));
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[3]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n62535));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n62535_bdd_4_lut (.I0(n62535), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[1]), 
            .I3(r_Bit_Index[1]), .O(n62538));
    defparam n62535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Clock_Count_1945_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n46250), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_3 (.CI(n46250), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n46251));
    SB_LUT4 r_Clock_Count_1945_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1945_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1945_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n46250));
    SB_LUT4 i1_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n32));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut (.I0(n23), .I1(\o_Rx_DV_N_3464[12] ), .I2(n4858), 
            .I3(n32), .O(n55456));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1125 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n27), .I2(n29), 
            .I3(n55456), .O(n6_c));
    defparam i1_4_lut_adj_1125.LUT_INIT = 16'h0100;
    SB_LUT4 i23_3_lut (.I0(\r_SM_Main_2__N_3521[0] ), .I1(n6_c), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3512[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n48693));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38455_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53304));
    defparam i38455_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24907107_i1_3_lut (.I0(n62424), .I1(n62538), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n5));
    defparam i24907107_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n5), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i2_3_lut_4_lut (.I0(\r_SM_Main_2__N_3521[0] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n20187));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut (.I0(n4858), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n55564));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1126 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3464[12] ), 
            .I3(n55564), .O(n55570));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'h0100;
    SB_LUT4 i6511_4_lut (.I0(\o_Rx_DV_N_3464[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n55570), .O(n3_adj_5252));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i6511_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut_47610 (.I0(r_Bit_Index[2]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[6]), .I3(r_Bit_Index[1]), .O(n62421));
    defparam r_Bit_Index_2__bdd_4_lut_47610.LUT_INIT = 16'he4aa;
    SB_LUT4 n62421_bdd_4_lut (.I0(n62421), .I1(r_Tx_Data[4]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n62424));
    defparam n62421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i47432_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(\r_SM_Main_2__N_3512[1] ), 
            .I3(r_SM_Main[0]), .O(n35561));
    defparam i47432_4_lut.LUT_INIT = 16'h0515;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n53934), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3521[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1127 (.I0(n6_c), .I1(n53304), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n52322));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_3_lut_adj_1127.LUT_INIT = 16'h2323;
    SB_LUT4 i21959_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i21959_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut_adj_1128 (.I0(r_SM_Main[1]), .I1(n53907), .I2(n53304), 
            .I3(n32), .O(n53939));
    defparam i1_4_lut_adj_1128.LUT_INIT = 16'h0301;
    SB_LUT4 i11_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45371_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n59203));   // verilog/uart_tx.v(32[16:25])
    defparam i45371_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i47324_2_lut_4_lut (.I0(\r_SM_Main_2__N_3512[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n53390));
    defparam i47324_2_lut_4_lut.LUT_INIT = 16'h0007;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, n27247, rx_data, clk16MHz, baudrate, \o_Rx_DV_N_3464[24] , 
            n29, n23, n55830, VCC_net, n27246, n27245, n27243, 
            n27242, \o_Rx_DV_N_3464[8] , \o_Rx_DV_N_3464[12] , n4855, 
            n52352, r_SM_Main, n27, n25039, n27241, n27240, \r_SM_Main[2] , 
            n55782, r_Clock_Count, n55798, n55750, n55766, r_Rx_Data, 
            RX_N_2, n22878, \o_Rx_DV_N_3464[7] , \o_Rx_DV_N_3464[6] , 
            \o_Rx_DV_N_3464[5] , \o_Rx_DV_N_3464[4] , \o_Rx_DV_N_3464[3] , 
            \o_Rx_DV_N_3464[2] , \o_Rx_DV_N_3464[1] , \o_Rx_DV_N_3464[0] , 
            n25264, n27583, n48661, rx_data_ready, n27579, r_Bit_Index, 
            n53350, n55734, n55846, n55814, n4858, \r_SM_Main_2__N_3512[1] , 
            \r_SM_Main[0]_adj_7 , n53934) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n27247;
    output [7:0]rx_data;
    input clk16MHz;
    input [31:0]baudrate;
    output \o_Rx_DV_N_3464[24] ;
    output n29;
    output n23;
    output n55830;
    input VCC_net;
    input n27246;
    input n27245;
    input n27243;
    input n27242;
    output \o_Rx_DV_N_3464[8] ;
    output \o_Rx_DV_N_3464[12] ;
    input n4855;
    input n52352;
    output [2:0]r_SM_Main;
    output n27;
    output n25039;
    input n27241;
    input n27240;
    output \r_SM_Main[2] ;
    output n55782;
    output [7:0]r_Clock_Count;
    output n55798;
    output n55750;
    output n55766;
    output r_Rx_Data;
    input RX_N_2;
    output n22878;
    output \o_Rx_DV_N_3464[7] ;
    output \o_Rx_DV_N_3464[6] ;
    output \o_Rx_DV_N_3464[5] ;
    output \o_Rx_DV_N_3464[4] ;
    output \o_Rx_DV_N_3464[3] ;
    output \o_Rx_DV_N_3464[2] ;
    output \o_Rx_DV_N_3464[1] ;
    output \o_Rx_DV_N_3464[0] ;
    output n25264;
    input n27583;
    input n48661;
    output rx_data_ready;
    input n27579;
    output [2:0]r_Bit_Index;
    output n53350;
    output n55734;
    output n55846;
    output n55814;
    input n4858;
    output \r_SM_Main_2__N_3512[1] ;
    input \r_SM_Main[0]_adj_7 ;
    output n53934;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n7589;
    
    wire n1411, n1460, n45839;
    wire [23:0]n7953;
    
    wire n3171, n698, n46038, n45840, n46039, n1412, n1011, n45838, 
        n3172, n858, n46037, n1413, n856, n45837, n61424, n37, 
        n60660, n55376, n538, n46036, n53438, n55824, n1414, n45836;
    wire [23:0]n7927;
    
    wire n3046, n3082, n46035, n3047, n3188, n46034, n3048, n3084, 
        n46033, n1415, n45835, n3049, n2977, n46032, n56481, n56148, 
        n56479, n56102, n56537, n53446, n14, n25, n22, n56162, 
        n55316, n55314, n56152, n22959, n59276, n53458, n59273;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(37[17:26])
    
    wire n3154;
    wire [23:0]n294;
    
    wire n41, n3155, n39, n55770, n55776, n3158, n33, n3157, 
        n35, n3156, n37_adj_4979, n3160, n29_adj_4980, n3159, n31, 
        n3163, n23_adj_4981, n62842, n12, n59813, n61919, n3162, 
        n25_adj_4982, n7, n3152, n45, n3153, n43, n3170, n9, 
        n3166, n17, n3165, n19, n3164, n21, n3169, n11, n3168, 
        n13, n3167, n15, n3161, n27_adj_4983, n59582, n59594, 
        n16, n55354, n48;
    wire [7:0]n1;
    
    wire n25247, n26549, n6, n59536, n8, n24, n27_adj_4985, n61920, 
        n3274, n59606, n60448, n55786, n55792, n60444, n55356, 
        n53488, n61743, n61133, n61947, n12_adj_4986, n56533, n53496, 
        n48_adj_4987, n4, n61641, n3050, n2867, n46031, n55738, 
        n55744, n61642, n59570, n10, n30, n59574, n61994, n61560, 
        n62138, n3051, n2754, n46030, n62139, n6_adj_4988, n61643, 
        n61644, n22971, n53442, n59540, n61225, n61558, n62113, 
        n59546, n2831, n39_adj_4989, n2832, n37_adj_4990, n61817, 
        n40, n2829, n43_adj_4991, n2830, n41_adj_4992, n2835, n31_adj_4993, 
        n2834, n33_adj_4994, n2838, n25_adj_4995, n2837, n27_adj_4996, 
        n2836, n29_adj_4997, n55328, n3151, n3253, n3052, n2638, 
        n46029, n3053, n2519, n46028, n61819, n56260, n56108, 
        n56104, n55336, n2841, n19_adj_4998;
    wire [23:0]n7563;
    
    wire n1261, n1602, n45834, n2840, n21_adj_4999, n1262, n1459, 
        n45833, n2839, n23_adj_5000, n1263, n45832, n2833, n35_adj_5001, 
        n54288, n1264, n45831, n2843, n15_adj_5002, n2842, n17_adj_5003, 
        n59871, n2844, n60801, n61281, n3054, n2397, n46027, n61273, 
        n59878, n55754, n55760, n2845, n12_adj_5004, n3055, n2272, 
        n46026, n61427, n1265, n45830, n20, n38, n61428, n3, 
        n3056, n2144, n46025, r_Rx_Data_R, n59859, n1266, n45829, 
        n33_adj_5005, n18, n59853, n61857, n2939;
    wire [23:0]n7901;
    
    wire n60654, n3057, n2013, n46024, n2940, n16_adj_5006, n24_adj_5007, 
        n14_adj_5008, n59896, n61903, n61904, n31_adj_5009, n37_adj_5010, 
        n35_adj_5011, n3058, n1879, n46023, n61736, n61611, n25_adj_5012, 
        n1267, n45828, n62118, n60652, n3059, n1742, n46022, n62144, 
        n2941, n2828, n62145, n27_adj_5013, n2957, n3065, n21_adj_5014, 
        n3060, n46021, n2716, n41_adj_5015, n3061, n46020, n23_adj_5016, 
        n2714, n45_adj_5017, n2717, n39_adj_5018, n2715, n43_adj_5019, 
        n2720, n33_adj_5020, n9_adj_5021, n2719, n35_adj_5022, n2723, 
        n27_adj_5023, n53492, n2722, n29_adj_5024, n2721, n31_adj_5025, 
        n2728, n17_adj_5026, n2727, n19_adj_5027, n2726, n21_adj_5028, 
        n2725, n23_adj_5029, n3062, n46019, n2724, n25_adj_5030, 
        n2718, n37_adj_5031, n59948, n2729, n60847, n61309, n3064, 
        n61305, n11_adj_5032, n3063, n46018, n59950;
    wire [23:0]n7537;
    
    wire n1111, n45827, n19_adj_5033, n2730, n14_adj_5034, n61433, 
        n61434, n1112, n45826, n46017, n1113, n45825, n46016, 
        n1114, n45824, n22_adj_5035, n40_adj_5036, n3066, n46015, 
        n59938, n13_adj_5037, n15_adj_5038, n20_adj_5039, n59934, 
        n61535, n60648, n55374, n17_adj_5040, n18_adj_5041, n26, 
        n16_adj_5042, n59960, n61901, n61902, n61740, n61625, n29_adj_5043, 
        n59633, n61973, n60558, n60646, n61975, n61179, n61177, 
        n59639;
    wire [23:0]n7875;
    
    wire n2956, n6_adj_5044, n61649, n2601, n37_adj_5045, n2938, 
        n46014, n1115, n45823, n46013, n46012, n1116, n45822, 
        n46011, n14_adj_5046, n32, n2942, n46010, n55352, n2943, 
        n46009, n2944, n46008, n61650, n2945, n46007, n2598, n43_adj_5047, 
        n2946, n46006, n2599, n41_adj_5048, n59628, n12_adj_5049, 
        n59625, n61990, n2600, n39_adj_5050, n61550, n2947, n46005, 
        n2948, n46004, n2604, n31_adj_5051, n8_adj_5052, n61651, 
        n61652, n2603, n33_adj_5053, n2949, n46003, n2602, n35_adj_5054, 
        n59661, n60540, n10_adj_5055, n61223, n61548, n2950, n46002, 
        n61472, n62136, n2951, n46001, n2606, n27_adj_5056, n2952, 
        n46000, n61645, n62152, n2605, n29_adj_5057, n2610, n19_adj_5058, 
        n2609, n21_adj_5059, n62153, n62143, n2608, n23_adj_5060, 
        n2607, n25_adj_5061, n61911, n2611, n17_adj_5062, n2953, 
        n45999, n61912, n60014, n2954, n45998, n60010, n61635, 
        n2612, n16_adj_5063, n2955, n45997, n61439, n45996, n61440, 
        n60012, n60861, n22_adj_5064, n61533, n60636, n20_adj_5065, 
        n28, n45995, n18_adj_5066, n60008, n61899, n61900, n61746, 
        n60867, n61741, n55372, n60634, n62016, n2827, n45994, 
        n2597, n62017, n45993, n45992;
    wire [23:0]n7849;
    
    wire n45991, n45990, n45989, n2480, n39_adj_5067, n2477, n45_adj_5068, 
        n45988, n2479, n41_adj_5069, n2478, n43_adj_5070, n2485, 
        n29_adj_5071, n2484, n31_adj_5072, n2483, n33_adj_5073, n2482, 
        n35_adj_5074, n2481, n37_adj_5075, n2489, n21_adj_5076, n2488, 
        n23_adj_5077, n45987, n45986, n2487, n25_adj_5078, n2486, 
        n27_adj_5079, n2490, n19_adj_5080, n60063, n60055, n45985, 
        n45671, n45670, n55340, n45984, n56571, n45669, n55416, 
        n61669, n2491, n18_adj_5081, n45668;
    wire [24:0]o_Rx_DV_N_3464;
    
    wire n45667, n55414, n43_adj_5082, n45983, n61445, n45982, n61446, 
        n45666, n55412, n45665, n45981, n60057, n60887, n45664, 
        n55410, n45663, n55408, n45980, n24_adj_5083, n26_adj_5084, 
        n60630, n45979, n45978, n45662, n55338, n45661, n55406, 
        n45660, n45977, n45659, n45658, n45657, n45976, n55370, 
        n53450, n45656, n2713, n45975, n45974, n45655, n22_adj_5085, 
        n30_adj_5086, n20_adj_5087, n60045, n61897, n61898, n45654, 
        n45973, n61748, n60893, n45653, n45652, n45972, n45651, 
        n45971, n61530, n60628, n45650, n45970, n45649, n45969, 
        n45648, n22965, n61532;
    wire [23:0]n7823;
    
    wire n45968, n45967, n29_adj_5088, n61732, n39_adj_5089, n35_adj_5090, 
        n59790, n61577, n38_adj_5091, n2356, n41_adj_5092, n40_adj_5093, 
        n42, n2357, n39_adj_5094, n2358, n37_adj_5095, n2359, n35_adj_5096, 
        n59521, n61683, n2362, n29_adj_5097, n2361, n31_adj_5098, 
        n2360, n33_adj_5099, n61684, n2365, n23_adj_5100, n2364, 
        n25_adj_5101, n2363, n27_adj_5102, n2366, n21_adj_5103, n60134, 
        n60123, n2367, n20_adj_5104, n26_adj_5105, n28_adj_5106, n24_adj_5107, 
        n32_adj_5108, n22_adj_5109, n60121, n61891, n61892, n61752, 
        n61701, n60129, n61986, n60624, n62056, n2355, n62057, 
        n2354, n62029;
    wire [23:0]n7797;
    
    wire n2229, n43_adj_5110, n2231, n39_adj_5111, n2230, n41_adj_5112, 
        n2232, n37_adj_5113, n2235, n31_adj_5114, n2234, n33_adj_5115, 
        n2233, n35_adj_5116, n2238, n25_adj_5117, n2237, n27_adj_5118, 
        n45966, n45965, n2236, n29_adj_5119, n16_adj_5120, n2239, 
        n23_adj_5121, n60208, n45964, n60180, n45963, n61921, n41_adj_5122, 
        n59781, n62090, n31_adj_5123, n60658, n2240, n22_adj_5124, 
        n62156, n62157, n28_adj_5125, n30_adj_5126, n45962, n45961, 
        n62149, n45960, n45959, n1556, n45958, n26_adj_5127, n34, 
        n24_adj_5128, n60178, n61889, n61890, n61754, n61711, n60194, 
        n61663, n60620, n55368, n53454, n56150, n61861, n2228, 
        n61862, n2596, n45957;
    wire [2:0]r_SM_Main_2__N_3422;
    
    wire n45956, n55892, n45955;
    wire [23:0]n7771;
    
    wire n55884, n55888, n45954, n45953, n55890, n56310, n45952, 
        n45951, n56313, n55886, n56505, n56154, n56002, n45950, 
        n56417, n53248, n56567, n56124, n56086, n56084, n56024, 
        n59296, n62174, n48_adj_5129, n46;
    wire [23:0]n7615;
    
    wire n1697, n59776, n53212, n48_adj_5130, n56082, n56036, n45949, 
        n45948, n56028, n56164, n22999, n805, n55894, n42_adj_5131, 
        n804, n61687, n803, n61688, n53214, n48_adj_5132, n962, 
        n40_adj_5133, n961, n56066, n38068, n18_adj_5134, n45947, 
        n45946, n45945, n55684, n45944, n45943, n56491, n55712, 
        n56421, n56561, n45942, n56549, n59667;
    wire [23:0]n7641;
    
    wire n1835, n45941;
    wire [23:0]n7667;
    
    wire n1970, n44;
    wire [23:0]n7693;
    
    wire n2102;
    wire [23:0]n7719;
    
    wire n55366, n2476, n45940, n45939, n45938;
    wire [23:0]n7745;
    
    wire n45937, n22983, n59671, n19287, n45936, n42_adj_5135, n960, 
        n9427, n19289, n19237, n9263, n44_adj_5136, n959, n44_adj_5137, 
        n56156, n56080, n45935, n56431, n45934, n45933, n45932, 
        n45931;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index_c;   // verilog/uart_rx.v(34[17:28])
    
    wire n45930, n45929, n45928, n55860, n45927, n45926, n2104, 
        n35_adj_5145, n39_adj_5146, n2103, n37_adj_5147, n2101, n41_adj_5148, 
        n39_adj_5149, n2107, n29_adj_5150, n45925, n2106, n31_adj_5151, 
        n55364, n53462, n2353, n45924, n2105, n33_adj_5152, n2108, 
        n27_adj_5153, n45923, n60259, n45922, n45921, n45920, n45919, 
        n45918, n45917, n3_adj_5154, n30_adj_5155, n38_adj_5156, n53473, 
        n2109, n26_adj_5157, n61466, n61467, n45916, n60235, n28_adj_5158, 
        n60233, n61885, n60610, n62077, n56262, n56056, n2100, 
        n62078, n45915, n45914, n31_adj_5159, n19_adj_5160, n17_adj_5161, 
        n15_adj_5162, n59717, n13_adj_5163, n11_adj_5164, n60671, 
        n61215, n25_adj_5165, n23_adj_5166, n21_adj_5167, n61203, 
        n2099, n62023, n2098, n48_adj_5168, n55896, n38066, n55292, 
        n56158, n56106, n56166, n22947, n45913, n29_adj_5169, n27_adj_5170, 
        n59725, n8_adj_5171, n1971, n37_adj_5172, n54410, n45912, 
        n1972, n35_adj_5173, n1969, n41_adj_5174, n39_adj_5175, n1975, 
        n29_adj_5176, n56264, n1974, n31_adj_5177, n1973, n33_adj_5178, 
        n1976, n27_adj_5179, n59408, n56266, n22974, n30_adj_5180, 
        n38_adj_5181, n1977, n26_adj_5182, n61470, n61471, n60286, 
        n28_adj_5183, n60284, n61883, n60602, n62058, n1968, n62059, 
        n1967, n62027, n1966, n48_adj_5184, n2110, n46249, n45911, 
        n46248, n46247, n61657, n33_adj_5185, n61658, n46246, n45910, 
        n55362, n53466, n46245, n2227, n45909, n45908, n45907, 
        n45906, n46244, n45905, n45904, n46243, n45903, n45902, 
        n45901, n45900, n45899, n45898, n45897, n45896, n55360, 
        n53470, n45895, n45894, n45893, n45892, n45891, n45890, 
        n45889, n45888, n16_adj_5186, n34_adj_5187, n37_adj_5188, 
        n35_adj_5189, n59710, n45887, n55628, n45886, n45885, n45884, 
        n45883, n55646, n45882, n45881, n45880, n45879, n45878, 
        n45877, n45876, n45875, n45874, n45873, n45872, n3186, 
        n46058, n46057, n1831, n45871, n1832, n45870, n46056, 
        n46055, n1833, n45869, n46054, n1834, n45868, n46053, 
        n45867, n1836, n45866, n1837, n45865, n46052, n1838, n45864, 
        n14_adj_5190, n59697, n61988, n1839, n45863, n46051, n1840, 
        n45862, n1841, n45861, n46050, n55358, n53479, n1693, 
        n45860, n46049, n1694, n45859, n1695, n45858, n1696, n45857, 
        n46048, n45856, n46047, n1698, n45855, n1699, n45854, 
        n1700, n45853, n46046, n1701, n45852, n46045, n1702, n1552, 
        n45851, n1553, n45850, n46044, n1554, n45849, n1555, n45848, 
        n45847, n46043, n46042, n1557, n45846, n1558, n45845, 
        n1559, n45844, n46041, n1560, n45843, n56497, n56563, 
        n46040, n1408, n45842, n1409, n45841, n1410, n17_adj_5191, 
        n33_adj_5192, n21_adj_5193, n19_adj_5194, n15_adj_5195, n23_adj_5196, 
        n13_adj_5197, n19207, n41_adj_5198, n61672, n22938, n4_adj_5199, 
        n55802, n55834, n55722, n56503, n56292, n56529, n39_adj_5200, 
        n37_adj_5201, n43_adj_5202, n41_adj_5203, n31_adj_5204, n33_adj_5205, 
        n35_adj_5206, n29_adj_5207, n59432, n32_adj_5208, n40_adj_5209, 
        n28_adj_5210, n61667, n61668, n59428, n30_adj_5211, n59424, 
        n61665, n61523, n62037, n62038, n43_adj_5212, n37_adj_5213, 
        n41_adj_5214, n39_adj_5215, n53482, n32_adj_5216, n61675, 
        n61676, n59457, n60340, n34_adj_5217, n61209, n61519, n53990, 
        n61671, n48_adj_5218, n56134, n56136, n61544, n56290, n54622, 
        n55482, n55488, n53499, n42_adj_5219, n52133, n56453, n56555, 
        n2, n9643, n61685, n61686, n53216, n48_adj_5220, n43_adj_5221, 
        n37_adj_5222, n41_adj_5223, n39_adj_5224, n56094, n56092, 
        n22990, n32_adj_5225, n61679, n61680, n59476, n60358, n34_adj_5226, 
        n61207, n61515, n61677, n61678, n48_adj_5227, n10_adj_5228, 
        n61659, n56280, n61660, n59750, n60592, n12_adj_5229, n20_adj_5230, 
        n26_adj_5231, n34_adj_5232, n45_adj_5233, n39_adj_5234, n41_adj_5235, 
        n43_adj_5236, n61681, n61682, n59496, n60366, n36, n38_adj_5237, 
        n61494, n44_adj_5238, n61205, n62134, n55906, n61219, n55908, 
        n62154, n22962, n62155, n62141, n61221, n55950, n59234, 
        n59235, n42_adj_5239, n38_adj_5240, n59508, n56044, n3_adj_5241, 
        n9434, n56048, n5, n56052, n8_adj_5242, n55346, n59335, 
        n59332, n59329, n55440, n55446, n46_adj_5243, n55818, n59223, 
        n59229, n59220, n59226, n46_adj_5244, n14_adj_5245, n15_adj_5246, 
        n55880, n36_adj_5247, n40_adj_5248, n61984, n61985, n59786, 
        n60721, n55728, n61868, n61247, n61243, n10_adj_5249, n61423, 
        n55840, n55808, n55390, n55422, n36_adj_5251;
    
    SB_LUT4 add_2639_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n45839), 
            .O(n7589[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n46038), 
            .O(n7953[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_7 (.CI(n45839), .I0(n1411), .I1(n1460), .CO(n45840));
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n27247));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2653_5 (.CI(n46038), .I0(n3171), .I1(n698), .CO(n46039));
    SB_LUT4 add_2639_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n45838), 
            .O(n7589[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n46037), 
            .O(n7953[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_4 (.CI(n46037), .I0(n3172), .I1(n858), .CO(n46038));
    SB_CARRY add_2639_6 (.CI(n45838), .I0(n1412), .I1(n1011), .CO(n45839));
    SB_LUT4 add_2639_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n45837), 
            .O(n7589[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45760_3_lut (.I0(n61424), .I1(baudrate[15]), .I2(n37), .I3(GND_net), 
            .O(n60660));   // verilog/uart_rx.v(119[33:55])
    defparam i45760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2653_3_lut (.I0(n53438), .I1(GND_net), .I2(n538), .I3(n46036), 
            .O(n55376)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), .I3(n55824), 
            .O(n55830));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2653_3 (.CI(n46036), .I0(GND_net), .I1(n538), .CO(n46037));
    SB_CARRY add_2639_5 (.CI(n45837), .I0(n1413), .I1(n856), .CO(n45838));
    SB_LUT4 add_2639_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n45836), 
            .O(n7589[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_4 (.CI(n45836), .I0(n1414), .I1(n698), .CO(n45837));
    SB_CARRY add_2653_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n46036));
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2652_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n46035), 
            .O(n7927[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n27246));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2652_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n46034), 
            .O(n7927[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_22_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n27245));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2652_22 (.CI(n46034), .I0(n3047), .I1(n3188), .CO(n46035));
    SB_LUT4 add_2652_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n46033), 
            .O(n7927[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2639_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n45835), 
            .O(n7589[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_3 (.CI(n45835), .I0(n1415), .I1(n858), .CO(n45836));
    SB_CARRY add_2652_21 (.CI(n46033), .I0(n3048), .I1(n3084), .CO(n46034));
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n27243));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2652_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n46032), 
            .O(n7927[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41590_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n56481));
    defparam i41590_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i41646_4_lut (.I0(n56481), .I1(n56148), .I2(n56479), .I3(n56102), 
            .O(n56537));
    defparam i41646_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i41647_1_lut (.I0(n56537), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53446));
    defparam i41647_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n27242));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14), .I1(baudrate[9]), 
            .I2(n25), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(n56162), .I1(n55316), .I2(n55314), 
            .I3(n56152), .O(n22959));
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 i45340_4_lut (.I0(\o_Rx_DV_N_3464[8] ), .I1(\o_Rx_DV_N_3464[12] ), 
            .I2(n4855), .I3(n52352), .O(n59276));
    defparam i45340_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i38602_1_lut (.I0(n22959), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53458));
    defparam i38602_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45337_4_lut (.I0(n59276), .I1(\o_Rx_DV_N_3464[24] ), .I2(n29), 
            .I3(n23), .O(n59273));
    defparam i45337_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(r_SM_Main[1]), .I1(n59273), .I2(r_SM_Main_c[0]), 
            .I3(n27), .O(n25039));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n27241));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n27240));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n7953[20]), .I3(n294[1]), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n7953[19]), .I3(n294[1]), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55770), .O(n55776));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n7953[16]), .I3(n294[1]), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n7953[17]), .I3(n294[1]), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n7953[18]), .I3(n294[1]), .O(n37_adj_4979));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n7953[14]), .I3(n294[1]), .O(n29_adj_4980));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n7953[15]), .I3(n294[1]), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n7953[11]), .I3(n294[1]), .O(n23_adj_4981));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n62842));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i1_4_lut_adj_1009 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55776), .O(n55782));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hfffe;
    SB_LUT4 i47019_4_lut (.I0(n22), .I1(n12), .I2(n25), .I3(n59813), 
            .O(n61919));   // verilog/uart_rx.v(119[33:55])
    defparam i47019_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n7953[12]), .I3(n294[1]), .O(n25_adj_4982));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n7953[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n7953[22]), .I3(n294[1]), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n7953[21]), .I3(n294[1]), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n7953[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n7953[8]), .I3(n294[1]), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n7953[9]), .I3(n294[1]), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n7953[10]), .I3(n294[1]), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n7953[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n7953[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n7953[7]), .I3(n294[1]), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n7953[13]), .I3(n294[1]), .O(n27_adj_4983));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i44682_4_lut (.I0(n27_adj_4983), .I1(n15), .I2(n13), .I3(n11), 
            .O(n59582));
    defparam i44682_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i44694_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n59594));
    defparam i44694_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n55354), .I1(n48), .I2(GND_net), .I3(GND_net), 
            .O(n1415));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR r_Clock_Count_1943__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n25247), .D(n1[0]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_c[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i44636_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n59536));
    defparam i44636_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2652_20 (.CI(n46032), .I0(n3049), .I1(n2977), .CO(n46033));
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47020_3_lut (.I0(n61919), .I1(baudrate[10]), .I2(n27_adj_4985), 
            .I3(GND_net), .O(n61920));   // verilog/uart_rx.v(119[33:55])
    defparam i47020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n7953[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44706_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n59606));
    defparam i44706_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i45548_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n59606), 
            .O(n60448));
    defparam i45548_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_4_lut_adj_1010 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55786), .O(n55792));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 i45544_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n60448), 
            .O(n60444));
    defparam i45544_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55792), .O(n55798));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2639_2_lut (.I0(n53488), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55356)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i46843_4_lut (.I0(n25_adj_4982), .I1(n23_adj_4981), .I2(n21), 
            .I3(n60444), .O(n61743));
    defparam i46843_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2639_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45835));
    SB_LUT4 i46233_4_lut (.I0(n31), .I1(n29_adj_4980), .I2(n27_adj_4983), 
            .I3(n61743), .O(n61133));
    defparam i46233_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47047_4_lut (.I0(n37_adj_4979), .I1(n35), .I2(n33), .I3(n61133), 
            .O(n61947));
    defparam i47047_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33), .I3(GND_net), .O(n12_adj_4986));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41643_1_lut (.I0(n56533), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53496));
    defparam i41643_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n55376), .I3(n48_adj_4987), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i46741_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_adj_4983), 
            .I3(GND_net), .O(n61641));   // verilog/uart_rx.v(119[33:55])
    defparam i46741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n46031), 
            .O(n7927[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_19 (.CI(n46031), .I0(n3050), .I1(n2867), .CO(n46032));
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55738), .O(n55744));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i46742_3_lut (.I0(n61641), .I1(baudrate[14]), .I2(n29_adj_4980), 
            .I3(GND_net), .O(n61642));   // verilog/uart_rx.v(119[33:55])
    defparam i46742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44670_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n59570));
    defparam i44670_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55744), .O(n55750));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_4986), .I1(baudrate[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44674_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4980), .I3(n59582), 
            .O(n59574));
    defparam i44674_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47094_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n59570), 
            .O(n61994));   // verilog/uart_rx.v(119[33:55])
    defparam i47094_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46660_3_lut (.I0(n61642), .I1(baudrate[15]), .I2(n31), .I3(GND_net), 
            .O(n61560));   // verilog/uart_rx.v(119[33:55])
    defparam i46660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47238_4_lut (.I0(n61560), .I1(n61994), .I2(n35), .I3(n59574), 
            .O(n62138));   // verilog/uart_rx.v(119[33:55])
    defparam i47238_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2652_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n46030), 
            .O(n7927[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_18 (.CI(n46030), .I0(n3051), .I1(n2754), .CO(n46031));
    SB_LUT4 i47239_3_lut (.I0(n62138), .I1(baudrate[18]), .I2(n37_adj_4979), 
            .I3(GND_net), .O(n62139));   // verilog/uart_rx.v(119[33:55])
    defparam i47239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_4988));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46743_3_lut (.I0(n6_adj_4988), .I1(baudrate[10]), .I2(n21), 
            .I3(GND_net), .O(n61643));   // verilog/uart_rx.v(119[33:55])
    defparam i46743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46744_3_lut (.I0(n61643), .I1(baudrate[11]), .I2(n23_adj_4981), 
            .I3(GND_net), .O(n61644));   // verilog/uart_rx.v(119[33:55])
    defparam i46744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38586_1_lut (.I0(n22971), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53442));
    defparam i38586_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i44640_4_lut (.I0(n43), .I1(n25_adj_4982), .I2(n23_adj_4981), 
            .I3(n59594), .O(n59540));
    defparam i44640_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46325_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n59536), 
            .O(n61225));   // verilog/uart_rx.v(119[33:55])
    defparam i46325_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46658_3_lut (.I0(n61644), .I1(baudrate[12]), .I2(n25_adj_4982), 
            .I3(GND_net), .O(n61558));   // verilog/uart_rx.v(119[33:55])
    defparam i46658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47213_3_lut (.I0(n62139), .I1(baudrate[19]), .I2(n39), .I3(GND_net), 
            .O(n62113));   // verilog/uart_rx.v(119[33:55])
    defparam i47213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44646_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n61947), 
            .O(n59546));
    defparam i44646_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4989));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4990));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46917_4_lut (.I0(n61558), .I1(n61225), .I2(n45), .I3(n59540), 
            .O(n61817));   // verilog/uart_rx.v(119[33:55])
    defparam i46917_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47153_3_lut (.I0(n62113), .I1(baudrate[20]), .I2(n41), .I3(GND_net), 
            .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam i47153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4991));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4992));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4993));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4994));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4995));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4996));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4997));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n55328));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n7953[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n46029), 
            .O(n7927[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_17 (.CI(n46029), .I0(n3052), .I1(n2638), .CO(n46030));
    SB_LUT4 add_2652_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n46028), 
            .O(n7927[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46919_4_lut (.I0(n40), .I1(n61817), .I2(n45), .I3(n59546), 
            .O(n61819));   // verilog/uart_rx.v(119[33:55])
    defparam i46919_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(n56260), .I1(n56108), .I2(n55328), 
            .I3(n56104), .O(n55336));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4998));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2638_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n45834), 
            .O(n7563[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4999));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2638_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n45833), 
            .O(n7563[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5000));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2638_8 (.CI(n45833), .I0(n1262), .I1(n1459), .CO(n45834));
    SB_CARRY add_2652_16 (.CI(n46028), .I0(n3053), .I1(n2519), .CO(n46029));
    SB_LUT4 add_2638_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n45832), 
            .O(n7563[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5001));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2638_7 (.CI(n45832), .I0(n1263), .I1(n1460), .CO(n45833));
    SB_LUT4 i47405_4_lut (.I0(n55336), .I1(n61819), .I2(baudrate[23]), 
            .I3(n3253), .O(n54288));   // verilog/uart_rx.v(119[33:55])
    defparam i47405_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 add_2638_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n45831), 
            .O(n7563[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5002));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5003));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44971_4_lut (.I0(n35_adj_5001), .I1(n23_adj_5000), .I2(n21_adj_4999), 
            .I3(n19_adj_4998), .O(n59871));
    defparam i44971_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45901_4_lut (.I0(n17_adj_5003), .I1(n15_adj_5002), .I2(n2844), 
            .I3(baudrate[2]), .O(n60801));
    defparam i45901_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i46381_4_lut (.I0(n23_adj_5000), .I1(n21_adj_4999), .I2(n19_adj_4998), 
            .I3(n60801), .O(n61281));
    defparam i46381_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_2652_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n46027), 
            .O(n7927[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46373_4_lut (.I0(n29_adj_4997), .I1(n27_adj_4996), .I2(n25_adj_4995), 
            .I3(n61281), .O(n61273));
    defparam i46373_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i44978_4_lut (.I0(n35_adj_5001), .I1(n33_adj_4994), .I2(n31_adj_4993), 
            .I3(n61273), .O(n59878));
    defparam i44978_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55754), .O(n55760));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5004));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55760), .O(n55766));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hfffe;
    SB_CARRY add_2652_15 (.CI(n46027), .I0(n3054), .I1(n2397), .CO(n46028));
    SB_LUT4 add_2652_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n46026), 
            .O(n7927[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n7927[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46527_3_lut (.I0(n12_adj_5004), .I1(baudrate[13]), .I2(n35_adj_5001), 
            .I3(GND_net), .O(n61427));   // verilog/uart_rx.v(119[33:55])
    defparam i46527_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2638_6 (.CI(n45831), .I0(n1264), .I1(n1011), .CO(n45832));
    SB_LUT4 add_2638_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n45830), 
            .O(n7563[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n7927[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n7927[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2652_14 (.CI(n46026), .I0(n3055), .I1(n2272), .CO(n46027));
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20), .I1(baudrate[17]), 
            .I2(n43_adj_4991), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46528_3_lut (.I0(n61427), .I1(baudrate[14]), .I2(n37_adj_4990), 
            .I3(GND_net), .O(n61428));   // verilog/uart_rx.v(119[33:55])
    defparam i46528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n7927[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n7927[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2638_5 (.CI(n45830), .I0(n1265), .I1(n856), .CO(n45831));
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n7927[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n46025), 
            .O(n7927[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 i44959_4_lut (.I0(n41_adj_4992), .I1(n39_adj_4989), .I2(n37_adj_4990), 
            .I3(n59871), .O(n59859));
    defparam i44959_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2638_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n45829), 
            .O(n7563[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_4 (.CI(n45829), .I0(n1266), .I1(n698), .CO(n45830));
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2652_13 (.CI(n46025), .I0(n3056), .I1(n2144), .CO(n46026));
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n7927[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5005));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46957_4_lut (.I0(n38), .I1(n18), .I2(n43_adj_4991), .I3(n59853), 
            .O(n61857));   // verilog/uart_rx.v(119[33:55])
    defparam i46957_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n7901[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n7927[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45754_3_lut (.I0(n61428), .I1(baudrate[15]), .I2(n39_adj_4989), 
            .I3(GND_net), .O(n60654));   // verilog/uart_rx.v(119[33:55])
    defparam i45754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n46024), 
            .O(n7927[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n7901[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5006), .I1(baudrate[9]), 
            .I2(n27_adj_4996), .I3(GND_net), .O(n24_adj_5007));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47003_4_lut (.I0(n24_adj_5007), .I1(n14_adj_5008), .I2(n27_adj_4996), 
            .I3(n59896), .O(n61903));   // verilog/uart_rx.v(119[33:55])
    defparam i47003_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47004_3_lut (.I0(n61903), .I1(baudrate[10]), .I2(n29_adj_4997), 
            .I3(GND_net), .O(n61904));   // verilog/uart_rx.v(119[33:55])
    defparam i47004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5009));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n7927[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2652_12 (.CI(n46024), .I0(n3057), .I1(n2013), .CO(n46025));
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5010));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n7927[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2652_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n46023), 
            .O(n7927[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n7927[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n7927[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46836_3_lut (.I0(n61904), .I1(baudrate[11]), .I2(n31_adj_4993), 
            .I3(GND_net), .O(n61736));   // verilog/uart_rx.v(119[33:55])
    defparam i46836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46711_4_lut (.I0(n41_adj_4992), .I1(n39_adj_4989), .I2(n37_adj_4990), 
            .I3(n59878), .O(n61611));
    defparam i46711_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2652_11 (.CI(n46023), .I0(n3058), .I1(n1879), .CO(n46024));
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5012));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2638_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n45828), 
            .O(n7563[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_3 (.CI(n45828), .I0(n1267), .I1(n858), .CO(n45829));
    SB_LUT4 i47218_4_lut (.I0(n60654), .I1(n61857), .I2(n43_adj_4991), 
            .I3(n59859), .O(n62118));   // verilog/uart_rx.v(119[33:55])
    defparam i47218_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45752_3_lut (.I0(n61736), .I1(baudrate[12]), .I2(n33_adj_4994), 
            .I3(GND_net), .O(n60652));   // verilog/uart_rx.v(119[33:55])
    defparam i45752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n46022), 
            .O(n7927[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47244_4_lut (.I0(n60652), .I1(n62118), .I2(n43_adj_4991), 
            .I3(n61611), .O(n62144));   // verilog/uart_rx.v(119[33:55])
    defparam i47244_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n7901[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47245_3_lut (.I0(n62144), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n62145));   // verilog/uart_rx.v(119[33:55])
    defparam i47245_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n7927[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n7901[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n7927[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2652_10 (.CI(n46022), .I0(n3059), .I1(n1742), .CO(n46023));
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2652_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n46021), 
            .O(n7927[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2652_9 (.CI(n46021), .I0(n3060), .I1(n1602), .CO(n46022));
    SB_LUT4 add_2652_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n46020), 
            .O(n7927[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5018));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5019));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n7927[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n7927[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2638_2_lut (.I0(n53492), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55354)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2652_8 (.CI(n46020), .I0(n3061), .I1(n1459), .CO(n46021));
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2652_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n46019), 
            .O(n7927[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45048_4_lut (.I0(n37_adj_5031), .I1(n25_adj_5030), .I2(n23_adj_5029), 
            .I3(n21_adj_5028), .O(n59948));
    defparam i45048_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45947_4_lut (.I0(n19_adj_5027), .I1(n17_adj_5026), .I2(n2729), 
            .I3(baudrate[2]), .O(n60847));
    defparam i45947_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i46409_4_lut (.I0(n25_adj_5030), .I1(n23_adj_5029), .I2(n21_adj_5028), 
            .I3(n60847), .O(n61309));
    defparam i46409_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2652_7 (.CI(n46019), .I0(n3062), .I1(n1460), .CO(n46020));
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n7927[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46405_4_lut (.I0(n31_adj_5025), .I1(n29_adj_5024), .I2(n27_adj_5023), 
            .I3(n61309), .O(n61305));
    defparam i46405_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2652_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n46018), 
            .O(n7927[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45050_4_lut (.I0(n37_adj_5031), .I1(n35_adj_5022), .I2(n33_adj_5020), 
            .I3(n61305), .O(n59950));
    defparam i45050_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2652_6 (.CI(n46018), .I0(n3063), .I1(n1011), .CO(n46019));
    SB_CARRY add_2638_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45828));
    SB_LUT4 add_2637_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n45827), 
            .O(n7537[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n7927[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46533_3_lut (.I0(n14_adj_5034), .I1(baudrate[13]), .I2(n37_adj_5031), 
            .I3(GND_net), .O(n61433));   // verilog/uart_rx.v(119[33:55])
    defparam i46533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n7927[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46534_3_lut (.I0(n61433), .I1(baudrate[14]), .I2(n39_adj_5018), 
            .I3(GND_net), .O(n61434));   // verilog/uart_rx.v(119[33:55])
    defparam i46534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n7927[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2637_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n45826), 
            .O(n7537[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2652_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n46017), 
            .O(n7927[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_5 (.CI(n46017), .I0(n3064), .I1(n856), .CO(n46018));
    SB_CARRY add_2637_7 (.CI(n45826), .I0(n1112), .I1(n1460), .CO(n45827));
    SB_LUT4 add_2637_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n45825), 
            .O(n7537[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2652_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n46016), 
            .O(n7927[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2637_6 (.CI(n45825), .I0(n1113), .I1(n1011), .CO(n45826));
    SB_LUT4 add_2637_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n45824), 
            .O(n7537[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5035), .I1(baudrate[17]), 
            .I2(n45_adj_5017), .I3(GND_net), .O(n40_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2652_4 (.CI(n46016), .I0(n3065), .I1(n698), .CO(n46017));
    SB_LUT4 add_2652_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n46015), 
            .O(n7927[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45038_4_lut (.I0(n43_adj_5019), .I1(n41_adj_5015), .I2(n39_adj_5018), 
            .I3(n59948), .O(n59938));
    defparam i45038_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2652_3 (.CI(n46015), .I0(n3066), .I1(n858), .CO(n46016));
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46635_4_lut (.I0(n40_adj_5036), .I1(n20_adj_5039), .I2(n45_adj_5017), 
            .I3(n59934), .O(n61535));   // verilog/uart_rx.v(119[33:55])
    defparam i46635_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45748_3_lut (.I0(n61434), .I1(baudrate[15]), .I2(n41_adj_5015), 
            .I3(GND_net), .O(n60648));   // verilog/uart_rx.v(119[33:55])
    defparam i45748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2652_2_lut (.I0(n53442), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55374)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2652_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46015));
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5041), .I1(baudrate[9]), 
            .I2(n29_adj_5024), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47001_4_lut (.I0(n26), .I1(n16_adj_5042), .I2(n29_adj_5024), 
            .I3(n59960), .O(n61901));   // verilog/uart_rx.v(119[33:55])
    defparam i47001_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47002_3_lut (.I0(n61901), .I1(baudrate[10]), .I2(n31_adj_5025), 
            .I3(GND_net), .O(n61902));   // verilog/uart_rx.v(119[33:55])
    defparam i47002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46840_3_lut (.I0(n61902), .I1(baudrate[11]), .I2(n33_adj_5020), 
            .I3(GND_net), .O(n61740));   // verilog/uart_rx.v(119[33:55])
    defparam i46840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46725_4_lut (.I0(n43_adj_5019), .I1(n41_adj_5015), .I2(n39_adj_5018), 
            .I3(n59950), .O(n61625));
    defparam i46725_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44733_4_lut (.I0(n29_adj_5043), .I1(n17_adj_5040), .I2(n15_adj_5038), 
            .I3(n13_adj_5037), .O(n59633));
    defparam i44733_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47073_4_lut (.I0(n60648), .I1(n61535), .I2(n45_adj_5017), 
            .I3(n59938), .O(n61973));   // verilog/uart_rx.v(119[33:55])
    defparam i47073_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45658_4_lut (.I0(n11_adj_5032), .I1(n9_adj_5021), .I2(n3171), 
            .I3(baudrate[2]), .O(n60558));
    defparam i45658_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i45746_3_lut (.I0(n61740), .I1(baudrate[12]), .I2(n35_adj_5022), 
            .I3(GND_net), .O(n60646));   // verilog/uart_rx.v(119[33:55])
    defparam i45746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47075_4_lut (.I0(n60646), .I1(n61973), .I2(n45_adj_5017), 
            .I3(n61625), .O(n61975));   // verilog/uart_rx.v(119[33:55])
    defparam i47075_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46279_4_lut (.I0(n17_adj_5040), .I1(n15_adj_5038), .I2(n13_adj_5037), 
            .I3(n60558), .O(n61179));
    defparam i46279_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46277_4_lut (.I0(n23_adj_5016), .I1(n21_adj_5014), .I2(n19_adj_5033), 
            .I3(n61179), .O(n61177));
    defparam i46277_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i44739_4_lut (.I0(n29_adj_5043), .I1(n27_adj_5013), .I2(n25_adj_5012), 
            .I3(n61177), .O(n59639));
    defparam i44739_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n7875[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n7901[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46749_3_lut (.I0(n6_adj_5044), .I1(baudrate[13]), .I2(n29_adj_5043), 
            .I3(GND_net), .O(n61649));   // verilog/uart_rx.v(119[33:55])
    defparam i46749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2651_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n46014), 
            .O(n7901[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2637_5 (.CI(n45824), .I0(n1114), .I1(n856), .CO(n45825));
    SB_LUT4 add_2637_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n45823), 
            .O(n7537[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2651_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n46013), 
            .O(n7901[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2637_4 (.CI(n45823), .I0(n1115), .I1(n698), .CO(n45824));
    SB_CARRY add_2651_21 (.CI(n46013), .I0(n2939), .I1(n3084), .CO(n46014));
    SB_LUT4 add_2651_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n46012), 
            .O(n7901[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2637_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n45822), 
            .O(n7537[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_20 (.CI(n46012), .I0(n2940), .I1(n2977), .CO(n46013));
    SB_LUT4 add_2651_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n46011), 
            .O(n7901[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_19 (.CI(n46011), .I0(n2941), .I1(n2867), .CO(n46012));
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5046), .I1(baudrate[17]), 
            .I2(n37_adj_5010), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2637_3 (.CI(n45822), .I0(n1116), .I1(n858), .CO(n45823));
    SB_LUT4 add_2651_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n46010), 
            .O(n7901[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2637_2_lut (.I0(n53496), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55352)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2637_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2651_18 (.CI(n46010), .I0(n2942), .I1(n2754), .CO(n46011));
    SB_LUT4 add_2651_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n46009), 
            .O(n7901[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_17 (.CI(n46009), .I0(n2943), .I1(n2638), .CO(n46010));
    SB_LUT4 add_2651_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n46008), 
            .O(n7901[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_16 (.CI(n46008), .I0(n2944), .I1(n2519), .CO(n46009));
    SB_LUT4 i46750_3_lut (.I0(n61649), .I1(baudrate[14]), .I2(n31_adj_5009), 
            .I3(GND_net), .O(n61650));   // verilog/uart_rx.v(119[33:55])
    defparam i46750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2651_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n46007), 
            .O(n7901[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2637_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45822));
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2651_15 (.CI(n46007), .I0(n2945), .I1(n2397), .CO(n46008));
    SB_LUT4 add_2651_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n46006), 
            .O(n7901[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_14 (.CI(n46006), .I0(n2946), .I1(n2272), .CO(n46007));
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44728_4_lut (.I0(n35_adj_5011), .I1(n33_adj_5005), .I2(n31_adj_5009), 
            .I3(n59633), .O(n59628));
    defparam i44728_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47090_4_lut (.I0(n32), .I1(n12_adj_5049), .I2(n37_adj_5010), 
            .I3(n59625), .O(n61990));   // verilog/uart_rx.v(119[33:55])
    defparam i47090_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46650_3_lut (.I0(n61650), .I1(baudrate[15]), .I2(n33_adj_5005), 
            .I3(GND_net), .O(n61550));   // verilog/uart_rx.v(119[33:55])
    defparam i46650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2651_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n46005), 
            .O(n7901[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_13 (.CI(n46005), .I0(n2947), .I1(n2144), .CO(n46006));
    SB_LUT4 add_2651_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n46004), 
            .O(n7901[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46751_3_lut (.I0(n8_adj_5052), .I1(baudrate[10]), .I2(n23_adj_5016), 
            .I3(GND_net), .O(n61651));   // verilog/uart_rx.v(119[33:55])
    defparam i46751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46752_3_lut (.I0(n61651), .I1(baudrate[11]), .I2(n25_adj_5012), 
            .I3(GND_net), .O(n61652));   // verilog/uart_rx.v(119[33:55])
    defparam i46752_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2651_12 (.CI(n46004), .I0(n2948), .I1(n2013), .CO(n46005));
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2651_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n46003), 
            .O(n7901[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45640_4_lut (.I0(n25_adj_5012), .I1(n23_adj_5016), .I2(n21_adj_5014), 
            .I3(n59661), .O(n60540));
    defparam i45640_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46323_3_lut (.I0(n10_adj_5055), .I1(baudrate[9]), .I2(n21_adj_5014), 
            .I3(GND_net), .O(n61223));   // verilog/uart_rx.v(119[33:55])
    defparam i46323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46648_3_lut (.I0(n61652), .I1(baudrate[12]), .I2(n27_adj_5013), 
            .I3(GND_net), .O(n61548));   // verilog/uart_rx.v(119[33:55])
    defparam i46648_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2651_11 (.CI(n46003), .I0(n2949), .I1(n1879), .CO(n46004));
    SB_LUT4 add_2651_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n46002), 
            .O(n7901[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46572_4_lut (.I0(n35_adj_5011), .I1(n33_adj_5005), .I2(n31_adj_5009), 
            .I3(n59639), .O(n61472));
    defparam i46572_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2651_10 (.CI(n46002), .I0(n2950), .I1(n1742), .CO(n46003));
    SB_LUT4 i47236_4_lut (.I0(n61550), .I1(n61990), .I2(n37_adj_5010), 
            .I3(n59628), .O(n62136));   // verilog/uart_rx.v(119[33:55])
    defparam i47236_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2651_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n46001), 
            .O(n7901[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_9 (.CI(n46001), .I0(n2951), .I1(n1602), .CO(n46002));
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2651_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n46000), 
            .O(n7901[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46745_4_lut (.I0(n61548), .I1(n61223), .I2(n27_adj_5013), 
            .I3(n60540), .O(n61645));   // verilog/uart_rx.v(119[33:55])
    defparam i46745_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47252_4_lut (.I0(n61645), .I1(n62136), .I2(n37_adj_5010), 
            .I3(n61472), .O(n62152));   // verilog/uart_rx.v(119[33:55])
    defparam i47252_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47253_3_lut (.I0(n62152), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n62153));   // verilog/uart_rx.v(119[33:55])
    defparam i47253_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47243_3_lut (.I0(n62153), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n62143));   // verilog/uart_rx.v(119[33:55])
    defparam i47243_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2651_8 (.CI(n46000), .I0(n2952), .I1(n1459), .CO(n46001));
    SB_LUT4 i47011_3_lut (.I0(n62143), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n61911));   // verilog/uart_rx.v(119[33:55])
    defparam i47011_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2651_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n45999), 
            .O(n7901[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47012_3_lut (.I0(n61911), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n61912));   // verilog/uart_rx.v(119[33:55])
    defparam i47012_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46656_3_lut (.I0(n61912), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_4987));   // verilog/uart_rx.v(119[33:55])
    defparam i46656_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45114_4_lut (.I0(n23_adj_5060), .I1(n21_adj_5059), .I2(n19_adj_5058), 
            .I3(n17_adj_5062), .O(n60014));
    defparam i45114_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2651_7 (.CI(n45999), .I0(n2953), .I1(n1460), .CO(n46000));
    SB_LUT4 add_2651_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n45998), 
            .O(n7901[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45110_4_lut (.I0(n29_adj_5057), .I1(n27_adj_5056), .I2(n25_adj_5061), 
            .I3(n60014), .O(n60010));
    defparam i45110_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46735_4_lut (.I0(n35_adj_5054), .I1(n33_adj_5053), .I2(n31_adj_5051), 
            .I3(n60010), .O(n61635));
    defparam i46735_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2651_6 (.CI(n45998), .I0(n2954), .I1(n1011), .CO(n45999));
    SB_LUT4 add_2651_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n45997), 
            .O(n7901[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46539_3_lut (.I0(n16_adj_5063), .I1(baudrate[13]), .I2(n39_adj_5050), 
            .I3(GND_net), .O(n61439));   // verilog/uart_rx.v(119[33:55])
    defparam i46539_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2651_5 (.CI(n45997), .I0(n2955), .I1(n856), .CO(n45998));
    SB_LUT4 add_2651_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n45996), 
            .O(n7901[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_4 (.CI(n45996), .I0(n2956), .I1(n698), .CO(n45997));
    SB_LUT4 i46540_3_lut (.I0(n61439), .I1(baudrate[14]), .I2(n41_adj_5048), 
            .I3(GND_net), .O(n61440));   // verilog/uart_rx.v(119[33:55])
    defparam i46540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45961_4_lut (.I0(n41_adj_5048), .I1(n39_adj_5050), .I2(n27_adj_5056), 
            .I3(n60012), .O(n60861));
    defparam i45961_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46633_3_lut (.I0(n22_adj_5064), .I1(baudrate[7]), .I2(n27_adj_5056), 
            .I3(GND_net), .O(n61533));   // verilog/uart_rx.v(119[33:55])
    defparam i46633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45736_3_lut (.I0(n61440), .I1(baudrate[15]), .I2(n43_adj_5047), 
            .I3(GND_net), .O(n60636));   // verilog/uart_rx.v(119[33:55])
    defparam i45736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5065), .I1(baudrate[9]), 
            .I2(n31_adj_5051), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2651_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n45995), 
            .O(n7901[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46999_4_lut (.I0(n28), .I1(n18_adj_5066), .I2(n31_adj_5051), 
            .I3(n60008), .O(n61899));   // verilog/uart_rx.v(119[33:55])
    defparam i46999_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47000_3_lut (.I0(n61899), .I1(baudrate[10]), .I2(n33_adj_5053), 
            .I3(GND_net), .O(n61900));   // verilog/uart_rx.v(119[33:55])
    defparam i47000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46846_3_lut (.I0(n61900), .I1(baudrate[11]), .I2(n35_adj_5054), 
            .I3(GND_net), .O(n61746));   // verilog/uart_rx.v(119[33:55])
    defparam i46846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45967_4_lut (.I0(n41_adj_5048), .I1(n39_adj_5050), .I2(n37_adj_5045), 
            .I3(n61635), .O(n60867));
    defparam i45967_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2651_3 (.CI(n45995), .I0(n2957), .I1(n858), .CO(n45996));
    SB_LUT4 i46841_4_lut (.I0(n60636), .I1(n61533), .I2(n43_adj_5047), 
            .I3(n60861), .O(n61741));   // verilog/uart_rx.v(119[33:55])
    defparam i46841_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2651_2_lut (.I0(n53446), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55372)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i45734_3_lut (.I0(n61746), .I1(baudrate[12]), .I2(n37_adj_5045), 
            .I3(GND_net), .O(n60634));   // verilog/uart_rx.v(119[33:55])
    defparam i45734_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2651_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45995));
    SB_LUT4 i47116_4_lut (.I0(n60634), .I1(n61741), .I2(n43_adj_5047), 
            .I3(n60867), .O(n62016));   // verilog/uart_rx.v(119[33:55])
    defparam i47116_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2650_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n45994), 
            .O(n7875[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47117_3_lut (.I0(n62016), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n62017));   // verilog/uart_rx.v(119[33:55])
    defparam i47117_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2650_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n45993), 
            .O(n7875[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_20 (.CI(n45993), .I0(n2828), .I1(n2977), .CO(n45994));
    SB_LUT4 add_2650_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n45992), 
            .O(n7875[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_19 (.CI(n45992), .I0(n2829), .I1(n2867), .CO(n45993));
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n7849[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n7875[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2650_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n45991), 
            .O(n7875[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_18 (.CI(n45991), .I0(n2830), .I1(n2754), .CO(n45992));
    SB_LUT4 add_2650_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n45990), 
            .O(n7875[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_17 (.CI(n45990), .I0(n2831), .I1(n2638), .CO(n45991));
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n7901[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2650_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n45989), 
            .O(n7875[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_16 (.CI(n45989), .I0(n2832), .I1(n2519), .CO(n45990));
    SB_LUT4 add_2650_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n45988), 
            .O(n7875[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_15 (.CI(n45988), .I0(n2833), .I1(n2397), .CO(n45989));
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2650_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n45987), 
            .O(n7875[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_14 (.CI(n45987), .I0(n2834), .I1(n2272), .CO(n45988));
    SB_LUT4 add_2650_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n45986), 
            .O(n7875[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_13 (.CI(n45986), .I0(n2835), .I1(n2144), .CO(n45987));
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45163_4_lut (.I0(n25_adj_5078), .I1(n23_adj_5077), .I2(n21_adj_5076), 
            .I3(n19_adj_5080), .O(n60063));
    defparam i45163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45155_4_lut (.I0(n31_adj_5072), .I1(n29_adj_5071), .I2(n27_adj_5079), 
            .I3(n60063), .O(n60055));
    defparam i45155_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2650_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n45985), 
            .O(n7875[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n45671), .O(\o_Rx_DV_N_3464[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n55340), .I1(n22878), .I2(VCC_net), 
            .I3(n45670), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n45670), .I0(n22878), .I1(VCC_net), 
            .CO(n45671));
    SB_CARRY add_2650_12 (.CI(n45985), .I0(n2836), .I1(n2013), .CO(n45986));
    SB_LUT4 add_2650_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n45984), 
            .O(n7875[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n55416), .I1(n56571), .I2(VCC_net), 
            .I3(n45669), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_24 (.CI(n45669), .I0(n56571), .I1(VCC_net), 
            .CO(n45670));
    SB_CARRY add_2650_11 (.CI(n45984), .I0(n2837), .I1(n1879), .CO(n45985));
    SB_LUT4 i46769_4_lut (.I0(n37_adj_5075), .I1(n35_adj_5074), .I2(n33_adj_5073), 
            .I3(n60055), .O(n61669));
    defparam i46769_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3464[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n45668), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n45668), .I0(n294[21]), .I1(VCC_net), 
            .CO(n45669));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n55414), .I1(n294[20]), .I2(VCC_net), 
            .I3(n45667), .O(n55416)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_22 (.CI(n45667), .I0(n294[20]), .I1(VCC_net), 
            .CO(n45668));
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2650_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n45983), 
            .O(n7875[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46545_3_lut (.I0(n18_adj_5081), .I1(baudrate[13]), .I2(n41_adj_5069), 
            .I3(GND_net), .O(n61445));   // verilog/uart_rx.v(119[33:55])
    defparam i46545_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2650_10 (.CI(n45983), .I0(n2838), .I1(n1742), .CO(n45984));
    SB_LUT4 add_2650_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n45982), 
            .O(n7875[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46546_3_lut (.I0(n61445), .I1(baudrate[14]), .I2(n43_adj_5070), 
            .I3(GND_net), .O(n61446));   // verilog/uart_rx.v(119[33:55])
    defparam i46546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n55412), .I1(n294[19]), .I2(VCC_net), 
            .I3(n45666), .O(n55414)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2650_9 (.CI(n45982), .I0(n2839), .I1(n1602), .CO(n45983));
    SB_CARRY sub_38_add_2_21 (.CI(n45666), .I0(n294[19]), .I1(VCC_net), 
            .CO(n45667));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n45665), .O(o_Rx_DV_N_3464[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n45665), .I0(n294[18]), .I1(VCC_net), 
            .CO(n45666));
    SB_LUT4 add_2650_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n45981), 
            .O(n7875[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45987_4_lut (.I0(n43_adj_5070), .I1(n41_adj_5069), .I2(n29_adj_5071), 
            .I3(n60057), .O(n60887));
    defparam i45987_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2650_8 (.CI(n45981), .I0(n2840), .I1(n1459), .CO(n45982));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n55410), .I1(n294[17]), .I2(VCC_net), 
            .I3(n45664), .O(n55412)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_19 (.CI(n45664), .I0(n294[17]), .I1(VCC_net), 
            .CO(n45665));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n55408), .I1(n294[16]), .I2(VCC_net), 
            .I3(n45663), .O(n55410)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2650_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n45980), 
            .O(n7875[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_7 (.CI(n45980), .I0(n2841), .I1(n1460), .CO(n45981));
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5083), .I1(baudrate[7]), 
            .I2(n29_adj_5071), .I3(GND_net), .O(n26_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45730_3_lut (.I0(n61446), .I1(baudrate[15]), .I2(n45_adj_5068), 
            .I3(GND_net), .O(n60630));   // verilog/uart_rx.v(119[33:55])
    defparam i45730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2650_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n45979), 
            .O(n7875[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_6 (.CI(n45979), .I0(n2842), .I1(n1011), .CO(n45980));
    SB_LUT4 add_2650_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n45978), 
            .O(n7875[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_18 (.CI(n45663), .I0(n294[16]), .I1(VCC_net), 
            .CO(n45664));
    SB_LUT4 sub_38_add_2_17_lut (.I0(n55338), .I1(n294[15]), .I2(VCC_net), 
            .I3(n45662), .O(n55340)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n45662), .I0(n294[15]), .I1(VCC_net), 
            .CO(n45663));
    SB_CARRY add_2650_5 (.CI(n45978), .I0(n2843), .I1(n856), .CO(n45979));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n55406), .I1(n294[14]), .I2(VCC_net), 
            .I3(n45661), .O(n55408)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n45661), .I0(n294[14]), .I1(VCC_net), 
            .CO(n45662));
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3464[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n45660), .O(n55406)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2650_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n45977), 
            .O(n7875[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n45660), .I0(n294[13]), .I1(VCC_net), 
            .CO(n45661));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n45659), .O(\o_Rx_DV_N_3464[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_4 (.CI(n45977), .I0(n2844), .I1(n698), .CO(n45978));
    SB_CARRY sub_38_add_2_14 (.CI(n45659), .I0(n294[12]), .I1(VCC_net), 
            .CO(n45660));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3464[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n45658), .O(n55338)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n45658), .I0(n294[11]), .I1(VCC_net), 
            .CO(n45659));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n45657), .O(o_Rx_DV_N_3464[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2650_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n45976), 
            .O(n7875[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_3 (.CI(n45976), .I0(n2845), .I1(n858), .CO(n45977));
    SB_CARRY sub_38_add_2_12 (.CI(n45657), .I0(n294[10]), .I1(VCC_net), 
            .CO(n45658));
    SB_LUT4 add_2650_2_lut (.I0(n53450), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55370)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n45656), .O(o_Rx_DV_N_3464[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45976));
    SB_CARRY sub_38_add_2_11 (.CI(n45656), .I0(n294[9]), .I1(VCC_net), 
            .CO(n45657));
    SB_LUT4 add_2649_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n45975), 
            .O(n7849[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2649_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n45974), 
            .O(n7849[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n45655), .O(\o_Rx_DV_N_3464[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_19 (.CI(n45974), .I0(n2714), .I1(n2867), .CO(n45975));
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5085), .I1(baudrate[9]), 
            .I2(n33_adj_5073), .I3(GND_net), .O(n30_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46997_4_lut (.I0(n30_adj_5086), .I1(n20_adj_5087), .I2(n33_adj_5073), 
            .I3(n60045), .O(n61897));   // verilog/uart_rx.v(119[33:55])
    defparam i46997_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46998_3_lut (.I0(n61897), .I1(baudrate[10]), .I2(n35_adj_5074), 
            .I3(GND_net), .O(n61898));   // verilog/uart_rx.v(119[33:55])
    defparam i46998_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_10 (.CI(n45655), .I0(n294[8]), .I1(VCC_net), 
            .CO(n45656));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n45654), .O(\o_Rx_DV_N_3464[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n45654), .I0(n294[7]), .I1(VCC_net), 
            .CO(n45655));
    SB_LUT4 add_2649_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n45973), 
            .O(n7849[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_18 (.CI(n45973), .I0(n2715), .I1(n2754), .CO(n45974));
    SB_LUT4 i46848_3_lut (.I0(n61898), .I1(baudrate[11]), .I2(n37_adj_5075), 
            .I3(GND_net), .O(n61748));   // verilog/uart_rx.v(119[33:55])
    defparam i46848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45993_4_lut (.I0(n43_adj_5070), .I1(n41_adj_5069), .I2(n39_adj_5067), 
            .I3(n61669), .O(n60893));
    defparam i45993_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n45653), .O(\o_Rx_DV_N_3464[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n45653), .I0(n294[6]), .I1(VCC_net), 
            .CO(n45654));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n45652), .O(\o_Rx_DV_N_3464[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n45652), .I0(n294[5]), .I1(VCC_net), 
            .CO(n45653));
    SB_LUT4 add_2649_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n45972), 
            .O(n7849[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n45651), .O(\o_Rx_DV_N_3464[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_17 (.CI(n45972), .I0(n2716), .I1(n2638), .CO(n45973));
    SB_CARRY sub_38_add_2_6 (.CI(n45651), .I0(n294[4]), .I1(VCC_net), 
            .CO(n45652));
    SB_LUT4 add_2649_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n45971), 
            .O(n7849[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46630_4_lut (.I0(n60630), .I1(n26_adj_5084), .I2(n45_adj_5068), 
            .I3(n60887), .O(n61530));   // verilog/uart_rx.v(119[33:55])
    defparam i46630_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45728_3_lut (.I0(n61748), .I1(baudrate[12]), .I2(n39_adj_5067), 
            .I3(GND_net), .O(n60628));   // verilog/uart_rx.v(119[33:55])
    defparam i45728_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2649_16 (.CI(n45971), .I0(n2717), .I1(n2519), .CO(n45972));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n45650), .O(\o_Rx_DV_N_3464[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2649_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n45970), 
            .O(n7849[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n45650), .I0(n294[3]), .I1(VCC_net), 
            .CO(n45651));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n45649), .O(\o_Rx_DV_N_3464[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_15 (.CI(n45970), .I0(n2718), .I1(n2397), .CO(n45971));
    SB_LUT4 add_2649_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n45969), 
            .O(n7849[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n45649), .I0(n294[2]), .I1(VCC_net), 
            .CO(n45650));
    SB_CARRY add_2649_14 (.CI(n45969), .I0(n2719), .I1(n2272), .CO(n45970));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n45648), .O(\o_Rx_DV_N_3464[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n45648), .I0(n294[1]), .I1(VCC_net), 
            .CO(n45649));
    SB_LUT4 i38594_1_lut (.I0(n22965), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53450));
    defparam i38594_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n54288), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3464[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n54288), .I1(GND_net), 
            .CO(n45648));
    SB_LUT4 i46632_4_lut (.I0(n60628), .I1(n61530), .I2(n45_adj_5068), 
            .I3(n60893), .O(n61532));   // verilog/uart_rx.v(119[33:55])
    defparam i46632_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n7823[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2649_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n45968), 
            .O(n7849[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n7849[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n7875[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n7901[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2649_13 (.CI(n45968), .I0(n2720), .I1(n2144), .CO(n45969));
    SB_LUT4 add_2649_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n45967), 
            .O(n7849[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46832_3_lut (.I0(n61920), .I1(baudrate[11]), .I2(n29_adj_5088), 
            .I3(GND_net), .O(n61732));   // verilog/uart_rx.v(119[33:55])
    defparam i46832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46677_4_lut (.I0(n39_adj_5089), .I1(n37), .I2(n35_adj_5090), 
            .I3(n59790), .O(n61577));
    defparam i46677_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2649_12 (.CI(n45967), .I0(n2721), .I1(n2013), .CO(n45968));
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7537[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5093), .I1(baudrate[4]), 
            .I2(n43_adj_5082), .I3(GND_net), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46783_4_lut (.I0(n42), .I1(n38_adj_5091), .I2(n43_adj_5082), 
            .I3(n59521), .O(n61683));   // verilog/uart_rx.v(119[33:55])
    defparam i46783_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46784_3_lut (.I0(n61683), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n61684));   // verilog/uart_rx.v(119[33:55])
    defparam i46784_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45234_4_lut (.I0(n27_adj_5102), .I1(n25_adj_5101), .I2(n23_adj_5100), 
            .I3(n21_adj_5103), .O(n60134));
    defparam i45234_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7563[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45223_4_lut (.I0(n33_adj_5099), .I1(n31_adj_5098), .I2(n29_adj_5097), 
            .I3(n60134), .O(n60123));
    defparam i45223_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5105), .I1(baudrate[7]), 
            .I2(n31_adj_5098), .I3(GND_net), .O(n28_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5107), .I1(baudrate[9]), 
            .I2(n35_adj_5096), .I3(GND_net), .O(n32_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46991_4_lut (.I0(n32_adj_5108), .I1(n22_adj_5109), .I2(n35_adj_5096), 
            .I3(n60121), .O(n61891));   // verilog/uart_rx.v(119[33:55])
    defparam i46991_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46992_3_lut (.I0(n61891), .I1(baudrate[10]), .I2(n37_adj_5095), 
            .I3(GND_net), .O(n61892));   // verilog/uart_rx.v(119[33:55])
    defparam i46992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46852_3_lut (.I0(n61892), .I1(baudrate[11]), .I2(n39_adj_5094), 
            .I3(GND_net), .O(n61752));   // verilog/uart_rx.v(119[33:55])
    defparam i46852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46801_4_lut (.I0(n39_adj_5094), .I1(n37_adj_5095), .I2(n35_adj_5096), 
            .I3(n60123), .O(n61701));
    defparam i46801_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47086_4_lut (.I0(n28_adj_5106), .I1(n20_adj_5104), .I2(n31_adj_5098), 
            .I3(n60129), .O(n61986));   // verilog/uart_rx.v(119[33:55])
    defparam i47086_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45724_3_lut (.I0(n61752), .I1(baudrate[12]), .I2(n41_adj_5092), 
            .I3(GND_net), .O(n60624));   // verilog/uart_rx.v(119[33:55])
    defparam i45724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47156_4_lut (.I0(n60624), .I1(n61986), .I2(n41_adj_5092), 
            .I3(n61701), .O(n62056));   // verilog/uart_rx.v(119[33:55])
    defparam i47156_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47157_3_lut (.I0(n62056), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n62057));   // verilog/uart_rx.v(119[33:55])
    defparam i47157_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47129_3_lut (.I0(n62057), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n62029));   // verilog/uart_rx.v(119[33:55])
    defparam i47129_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n7797[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n7823[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n7849[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n7875[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n7901[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2649_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n45966), 
            .O(n7849[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_11 (.CI(n45966), .I0(n2722), .I1(n1879), .CO(n45967));
    SB_LUT4 add_2649_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n45965), 
            .O(n7849[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7563[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2649_10 (.CI(n45965), .I0(n2723), .I1(n1742), .CO(n45966));
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45308_4_lut (.I0(n29_adj_5119), .I1(n27_adj_5118), .I2(n25_adj_5117), 
            .I3(n23_adj_5121), .O(n60208));
    defparam i45308_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2649_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n45964), 
            .O(n7849[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45280_4_lut (.I0(n35_adj_5116), .I1(n33_adj_5115), .I2(n31_adj_5114), 
            .I3(n60208), .O(n60180));
    defparam i45280_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2649_9 (.CI(n45964), .I0(n2724), .I1(n1602), .CO(n45965));
    SB_LUT4 add_2649_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n45963), 
            .O(n7849[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47190_4_lut (.I0(n60660), .I1(n61921), .I2(n41_adj_5122), 
            .I3(n59781), .O(n62090));   // verilog/uart_rx.v(119[33:55])
    defparam i47190_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45758_3_lut (.I0(n61732), .I1(baudrate[12]), .I2(n31_adj_5123), 
            .I3(GND_net), .O(n60658));   // verilog/uart_rx.v(119[33:55])
    defparam i45758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47256_4_lut (.I0(n60658), .I1(n62090), .I2(n41_adj_5122), 
            .I3(n61577), .O(n62156));   // verilog/uart_rx.v(119[33:55])
    defparam i47256_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47257_3_lut (.I0(n62156), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n62157));   // verilog/uart_rx.v(119[33:55])
    defparam i47257_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5125), .I1(baudrate[7]), 
            .I2(n33_adj_5115), .I3(GND_net), .O(n30_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2649_8 (.CI(n45963), .I0(n2725), .I1(n1459), .CO(n45964));
    SB_LUT4 add_2649_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n45962), 
            .O(n7849[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_7 (.CI(n45962), .I0(n2726), .I1(n1460), .CO(n45963));
    SB_LUT4 add_2649_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n45961), 
            .O(n7849[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47249_3_lut (.I0(n62157), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n62149));   // verilog/uart_rx.v(119[33:55])
    defparam i47249_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2649_6 (.CI(n45961), .I0(n2727), .I1(n1011), .CO(n45962));
    SB_LUT4 add_2649_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n45960), 
            .O(n7849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_5 (.CI(n45960), .I0(n2728), .I1(n856), .CO(n45961));
    SB_LUT4 add_2649_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n45959), 
            .O(n7849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_4 (.CI(n45959), .I0(n2729), .I1(n698), .CO(n45960));
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7589[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2649_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n45958), 
            .O(n7849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5127), .I1(baudrate[9]), 
            .I2(n37_adj_5113), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n7927[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46989_4_lut (.I0(n34), .I1(n24_adj_5128), .I2(n37_adj_5113), 
            .I3(n60178), .O(n61889));   // verilog/uart_rx.v(119[33:55])
    defparam i46989_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n56148));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'heeee;
    SB_LUT4 i46990_3_lut (.I0(n61889), .I1(baudrate[10]), .I2(n39_adj_5111), 
            .I3(GND_net), .O(n61890));   // verilog/uart_rx.v(119[33:55])
    defparam i46990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46854_3_lut (.I0(n61890), .I1(baudrate[11]), .I2(n41_adj_5112), 
            .I3(GND_net), .O(n61754));   // verilog/uart_rx.v(119[33:55])
    defparam i46854_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2649_3 (.CI(n45958), .I0(n2730), .I1(n858), .CO(n45959));
    SB_LUT4 i46811_4_lut (.I0(n41_adj_5112), .I1(n39_adj_5111), .I2(n37_adj_5113), 
            .I3(n60180), .O(n61711));
    defparam i46811_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46763_4_lut (.I0(n30_adj_5126), .I1(n22_adj_5124), .I2(n33_adj_5115), 
            .I3(n60194), .O(n61663));   // verilog/uart_rx.v(119[33:55])
    defparam i46763_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45720_3_lut (.I0(n61754), .I1(baudrate[12]), .I2(n43_adj_5110), 
            .I3(GND_net), .O(n60620));   // verilog/uart_rx.v(119[33:55])
    defparam i45720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2649_2_lut (.I0(n53454), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55368)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2649_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45958));
    SB_LUT4 i1_2_lut_adj_1019 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n56150));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(baudrate[24]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n56108));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n56102));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'heeee;
    SB_LUT4 i46961_4_lut (.I0(n60620), .I1(n61663), .I2(n43_adj_5110), 
            .I3(n61711), .O(n61861));   // verilog/uart_rx.v(119[33:55])
    defparam i46961_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46962_3_lut (.I0(n61861), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n61862));   // verilog/uart_rx.v(119[33:55])
    defparam i46962_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2648_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n45957), 
            .O(n7823[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47305_2_lut_3_lut_4_lut (.I0(r_SM_Main_2__N_3422[1]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main_c[0]), .I3(\r_SM_Main[2] ), .O(n25264));
    defparam i47305_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 add_2648_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n45956), 
            .O(n7823[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_18 (.CI(n45956), .I0(n2597), .I1(n2754), .CO(n45957));
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n55892));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 add_2648_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n45955), 
            .O(n7823[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_17 (.CI(n45955), .I0(n2598), .I1(n2638), .CO(n45956));
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n7771[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n55884));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n55888));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n56152));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 add_2648_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n45954), 
            .O(n7823[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_16 (.CI(n45954), .I0(n2599), .I1(n2519), .CO(n45955));
    SB_LUT4 add_2648_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n45953), 
            .O(n7823[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_15 (.CI(n45953), .I0(n2600), .I1(n2397), .CO(n45954));
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n7797[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n55890));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'heeee;
    SB_LUT4 i41421_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n56310));
    defparam i41421_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n7823[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2648_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n45952), 
            .O(n7823[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_14 (.CI(n45952), .I0(n2601), .I1(n2272), .CO(n45953));
    SB_LUT4 add_2648_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n45951), 
            .O(n7823[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n7849[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2648_13 (.CI(n45951), .I0(n2602), .I1(n2144), .CO(n45952));
    SB_LUT4 i1_2_lut_adj_1027 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56313));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'heeee;
    SB_LUT4 i41614_4_lut (.I0(n55890), .I1(n55886), .I2(n55888), .I3(n55884), 
            .O(n56505));
    defparam i41614_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n56154));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n56002));
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2648_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n45950), 
            .O(n7823[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n7875[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n7901[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41676_4_lut (.I0(n56537), .I1(n56417), .I2(n53248), .I3(baudrate[4]), 
            .O(n56567));
    defparam i41676_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47402_4_lut (.I0(n56505), .I1(n56313), .I2(n56567), .I3(n56310), 
            .O(n56571));
    defparam i47402_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_2648_12 (.CI(n45950), .I0(n2603), .I1(n2013), .CO(n45951));
    SB_LUT4 i1_3_lut (.I0(n56002), .I1(n56162), .I2(n56124), .I3(GND_net), 
            .O(n22965));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n56086));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n56084));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n56024));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n59296), .I1(baudrate[2]), 
            .I2(n62174), .I3(n48_adj_5129), .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7615[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44876_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n59776));
    defparam i44876_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46), .I1(baudrate[3]), .I2(n53212), 
            .I3(GND_net), .O(n48_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(n56024), .I1(n56084), .I2(n56086), 
            .I3(n56082), .O(n56036));
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2648_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n45949), 
            .O(n7823[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_11 (.CI(n45949), .I0(n2604), .I1(n1879), .CO(n45950));
    SB_LUT4 add_2648_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n45948), 
            .O(n7823[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n56036), .I1(n22965), .I2(n56028), 
            .I3(n56164), .O(n22999));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1035 (.I0(n22999), .I1(n48_adj_5130), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1035.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n55894));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46787_3_lut (.I0(n42_adj_5131), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n61687));   // verilog/uart_rx.v(119[33:55])
    defparam i46787_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46788_3_lut (.I0(n61687), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n61688));   // verilog/uart_rx.v(119[33:55])
    defparam i46788_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46603_3_lut (.I0(n61688), .I1(baudrate[4]), .I2(n53214), 
            .I3(GND_net), .O(n48_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam i46603_3_lut.LUT_INIT = 16'he8e8;
    SB_CARRY add_2648_10 (.CI(n45948), .I0(n2605), .I1(n1742), .CO(n45949));
    SB_LUT4 i41588_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n56479));
    defparam i41588_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4093_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam i4093_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n56066));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5133), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i24480_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38068));
    defparam i24480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2648_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n45947), 
            .O(n7823[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_9 (.CI(n45947), .I0(n2606), .I1(n1602), .CO(n45948));
    SB_LUT4 add_2648_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n45946), 
            .O(n7823[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_8 (.CI(n45946), .I0(n2607), .I1(n1459), .CO(n45947));
    SB_LUT4 add_2648_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n45945), 
            .O(n7823[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_7 (.CI(n45945), .I0(n2608), .I1(n1460), .CO(n45946));
    SB_LUT4 i1_4_lut_adj_1037 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n55684));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h0100;
    SB_LUT4 add_2648_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n45944), 
            .O(n7823[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_6 (.CI(n45944), .I0(n2609), .I1(n1011), .CO(n45945));
    SB_LUT4 add_2648_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n45943), 
            .O(n7823[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41600_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n56491));
    defparam i41600_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(n53248), .I1(n55684), .I2(n56260), 
            .I3(baudrate[16]), .O(n55712));
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'h0004;
    SB_CARRY add_2648_5 (.CI(n45943), .I0(n2610), .I1(n856), .CO(n45944));
    SB_LUT4 i41670_4_lut (.I0(n56491), .I1(n56417), .I2(n56421), .I3(n56313), 
            .O(n56561));
    defparam i41670_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2648_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n45942), 
            .O(n7823[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47274_4_lut (.I0(n56549), .I1(n59667), .I2(n56561), .I3(n55712), 
            .O(n62174));
    defparam i47274_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n7641[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2648_4 (.CI(n45942), .I0(n2611), .I1(n698), .CO(n45943));
    SB_LUT4 add_2648_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n45941), 
            .O(n7823[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_3 (.CI(n45941), .I0(n2612), .I1(n858), .CO(n45942));
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n7667[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i535_4_lut (.I0(n62174), .I1(n44), .I2(n294[20]), .I3(baudrate[2]), 
            .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n7693[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n7719[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n27583));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n48661));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n27579));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2648_2_lut (.I0(n53458), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55366)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2648_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45941));
    SB_LUT4 add_2647_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n45940), 
            .O(n7797[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2647_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n45939), 
            .O(n7797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_17 (.CI(n45939), .I0(n2477), .I1(n2638), .CO(n45940));
    SB_LUT4 add_2647_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n45938), 
            .O(n7797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_16 (.CI(n45938), .I0(n2478), .I1(n2519), .CO(n45939));
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n7745[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2647_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n45937), 
            .O(n7797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45261_4_lut (.I0(n22983), .I1(n59671), .I2(n48_adj_5129), 
            .I3(baudrate[0]), .O(n804));
    defparam i45261_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i5883_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n19287));   // verilog/uart_rx.v(119[33:55])
    defparam i5883_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n7771[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2647_15 (.CI(n45937), .I0(n2479), .I1(n2397), .CO(n45938));
    SB_LUT4 add_2647_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n45936), 
            .O(n7797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5135), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n7797[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5884_4_lut (.I0(n960), .I1(n9427), .I2(n19287), .I3(baudrate[3]), 
            .O(n19289));   // verilog/uart_rx.v(119[33:55])
    defparam i5884_4_lut.LUT_INIT = 16'ha8aa;
    SB_CARRY add_2647_14 (.CI(n45936), .I0(n2480), .I1(n2272), .CO(n45937));
    SB_LUT4 i3937_2_lut (.I0(n19237), .I1(n9263), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam i3937_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n7823[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5136), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5137), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n7849[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n56156));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n56080));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n56082));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 add_2647_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n45935), 
            .O(n7797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_13 (.CI(n45935), .I0(n2481), .I1(n2144), .CO(n45936));
    SB_LUT4 i38399_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n53248));
    defparam i38399_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41541_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56431));
    defparam i41541_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n7875[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2647_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n45934), 
            .O(n7797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_12 (.CI(n45934), .I0(n2482), .I1(n2013), .CO(n45935));
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n7901[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2647_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n45933), 
            .O(n7797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41658_4_lut (.I0(n56431), .I1(n56028), .I2(n56082), .I3(baudrate[9]), 
            .O(n56549));
    defparam i41658_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2647_11 (.CI(n45933), .I0(n2483), .I1(n1879), .CO(n45934));
    SB_LUT4 add_2647_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n45932), 
            .O(n7797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_10 (.CI(n45932), .I0(n2484), .I1(n1742), .CO(n45933));
    SB_LUT4 add_2647_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n45931), 
            .O(n7797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_9 (.CI(n45931), .I0(n2485), .I1(n1602), .CO(n45932));
    SB_DFFESR r_Clock_Count_1943__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n25247), .D(n1[7]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n25247), .D(n1[6]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n25247), .D(n1[5]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n25247), .D(n1[4]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n25247), .D(n1[3]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n25247), .D(n1[2]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1943__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n25247), .D(n1[1]), .R(n26549));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(clk16MHz), .E(n25264), 
            .D(n479[1]), .R(n53350));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(clk16MHz), .E(n25264), 
            .D(n479[2]), .R(n53350));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2647_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n45930), 
            .O(n7797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_8 (.CI(n45930), .I0(n2486), .I1(n1459), .CO(n45931));
    SB_LUT4 add_2647_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n45929), 
            .O(n7797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_7 (.CI(n45929), .I0(n2487), .I1(n1460), .CO(n45930));
    SB_LUT4 add_2647_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n45928), 
            .O(n7797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_6 (.CI(n45928), .I0(n2488), .I1(n1011), .CO(n45929));
    SB_LUT4 i1_2_lut_adj_1042 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n55860));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'heeee;
    SB_LUT4 add_2647_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n45927), 
            .O(n7797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_5 (.CI(n45927), .I0(n2489), .I1(n856), .CO(n45928));
    SB_LUT4 add_2647_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n45926), 
            .O(n7797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2647_4 (.CI(n45926), .I0(n2490), .I1(n698), .CO(n45927));
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2647_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n45925), 
            .O(n7797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_3 (.CI(n45925), .I0(n2491), .I1(n858), .CO(n45926));
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2647_2_lut (.I0(n53462), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55364)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2647_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45925));
    SB_LUT4 add_2646_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n45924), 
            .O(n7771[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2646_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n45923), 
            .O(n7771[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45359_4_lut (.I0(n33_adj_5152), .I1(n31_adj_5151), .I2(n29_adj_5150), 
            .I3(n27_adj_5153), .O(n60259));
    defparam i45359_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2646_16 (.CI(n45923), .I0(n2354), .I1(n2519), .CO(n45924));
    SB_LUT4 add_2646_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n45922), 
            .O(n7771[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_15 (.CI(n45922), .I0(n2355), .I1(n2397), .CO(n45923));
    SB_LUT4 add_2646_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n45921), 
            .O(n7771[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_14 (.CI(n45921), .I0(n2356), .I1(n2272), .CO(n45922));
    SB_LUT4 add_2646_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n45920), 
            .O(n7771[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_13 (.CI(n45920), .I0(n2357), .I1(n2144), .CO(n45921));
    SB_LUT4 add_2646_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n45919), 
            .O(n7771[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n7901[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2646_12 (.CI(n45919), .I0(n2358), .I1(n2013), .CO(n45920));
    SB_LUT4 add_2646_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n45918), 
            .O(n7771[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_11 (.CI(n45918), .I0(n2359), .I1(n1879), .CO(n45919));
    SB_LUT4 add_2646_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n45917), 
            .O(n7771[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_10 (.CI(n45917), .I0(n2360), .I1(n1742), .CO(n45918));
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5154), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5155), .I1(baudrate[10]), 
            .I2(n41_adj_5148), .I3(GND_net), .O(n38_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24523_rep_4_2_lut (.I0(n7693[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n53473));   // verilog/uart_rx.v(119[33:55])
    defparam i24523_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n53473), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i46566_3_lut (.I0(n26_adj_5157), .I1(baudrate[6]), .I2(n33_adj_5152), 
            .I3(GND_net), .O(n61466));   // verilog/uart_rx.v(119[33:55])
    defparam i46566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46567_3_lut (.I0(n61466), .I1(baudrate[7]), .I2(n35_adj_5145), 
            .I3(GND_net), .O(n61467));   // verilog/uart_rx.v(119[33:55])
    defparam i46567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2646_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n45916), 
            .O(n7771[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45335_4_lut (.I0(n39_adj_5149), .I1(n37_adj_5147), .I2(n35_adj_5145), 
            .I3(n60259), .O(n60235));
    defparam i45335_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46985_4_lut (.I0(n38_adj_5156), .I1(n28_adj_5158), .I2(n41_adj_5148), 
            .I3(n60233), .O(n61885));   // verilog/uart_rx.v(119[33:55])
    defparam i46985_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45710_3_lut (.I0(n61467), .I1(baudrate[8]), .I2(n37_adj_5147), 
            .I3(GND_net), .O(n60610));   // verilog/uart_rx.v(119[33:55])
    defparam i45710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47177_4_lut (.I0(n60610), .I1(n61885), .I2(n41_adj_5148), 
            .I3(n60235), .O(n62077));   // verilog/uart_rx.v(119[33:55])
    defparam i47177_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n56262), .I1(n56066), .I2(n56148), 
            .I3(n56056), .O(n22971));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'hfffe;
    SB_LUT4 i47178_3_lut (.I0(n62077), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n62078));   // verilog/uart_rx.v(119[33:55])
    defparam i47178_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2646_9 (.CI(n45916), .I0(n2361), .I1(n1602), .CO(n45917));
    SB_LUT4 add_2646_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n45915), 
            .O(n7771[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_8 (.CI(n45915), .I0(n2362), .I1(n1459), .CO(n45916));
    SB_LUT4 add_2646_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n45914), 
            .O(n7771[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i44817_4_lut (.I0(n31_adj_5159), .I1(n19_adj_5160), .I2(n17_adj_5161), 
            .I3(n15_adj_5162), .O(n59717));
    defparam i44817_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45771_4_lut (.I0(n13_adj_5163), .I1(n11_adj_5164), .I2(n3065), 
            .I3(baudrate[2]), .O(n60671));
    defparam i45771_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i46315_4_lut (.I0(n19_adj_5160), .I1(n17_adj_5161), .I2(n15_adj_5162), 
            .I3(n60671), .O(n61215));
    defparam i46315_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46303_4_lut (.I0(n25_adj_5165), .I1(n23_adj_5166), .I2(n21_adj_5167), 
            .I3(n61215), .O(n61203));
    defparam i46303_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47123_3_lut (.I0(n62078), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n62023));   // verilog/uart_rx.v(119[33:55])
    defparam i47123_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45716_3_lut (.I0(n62023), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam i45716_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(baudrate[17]), .I1(n55896), .I2(baudrate[2]), 
            .I3(n38066), .O(n55292));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'h0100;
    SB_CARRY add_2646_7 (.CI(n45914), .I0(n2363), .I1(n1460), .CO(n45915));
    SB_LUT4 i1_4_lut_adj_1045 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n56158));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1046 (.I0(n56106), .I1(n56156), .I2(n55860), 
            .I3(GND_net), .O(n56166));
    defparam i1_3_lut_adj_1046.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(n56166), .I1(n56162), .I2(n56164), 
            .I3(n56158), .O(n22947));
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1048 (.I0(n22947), .I1(n48_adj_5168), .I2(n538), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1048.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n7745[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n7771[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n7797[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n7823[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n7849[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2646_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n45913), 
            .O(n7771[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n7875[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i44825_4_lut (.I0(n31_adj_5159), .I1(n29_adj_5169), .I2(n27_adj_5170), 
            .I3(n61203), .O(n59725));
    defparam i44825_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n7901[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2646_6 (.CI(n45913), .I0(n2364), .I1(n1011), .CO(n45914));
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(n56505), .I1(n55292), .I2(n22959), 
            .I3(n56417), .O(n54410));
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'h0004;
    SB_LUT4 add_2646_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n45912), 
            .O(n7771[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n56262));
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n56104));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n56264));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n56260));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44508_4_lut (.I0(n33_adj_5178), .I1(n31_adj_5177), .I2(n29_adj_5176), 
            .I3(n27_adj_5179), .O(n59408));
    defparam i44508_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1054 (.I0(n56264), .I1(n56266), .I2(n56104), 
            .I3(n56262), .O(n22974));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5180), .I1(baudrate[9]), 
            .I2(n41_adj_5174), .I3(GND_net), .O(n38_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46570_3_lut (.I0(n26_adj_5182), .I1(baudrate[5]), .I2(n33_adj_5178), 
            .I3(GND_net), .O(n61470));   // verilog/uart_rx.v(119[33:55])
    defparam i46570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46571_3_lut (.I0(n61470), .I1(baudrate[6]), .I2(n35_adj_5173), 
            .I3(GND_net), .O(n61471));   // verilog/uart_rx.v(119[33:55])
    defparam i46571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45386_4_lut (.I0(n39_adj_5175), .I1(n37_adj_5172), .I2(n35_adj_5173), 
            .I3(n59408), .O(n60286));
    defparam i45386_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46983_4_lut (.I0(n38_adj_5181), .I1(n28_adj_5183), .I2(n41_adj_5174), 
            .I3(n60284), .O(n61883));   // verilog/uart_rx.v(119[33:55])
    defparam i46983_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45702_3_lut (.I0(n61471), .I1(baudrate[7]), .I2(n37_adj_5172), 
            .I3(GND_net), .O(n60602));   // verilog/uart_rx.v(119[33:55])
    defparam i45702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47158_4_lut (.I0(n60602), .I1(n61883), .I2(n41_adj_5174), 
            .I3(n60286), .O(n62058));   // verilog/uart_rx.v(119[33:55])
    defparam i47158_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47159_3_lut (.I0(n62058), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n62059));   // verilog/uart_rx.v(119[33:55])
    defparam i47159_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47127_3_lut (.I0(n62059), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n62027));   // verilog/uart_rx.v(119[33:55])
    defparam i47127_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45708_3_lut (.I0(n62027), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam i45708_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n7719[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n7745[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n7771[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n7797[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n7823[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n7849[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n7875[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n7901[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2646_5 (.CI(n45912), .I0(n2365), .I1(n856), .CO(n45913));
    SB_LUT4 r_Clock_Count_1943_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n46249), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2646_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n45911), 
            .O(n7771[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1943_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n46248), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1943_add_4_8 (.CI(n46248), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n46249));
    SB_LUT4 r_Clock_Count_1943_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n46247), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_4 (.CI(n45911), .I0(n2366), .I1(n698), .CO(n45912));
    SB_CARRY r_Clock_Count_1943_add_4_7 (.CI(n46247), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n46248));
    SB_LUT4 i46757_3_lut (.I0(n8_adj_5171), .I1(baudrate[13]), .I2(n31_adj_5159), 
            .I3(GND_net), .O(n61657));   // verilog/uart_rx.v(119[33:55])
    defparam i46757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46758_3_lut (.I0(n61657), .I1(baudrate[14]), .I2(n33_adj_5185), 
            .I3(GND_net), .O(n61658));   // verilog/uart_rx.v(119[33:55])
    defparam i46758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1943_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n46246), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2646_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n45910), 
            .O(n7771[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1943_add_4_6 (.CI(n46246), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n46247));
    SB_CARRY add_2646_3 (.CI(n45910), .I0(n2367), .I1(n858), .CO(n45911));
    SB_LUT4 add_2646_2_lut (.I0(n53466), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55362)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 r_Clock_Count_1943_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n46245), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1943_add_4_5 (.CI(n46245), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n46246));
    SB_CARRY add_2646_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45910));
    SB_LUT4 add_2645_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n45909), 
            .O(n7745[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2645_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n45908), 
            .O(n7745[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_15 (.CI(n45908), .I0(n2228), .I1(n2397), .CO(n45909));
    SB_LUT4 add_2645_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n45907), 
            .O(n7745[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_14 (.CI(n45907), .I0(n2229), .I1(n2272), .CO(n45908));
    SB_LUT4 add_2645_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n45906), 
            .O(n7745[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1943_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n46244), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_13 (.CI(n45906), .I0(n2230), .I1(n2144), .CO(n45907));
    SB_LUT4 add_2645_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n45905), 
            .O(n7745[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_12 (.CI(n45905), .I0(n2231), .I1(n2013), .CO(n45906));
    SB_CARRY r_Clock_Count_1943_add_4_4 (.CI(n46244), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n46245));
    SB_LUT4 add_2645_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n45904), 
            .O(n7745[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1943_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n46243), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1943_add_4_3 (.CI(n46243), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n46244));
    SB_CARRY add_2645_11 (.CI(n45904), .I0(n2232), .I1(n1879), .CO(n45905));
    SB_LUT4 r_Clock_Count_1943_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1943_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2645_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n45903), 
            .O(n7745[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_10 (.CI(n45903), .I0(n2233), .I1(n1742), .CO(n45904));
    SB_LUT4 add_2645_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n45902), 
            .O(n7745[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1943_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n46243));
    SB_CARRY add_2645_9 (.CI(n45902), .I0(n2234), .I1(n1602), .CO(n45903));
    SB_LUT4 add_2645_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n45901), 
            .O(n7745[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_8 (.CI(n45901), .I0(n2235), .I1(n1459), .CO(n45902));
    SB_LUT4 add_2645_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n45900), 
            .O(n7745[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_7 (.CI(n45900), .I0(n2236), .I1(n1460), .CO(n45901));
    SB_LUT4 add_2645_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n45899), 
            .O(n7745[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_6 (.CI(n45899), .I0(n2237), .I1(n1011), .CO(n45900));
    SB_LUT4 add_2645_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n45898), 
            .O(n7745[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_5 (.CI(n45898), .I0(n2238), .I1(n856), .CO(n45899));
    SB_LUT4 add_2645_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n45897), 
            .O(n7745[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_4 (.CI(n45897), .I0(n2239), .I1(n698), .CO(n45898));
    SB_LUT4 add_2645_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n45896), 
            .O(n7745[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_3 (.CI(n45896), .I0(n2240), .I1(n858), .CO(n45897));
    SB_LUT4 add_2645_2_lut (.I0(n53470), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55360)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2645_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45896));
    SB_LUT4 add_2644_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n45895), 
            .O(n7719[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2644_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n45894), 
            .O(n7719[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_13 (.CI(n45894), .I0(n2099), .I1(n2272), .CO(n45895));
    SB_LUT4 add_2644_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n45893), 
            .O(n7719[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_12 (.CI(n45893), .I0(n2100), .I1(n2144), .CO(n45894));
    SB_LUT4 add_2644_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n45892), 
            .O(n7719[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_11 (.CI(n45892), .I0(n2101), .I1(n2013), .CO(n45893));
    SB_LUT4 add_2644_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n45891), 
            .O(n7719[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_10 (.CI(n45891), .I0(n2102), .I1(n1879), .CO(n45892));
    SB_LUT4 add_2644_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n45890), 
            .O(n7719[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41393_1_lut_2_lut (.I0(baudrate[17]), .I1(n22959), .I2(GND_net), 
            .I3(GND_net), .O(n53462));
    defparam i41393_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_CARRY add_2644_9 (.CI(n45890), .I0(n2103), .I1(n1742), .CO(n45891));
    SB_LUT4 add_2644_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n45889), 
            .O(n7719[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_8 (.CI(n45889), .I0(n2104), .I1(n1602), .CO(n45890));
    SB_LUT4 add_2644_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n45888), 
            .O(n7719[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5186), .I1(baudrate[17]), 
            .I2(n39_adj_5146), .I3(GND_net), .O(n34_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44810_4_lut (.I0(n37_adj_5188), .I1(n35_adj_5189), .I2(n33_adj_5185), 
            .I3(n59717), .O(n59710));
    defparam i44810_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2644_7 (.CI(n45888), .I0(n2105), .I1(n1459), .CO(n45889));
    SB_LUT4 add_2644_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n45887), 
            .O(n7719[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1055 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n38068), .O(n55628));
    defparam i1_4_lut_adj_1055.LUT_INIT = 16'h0100;
    SB_CARRY add_2644_6 (.CI(n45887), .I0(n2106), .I1(n1460), .CO(n45888));
    SB_LUT4 add_2644_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n45886), 
            .O(n7719[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_5 (.CI(n45886), .I0(n2107), .I1(n1011), .CO(n45887));
    SB_LUT4 add_2644_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n45885), 
            .O(n7719[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_4 (.CI(n45885), .I0(n2108), .I1(n856), .CO(n45886));
    SB_LUT4 add_2644_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n45884), 
            .O(n7719[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_3 (.CI(n45884), .I0(n2109), .I1(n698), .CO(n45885));
    SB_LUT4 add_2644_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n7719[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n45884));
    SB_LUT4 add_2643_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n45883), 
            .O(n7693[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47398_2_lut_4_lut (.I0(n62023), .I1(baudrate[13]), .I2(n2098), 
            .I3(n22947), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i47398_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n55628), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n55646));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'h0002;
    SB_LUT4 add_2643_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n45882), 
            .O(n7693[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_13 (.CI(n45882), .I0(n1967), .I1(n2144), .CO(n45883));
    SB_LUT4 add_2643_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n45881), 
            .O(n7693[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_12 (.CI(n45881), .I0(n1968), .I1(n2013), .CO(n45882));
    SB_LUT4 add_2643_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n45880), 
            .O(n7693[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_11 (.CI(n45880), .I0(n1969), .I1(n1879), .CO(n45881));
    SB_LUT4 add_2643_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n45879), 
            .O(n7693[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_10 (.CI(n45879), .I0(n1970), .I1(n1742), .CO(n45880));
    SB_LUT4 add_2643_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n45878), 
            .O(n7693[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_9 (.CI(n45878), .I0(n1971), .I1(n1602), .CO(n45879));
    SB_LUT4 add_2643_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n45877), 
            .O(n7693[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_8 (.CI(n45877), .I0(n1972), .I1(n1459), .CO(n45878));
    SB_LUT4 add_2643_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n45876), 
            .O(n7693[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_7 (.CI(n45876), .I0(n1973), .I1(n1460), .CO(n45877));
    SB_LUT4 add_2643_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n45875), 
            .O(n7693[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_6 (.CI(n45875), .I0(n1974), .I1(n1011), .CO(n45876));
    SB_LUT4 add_2643_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n45874), 
            .O(n7693[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_5 (.CI(n45874), .I0(n1975), .I1(n856), .CO(n45875));
    SB_LUT4 add_2643_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n45873), 
            .O(n7693[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_4 (.CI(n45873), .I0(n1976), .I1(n698), .CO(n45874));
    SB_LUT4 add_2643_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n45872), 
            .O(n7693[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_3 (.CI(n45872), .I0(n1977), .I1(n858), .CO(n45873));
    SB_LUT4 add_2643_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7693[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45872));
    SB_LUT4 add_2653_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n46058), 
            .O(n7953[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n46057), 
            .O(n7953[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2642_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n45871), 
            .O(n7667[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2642_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n45870), 
            .O(n7667[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_24 (.CI(n46057), .I0(n3152), .I1(n3082), .CO(n46058));
    SB_LUT4 add_2653_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n46056), 
            .O(n7953[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_23 (.CI(n46056), .I0(n3153), .I1(n3188), .CO(n46057));
    SB_LUT4 add_2653_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n46055), 
            .O(n7953[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_12 (.CI(n45870), .I0(n1832), .I1(n2013), .CO(n45871));
    SB_LUT4 add_2642_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n45869), 
            .O(n7667[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_22 (.CI(n46055), .I0(n3154), .I1(n3084), .CO(n46056));
    SB_LUT4 add_2653_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n46054), 
            .O(n7953[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_21 (.CI(n46054), .I0(n3155), .I1(n2977), .CO(n46055));
    SB_CARRY add_2642_11 (.CI(n45869), .I0(n1833), .I1(n1879), .CO(n45870));
    SB_LUT4 add_2642_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n45868), 
            .O(n7667[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_10 (.CI(n45868), .I0(n1834), .I1(n1742), .CO(n45869));
    SB_LUT4 add_2653_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n46053), 
            .O(n7953[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2642_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n45867), 
            .O(n7667[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_9 (.CI(n45867), .I0(n1835), .I1(n1602), .CO(n45868));
    SB_LUT4 add_2642_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n45866), 
            .O(n7667[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_8 (.CI(n45866), .I0(n1836), .I1(n1459), .CO(n45867));
    SB_CARRY add_2653_20 (.CI(n46053), .I0(n3156), .I1(n2867), .CO(n46054));
    SB_LUT4 add_2642_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n45865), 
            .O(n7667[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_7 (.CI(n45865), .I0(n1837), .I1(n1460), .CO(n45866));
    SB_LUT4 add_2653_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n46052), 
            .O(n7953[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2642_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n45864), 
            .O(n7667[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_6 (.CI(n45864), .I0(n1838), .I1(n1011), .CO(n45865));
    SB_CARRY add_2653_19 (.CI(n46052), .I0(n3157), .I1(n2754), .CO(n46053));
    SB_LUT4 i47088_4_lut (.I0(n34_adj_5187), .I1(n14_adj_5190), .I2(n39_adj_5146), 
            .I3(n59697), .O(n61988));   // verilog/uart_rx.v(119[33:55])
    defparam i47088_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2642_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n45863), 
            .O(n7667[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n46051), 
            .O(n7953[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_5 (.CI(n45863), .I0(n1839), .I1(n856), .CO(n45864));
    SB_LUT4 add_2642_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n45862), 
            .O(n7667[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_4 (.CI(n45862), .I0(n1840), .I1(n698), .CO(n45863));
    SB_LUT4 add_2642_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n45861), 
            .O(n7667[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_18 (.CI(n46051), .I0(n3158), .I1(n2638), .CO(n46052));
    SB_LUT4 add_2653_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n46050), 
            .O(n7953[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_3 (.CI(n45861), .I0(n1841), .I1(n858), .CO(n45862));
    SB_LUT4 add_2642_2_lut (.I0(n53479), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55358)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2653_17 (.CI(n46050), .I0(n3159), .I1(n2519), .CO(n46051));
    SB_CARRY add_2642_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45861));
    SB_LUT4 add_2641_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n45860), 
            .O(n7641[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n46049), 
            .O(n7953[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2641_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n45859), 
            .O(n7641[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_10 (.CI(n45859), .I0(n1694), .I1(n1879), .CO(n45860));
    SB_LUT4 add_2641_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n45858), 
            .O(n7641[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_9 (.CI(n45858), .I0(n1695), .I1(n1742), .CO(n45859));
    SB_CARRY add_2653_16 (.CI(n46049), .I0(n3160), .I1(n2397), .CO(n46050));
    SB_LUT4 add_2641_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n45857), 
            .O(n7641[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n46048), 
            .O(n7953[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_8 (.CI(n45857), .I0(n1696), .I1(n1602), .CO(n45858));
    SB_LUT4 add_2641_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n45856), 
            .O(n7641[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_15 (.CI(n46048), .I0(n3161), .I1(n2272), .CO(n46049));
    SB_CARRY add_2641_7 (.CI(n45856), .I0(n1697), .I1(n1459), .CO(n45857));
    SB_LUT4 add_2653_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n46047), 
            .O(n7953[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2641_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n45855), 
            .O(n7641[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_6 (.CI(n45855), .I0(n1698), .I1(n1460), .CO(n45856));
    SB_CARRY add_2653_14 (.CI(n46047), .I0(n3162), .I1(n2144), .CO(n46048));
    SB_LUT4 add_2641_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n45854), 
            .O(n7641[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_5 (.CI(n45854), .I0(n1699), .I1(n1011), .CO(n45855));
    SB_LUT4 add_2641_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n45853), 
            .O(n7641[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n46046), 
            .O(n7953[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_4 (.CI(n45853), .I0(n1700), .I1(n856), .CO(n45854));
    SB_CARRY add_2653_13 (.CI(n46046), .I0(n3163), .I1(n2013), .CO(n46047));
    SB_LUT4 add_2641_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n45852), 
            .O(n7641[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_3 (.CI(n45852), .I0(n1701), .I1(n698), .CO(n45853));
    SB_LUT4 add_2653_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n46045), 
            .O(n7953[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2641_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n7641[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n45852));
    SB_CARRY add_2653_12 (.CI(n46045), .I0(n3164), .I1(n1879), .CO(n46046));
    SB_LUT4 add_2640_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n45851), 
            .O(n7615[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2640_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n45850), 
            .O(n7615[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n46044), 
            .O(n7953[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_10 (.CI(n45850), .I0(n1553), .I1(n1742), .CO(n45851));
    SB_LUT4 add_2640_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n45849), 
            .O(n7615[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_11 (.CI(n46044), .I0(n3165), .I1(n1742), .CO(n46045));
    SB_CARRY add_2640_9 (.CI(n45849), .I0(n1554), .I1(n1602), .CO(n45850));
    SB_LUT4 add_2640_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n45848), 
            .O(n7615[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_8 (.CI(n45848), .I0(n1555), .I1(n1459), .CO(n45849));
    SB_LUT4 add_2640_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n45847), 
            .O(n7615[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n46043), 
            .O(n7953[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_10 (.CI(n46043), .I0(n3166), .I1(n1602), .CO(n46044));
    SB_LUT4 add_2653_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n46042), 
            .O(n7953[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_7 (.CI(n45847), .I0(n1556), .I1(n1460), .CO(n45848));
    SB_LUT4 add_2640_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n45846), 
            .O(n7615[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_6 (.CI(n45846), .I0(n1557), .I1(n1011), .CO(n45847));
    SB_LUT4 add_2640_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n45845), 
            .O(n7615[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_9 (.CI(n46042), .I0(n3167), .I1(n1459), .CO(n46043));
    SB_CARRY add_2640_5 (.CI(n45845), .I0(n1558), .I1(n856), .CO(n45846));
    SB_LUT4 add_2640_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n45844), 
            .O(n7615[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_4 (.CI(n45844), .I0(n1559), .I1(n698), .CO(n45845));
    SB_LUT4 add_2653_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n46041), 
            .O(n7953[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2640_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n45843), 
            .O(n7615[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_3 (.CI(n45843), .I0(n1560), .I1(n858), .CO(n45844));
    SB_CARRY add_2653_8 (.CI(n46041), .I0(n3168), .I1(n1460), .CO(n46042));
    SB_LUT4 i41672_4_lut (.I0(n56497), .I1(n56417), .I2(n56421), .I3(n56313), 
            .O(n56563));
    defparam i41672_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2640_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7615[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n45843));
    SB_LUT4 add_2653_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n46040), 
            .O(n7953[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2639_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n45842), 
            .O(n7589[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_7 (.CI(n46040), .I0(n3169), .I1(n1011), .CO(n46041));
    SB_LUT4 add_2639_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n45841), 
            .O(n7589[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n46039), 
            .O(n7953[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_9 (.CI(n45841), .I0(n1409), .I1(n1602), .CO(n45842));
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2639_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n45840), 
            .O(n7589[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2653_6 (.CI(n46039), .I0(n3170), .I1(n856), .CO(n46040));
    SB_CARRY add_2639_8 (.CI(n45840), .I0(n1410), .I1(n1459), .CO(n45841));
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4985));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n55896));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'heeee;
    SB_LUT4 i24478_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38066));
    defparam i24478_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5844_4_lut (.I0(n804), .I1(n38066), .I2(n19207), .I3(baudrate[2]), 
            .O(n19237));   // verilog/uart_rx.v(119[33:55])
    defparam i5844_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47395_2_lut_4_lut (.I0(n61672), .I1(baudrate[10]), .I2(n1693), 
            .I3(n22938), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i47395_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55802));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1058 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55834));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1058.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_3_lut_4_lut_adj_1059 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55722));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1059.LUT_INIT = 16'hffef;
    SB_LUT4 i1_3_lut_4_lut_adj_1060 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55770));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1060.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1061 (.I0(n55894), .I1(n56533), .I2(baudrate[0]), 
            .I3(n48_adj_5132), .O(n962));
    defparam i1_3_lut_4_lut_adj_1061.LUT_INIT = 16'h0010;
    SB_LUT4 i41613_1_lut (.I0(n56503), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53479));
    defparam i41613_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(n61862), .I1(baudrate[14]), .I2(n2227), 
            .I3(n55360), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i47466_2_lut_4_lut (.I0(n61862), .I1(baudrate[14]), .I2(n2227), 
            .I3(n56292), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i47466_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47487_2_lut_4_lut (.I0(n62149), .I1(baudrate[20]), .I2(n2938), 
            .I3(n56537), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i47487_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i41641_1_lut_2_lut (.I0(baudrate[8]), .I1(n56529), .I2(GND_net), 
            .I3(GND_net), .O(n53492));
    defparam i41641_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i41642_2_lut_3_lut (.I0(baudrate[8]), .I1(n56529), .I2(baudrate[7]), 
            .I3(GND_net), .O(n56533));
    defparam i41642_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47449_2_lut_3_lut (.I0(baudrate[8]), .I1(n56529), .I2(n48), 
            .I3(GND_net), .O(n294[16]));
    defparam i47449_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut_adj_1062 (.I0(n62149), .I1(baudrate[20]), .I2(n2938), 
            .I3(n55372), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1062.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44532_4_lut (.I0(n35_adj_5206), .I1(n33_adj_5205), .I2(n31_adj_5204), 
            .I3(n29_adj_5207), .O(n59432));
    defparam i44532_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5208), .I1(baudrate[9]), 
            .I2(n43_adj_5202), .I3(GND_net), .O(n40_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46767_3_lut (.I0(n28_adj_5210), .I1(baudrate[5]), .I2(n35_adj_5206), 
            .I3(GND_net), .O(n61667));   // verilog/uart_rx.v(119[33:55])
    defparam i46767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46768_3_lut (.I0(n61667), .I1(baudrate[6]), .I2(n37_adj_5201), 
            .I3(GND_net), .O(n61668));   // verilog/uart_rx.v(119[33:55])
    defparam i46768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44528_4_lut (.I0(n41_adj_5203), .I1(n39_adj_5200), .I2(n37_adj_5201), 
            .I3(n59432), .O(n59428));
    defparam i44528_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46765_4_lut (.I0(n40_adj_5209), .I1(n30_adj_5211), .I2(n43_adj_5202), 
            .I3(n59424), .O(n61665));   // verilog/uart_rx.v(119[33:55])
    defparam i46765_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46623_3_lut (.I0(n61668), .I1(baudrate[7]), .I2(n39_adj_5200), 
            .I3(GND_net), .O(n61523));   // verilog/uart_rx.v(119[33:55])
    defparam i46623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47137_4_lut (.I0(n61523), .I1(n61665), .I2(n43_adj_5202), 
            .I3(n59428), .O(n62037));   // verilog/uart_rx.v(119[33:55])
    defparam i47137_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47138_3_lut (.I0(n62037), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n62038));   // verilog/uart_rx.v(119[33:55])
    defparam i47138_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n7693[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n7719[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n7745[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n7771[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n7797[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n7823[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n7849[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n7875[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n7901[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n56106));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24518_rep_5_2_lut (.I0(n7615[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n53482));   // verilog/uart_rx.v(119[33:55])
    defparam i24518_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3930_2_lut_4_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam i3930_2_lut_4_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n53482), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i46775_3_lut (.I0(n32_adj_5216), .I1(baudrate[6]), .I2(n39_adj_5215), 
            .I3(GND_net), .O(n61675));   // verilog/uart_rx.v(119[33:55])
    defparam i46775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46776_3_lut (.I0(n61675), .I1(baudrate[7]), .I2(n41_adj_5214), 
            .I3(GND_net), .O(n61676));   // verilog/uart_rx.v(119[33:55])
    defparam i46776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45440_4_lut (.I0(n41_adj_5214), .I1(n39_adj_5215), .I2(n37_adj_5213), 
            .I3(n59457), .O(n60340));
    defparam i45440_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46309_3_lut (.I0(n34_adj_5217), .I1(baudrate[5]), .I2(n37_adj_5213), 
            .I3(GND_net), .O(n61209));   // verilog/uart_rx.v(119[33:55])
    defparam i46309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46619_3_lut (.I0(n61676), .I1(baudrate[8]), .I2(n43_adj_5212), 
            .I3(GND_net), .O(n61519));   // verilog/uart_rx.v(119[33:55])
    defparam i46619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(n56549), .I1(n56563), .I2(n53248), 
            .I3(n55646), .O(n53990));
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'h0100;
    SB_LUT4 i46771_4_lut (.I0(n61519), .I1(n61209), .I2(n43_adj_5212), 
            .I3(n60340), .O(n61671));   // verilog/uart_rx.v(119[33:55])
    defparam i46771_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46772_3_lut (.I0(n61671), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n61672));   // verilog/uart_rx.v(119[33:55])
    defparam i46772_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46621_3_lut (.I0(n61672), .I1(baudrate[10]), .I2(n1693), 
            .I3(GND_net), .O(n48_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam i46621_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1065 (.I0(n56148), .I1(n56104), .I2(n56106), 
            .I3(baudrate[11]), .O(n56134));
    defparam i1_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1066 (.I0(n56134), .I1(n56136), .I2(n56124), 
            .I3(n56080), .O(n22938));
    defparam i1_4_lut_adj_1066.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1067 (.I0(n62029), .I1(baudrate[15]), .I2(n2353), 
            .I3(n55362), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1067.LUT_INIT = 16'h7100;
    SB_LUT4 i1_3_lut_adj_1068 (.I0(n22938), .I1(n48_adj_5218), .I2(n538), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1068.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n7667[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n7693[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n7719[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n7745[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n7771[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n7797[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n7823[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1069 (.I0(n56156), .I1(n56152), .I2(n56154), 
            .I3(n56150), .O(n56136));
    defparam i1_4_lut_adj_1069.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n7849[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n7875[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46644_3_lut (.I0(n61658), .I1(baudrate[15]), .I2(n35_adj_5189), 
            .I3(GND_net), .O(n61544));   // verilog/uart_rx.v(119[33:55])
    defparam i46644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n7901[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47469_2_lut_4_lut (.I0(n62029), .I1(baudrate[15]), .I2(n2353), 
            .I3(n56290), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i47469_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n54622));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1070 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n54622), .O(n55482));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1070.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55482), .O(n55488));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'hfffe;
    SB_LUT4 i24486_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n53499));   // verilog/uart_rx.v(119[33:55])
    defparam i24486_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n53499), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i41562_2_lut (.I0(\o_Rx_DV_N_3464[12] ), .I1(n52133), .I2(GND_net), 
            .I3(GND_net), .O(n56453));
    defparam i41562_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41664_4_lut (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n56453), .O(n56555));
    defparam i41664_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n55488), .I1(r_SM_Main_2__N_3422[1]), 
            .I2(r_SM_Main_c[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n56555), 
            .I2(r_SM_Main_c[0]), .I3(n27), .O(n9643));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n9643), .I1(n2), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_2_lut_4_lut_adj_1072 (.I0(n61684), .I1(baudrate[6]), .I2(n1111), 
            .I3(n55352), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1072.LUT_INIT = 16'h7100;
    SB_LUT4 i46785_3_lut (.I0(n42_adj_5219), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n61685));   // verilog/uart_rx.v(119[33:55])
    defparam i46785_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46786_3_lut (.I0(n61685), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n61686));   // verilog/uart_rx.v(119[33:55])
    defparam i46786_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46605_3_lut (.I0(n61686), .I1(baudrate[5]), .I2(n53216), 
            .I3(GND_net), .O(n48_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam i46605_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47443_2_lut_4_lut (.I0(n61684), .I1(baudrate[6]), .I2(n1111), 
            .I3(n56533), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i47443_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1073 (.I0(n56094), .I1(n22971), .I2(n56136), 
            .I3(n56092), .O(n22990));
    defparam i1_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1074 (.I0(n22990), .I1(n48_adj_5220), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1074.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46779_3_lut (.I0(n32_adj_5225), .I1(baudrate[5]), .I2(n39_adj_5224), 
            .I3(GND_net), .O(n61679));   // verilog/uart_rx.v(119[33:55])
    defparam i46779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46780_3_lut (.I0(n61679), .I1(baudrate[6]), .I2(n41_adj_5223), 
            .I3(GND_net), .O(n61680));   // verilog/uart_rx.v(119[33:55])
    defparam i46780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45458_4_lut (.I0(n41_adj_5223), .I1(n39_adj_5224), .I2(n37_adj_5222), 
            .I3(n59476), .O(n60358));
    defparam i45458_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46307_3_lut (.I0(n34_adj_5226), .I1(baudrate[4]), .I2(n37_adj_5222), 
            .I3(GND_net), .O(n61207));   // verilog/uart_rx.v(119[33:55])
    defparam i46307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46615_3_lut (.I0(n61680), .I1(baudrate[7]), .I2(n43_adj_5221), 
            .I3(GND_net), .O(n61515));   // verilog/uart_rx.v(119[33:55])
    defparam i46615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7537[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46777_4_lut (.I0(n61515), .I1(n61207), .I2(n43_adj_5221), 
            .I3(n60358), .O(n61677));   // verilog/uart_rx.v(119[33:55])
    defparam i46777_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46778_3_lut (.I0(n61677), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n61678));   // verilog/uart_rx.v(119[33:55])
    defparam i46778_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46617_3_lut (.I0(n61678), .I1(baudrate[9]), .I2(n1552), .I3(GND_net), 
            .O(n48_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam i46617_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n7641[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n7667[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n7693[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n7719[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n7745[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41402_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), .I2(n22959), 
            .I3(GND_net), .O(n56290));
    defparam i41402_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n7771[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n7797[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1075 (.I0(n61532), .I1(baudrate[16]), .I2(n2476), 
            .I3(n55364), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1075.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n7823[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n7849[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7563[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47455_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n56503), .I3(n48_adj_5227), .O(n294[14]));
    defparam i47455_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i41638_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n56503), .I3(baudrate[9]), .O(n56529));
    defparam i41638_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n7875[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46759_3_lut (.I0(n10_adj_5228), .I1(baudrate[10]), .I2(n25_adj_5165), 
            .I3(GND_net), .O(n61659));   // verilog/uart_rx.v(119[33:55])
    defparam i46759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47473_2_lut_4_lut (.I0(n61532), .I1(baudrate[16]), .I2(n2476), 
            .I3(n56280), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i47473_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i46760_3_lut (.I0(n61659), .I1(baudrate[11]), .I2(n27_adj_5170), 
            .I3(GND_net), .O(n61660));   // verilog/uart_rx.v(119[33:55])
    defparam i46760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45692_4_lut (.I0(n27_adj_5170), .I1(n25_adj_5165), .I2(n23_adj_5166), 
            .I3(n59750), .O(n60592));
    defparam i45692_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n7901[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5229), .I1(baudrate[9]), 
            .I2(n23_adj_5166), .I3(GND_net), .O(n20_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46642_3_lut (.I0(n61660), .I1(baudrate[12]), .I2(n29_adj_5169), 
            .I3(GND_net), .O(n26_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam i46642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n55354), .I3(n48), .O(n34_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i41403_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n22959), .I3(GND_net), .O(n53466));
    defparam i41403_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1076 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n56094));
    defparam i1_2_lut_4_lut_adj_1076.LUT_INIT = 16'hfffe;
    SB_LUT4 i46781_3_lut (.I0(n34_adj_5232), .I1(baudrate[5]), .I2(n41_adj_5235), 
            .I3(GND_net), .O(n61681));   // verilog/uart_rx.v(119[33:55])
    defparam i46781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46782_3_lut (.I0(n61681), .I1(baudrate[6]), .I2(n43_adj_5236), 
            .I3(GND_net), .O(n61682));   // verilog/uart_rx.v(119[33:55])
    defparam i46782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45466_4_lut (.I0(n43_adj_5236), .I1(n41_adj_5235), .I2(n39_adj_5234), 
            .I3(n59496), .O(n60366));
    defparam i45466_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39_adj_5234), 
            .I3(GND_net), .O(n38_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46594_4_lut (.I0(n37_adj_5188), .I1(n35_adj_5189), .I2(n33_adj_5185), 
            .I3(n59725), .O(n61494));
    defparam i46594_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46613_3_lut (.I0(n61682), .I1(baudrate[7]), .I2(n45_adj_5233), 
            .I3(GND_net), .O(n44_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam i46613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46305_4_lut (.I0(n44_adj_5238), .I1(n38_adj_5237), .I2(n45_adj_5233), 
            .I3(n60366), .O(n61205));   // verilog/uart_rx.v(119[33:55])
    defparam i46305_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_adj_1077 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n56092));
    defparam i1_2_lut_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7615[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n7641[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n7667[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n7693[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n7719[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n7745[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n7771[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44524_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n59424));
    defparam i44524_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n7797[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n7823[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n7849[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1078 (.I0(n56082), .I1(n56503), .I2(n7615[14]), 
            .I3(n48_adj_5227), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1078.LUT_INIT = 16'h0010;
    SB_LUT4 i47234_4_lut (.I0(n61544), .I1(n61988), .I2(n39_adj_5146), 
            .I3(n59710), .O(n62134));   // verilog/uart_rx.v(119[33:55])
    defparam i47234_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n7875[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n7901[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47429_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n56533), .I3(n48_adj_5132), .O(n294[19]));
    defparam i47429_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i5815_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n19207));   // verilog/uart_rx.v(119[33:55])
    defparam i5815_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i41531_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n56421));
    defparam i41531_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7589[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7615[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n7641[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n7667[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(n55888), .I1(n55884), .I2(n55886), 
            .I3(n56313), .O(n55906));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'hfffe;
    SB_LUT4 i46319_4_lut (.I0(n26_adj_5231), .I1(n20_adj_5230), .I2(n29_adj_5169), 
            .I3(n60592), .O(n61219));   // verilog/uart_rx.v(119[33:55])
    defparam i46319_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n7693[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(n55896), .I1(n55892), .I2(n55894), 
            .I3(n55890), .O(n55908));
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n7719[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47254_4_lut (.I0(n61219), .I1(n62134), .I2(n39_adj_5146), 
            .I3(n61494), .O(n62154));   // verilog/uart_rx.v(119[33:55])
    defparam i47254_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n7745[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1081 (.I0(n55908), .I1(n22962), .I2(n55906), 
            .I3(GND_net), .O(n22983));
    defparam i1_3_lut_adj_1081.LUT_INIT = 16'hfefe;
    SB_LUT4 i47255_3_lut (.I0(n62154), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n62155));   // verilog/uart_rx.v(119[33:55])
    defparam i47255_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n7771[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47241_3_lut (.I0(n62155), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n62141));   // verilog/uart_rx.v(119[33:55])
    defparam i47241_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n7797[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46321_3_lut (.I0(n62141), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n61221));   // verilog/uart_rx.v(119[33:55])
    defparam i46321_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n7823[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n7849[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n7875[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n7901[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n53990), .I1(baudrate[2]), 
            .I2(n54410), .I3(GND_net), .O(n48_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7589[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7563[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41392_2_lut (.I0(baudrate[17]), .I1(n22959), .I2(GND_net), 
            .I3(GND_net), .O(n56280));
    defparam i41392_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7589[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7615[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n7641[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1082 (.I0(n55886), .I1(n56292), .I2(n7693[11]), 
            .I3(n48_adj_5184), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1082.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n7667[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41612_2_lut_3_lut (.I0(n55886), .I1(n56292), .I2(baudrate[12]), 
            .I3(GND_net), .O(n56503));
    defparam i41612_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n7693[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7615[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47332_2_lut (.I0(n48_adj_5129), .I1(n22983), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i47332_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n7719[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n7641[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47461_2_lut_3_lut (.I0(n55886), .I1(n56292), .I2(n48_adj_5184), 
            .I3(GND_net), .O(n294[11]));
    defparam i47461_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n7667[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n7745[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47386_2_lut (.I0(n48_adj_5130), .I1(n22999), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i47386_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n7771[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n7693[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n7797[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n7823[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n7849[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n7875[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n7901[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1083 (.I0(n56092), .I1(n56156), .I2(baudrate[16]), 
            .I3(n38066), .O(n55950));
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n7719[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45404_3_lut (.I0(n53990), .I1(n54410), .I2(baudrate[2]), 
            .I3(GND_net), .O(n59234));   // verilog/uart_rx.v(119[33:55])
    defparam i45404_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n7745[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n7771[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n7797[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1084 (.I0(n61221), .I1(baudrate[21]), .I2(n3046), 
            .I3(n55374), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1084.LUT_INIT = 16'h7100;
    SB_LUT4 i47490_2_lut_4_lut (.I0(n61221), .I1(baudrate[21]), .I2(n3046), 
            .I3(n22971), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i47490_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i45298_4_lut (.I0(n53248), .I1(n55950), .I2(n56094), .I3(n56024), 
            .O(n59235));   // verilog/uart_rx.v(119[33:55])
    defparam i45298_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_4_lut_adj_1085 (.I0(n61205), .I1(baudrate[8]), .I2(n1408), 
            .I3(n55356), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1085.LUT_INIT = 16'h7100;
    SB_LUT4 i47452_2_lut_4_lut (.I0(n61205), .I1(baudrate[8]), .I2(n1408), 
            .I3(n56529), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i47452_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i44596_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n59496));   // verilog/uart_rx.v(119[33:55])
    defparam i44596_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n7823[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n7849[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i427_4_lut (.I0(n59235), .I1(n59234), .I2(n294[21]), 
            .I3(n56280), .O(n53212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n7875[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4101_2_lut (.I0(n19287), .I1(n9427), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam i4101_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i44621_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n59521));   // verilog/uart_rx.v(119[33:55])
    defparam i44621_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5239), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i44576_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n59476));   // verilog/uart_rx.v(119[33:55])
    defparam i44576_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7537[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7589[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7615[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n7641[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n7667[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n7693[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n7719[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n7745[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n7771[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n7797[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n7823[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7563[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n7849[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n7875[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n7901[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n55886));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'heeee;
    SB_LUT4 i41639_1_lut (.I0(n56529), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53488));
    defparam i41639_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44557_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n59457));   // verilog/uart_rx.v(119[33:55])
    defparam i44557_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7589[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1087 (.I0(n62038), .I1(baudrate[11]), .I2(n1831), 
            .I3(n55358), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1087.LUT_INIT = 16'h7100;
    SB_LUT4 i47458_2_lut_4_lut (.I0(n62038), .I1(baudrate[11]), .I2(n1831), 
            .I3(n56503), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i47458_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7615[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44797_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n59697));
    defparam i44797_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i44608_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n59508));   // verilog/uart_rx.v(119[33:55])
    defparam i44608_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n7641[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n7667[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45384_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n60284));
    defparam i45384_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n56266));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n7693[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n7719[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n7745[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n7771[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i534_3_lut (.I0(n53212), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n53214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44850_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n59750));
    defparam i44850_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45333_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n60233));
    defparam i45333_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47389_2_lut (.I0(n48_adj_5220), .I1(n22990), .I2(GND_net), 
            .I3(GND_net), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i47389_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n7797[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1088 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n56028));
    defparam i1_2_lut_4_lut_adj_1088.LUT_INIT = 16'hfffe;
    SB_LUT4 i4108_2_lut_4_lut (.I0(n960), .I1(n9427), .I2(n19287), .I3(baudrate[3]), 
            .O(n44_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam i4108_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n7823[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1089 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3464[2] ), .I3(\o_Rx_DV_N_3464[1] ), .O(n56044));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_274_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3464[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5241));   // verilog/uart_rx.v(69[17:62])
    defparam equal_274_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4106_2_lut_3_lut (.I0(baudrate[3]), .I1(n19287), .I2(n9427), 
            .I3(GND_net), .O(n9434));   // verilog/uart_rx.v(119[33:55])
    defparam i4106_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(r_Clock_Count[3]), .I1(n3_adj_5241), 
            .I2(\o_Rx_DV_N_3464[4] ), .I3(n56044), .O(n56048));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'hffde;
    SB_LUT4 i4099_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9427));   // verilog/uart_rx.v(119[33:55])
    defparam i4099_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 equal_274_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3464[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_274_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44771_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5130), .I2(n22999), 
            .I3(GND_net), .O(n59671));   // verilog/uart_rx.v(119[33:55])
    defparam i44771_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3464[6] ), 
            .I3(n56048), .O(n56052));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'hffde;
    SB_LUT4 equal_274_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3464[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5242));   // verilog/uart_rx.v(69[17:62])
    defparam equal_274_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1092 (.I0(r_Clock_Count[6]), .I1(n8_adj_5242), 
            .I2(n56052), .I3(\o_Rx_DV_N_3464[7] ), .O(n52133));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1092.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_3_lut_4_lut_adj_1093 (.I0(n22983), .I1(n48_adj_5129), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44));
    defparam i1_3_lut_4_lut_adj_1093.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_1094 (.I0(n23), .I1(\o_Rx_DV_N_3464[12] ), .I2(n4855), 
            .I3(\o_Rx_DV_N_3464[8] ), .O(n55346));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1094.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1095 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n27), .I2(n29), 
            .I3(n55346), .O(r_SM_Main_2__N_3422[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1095.LUT_INIT = 16'hfffe;
    SB_LUT4 i45369_2_lut (.I0(n52133), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n59335));
    defparam i45369_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45366_4_lut (.I0(n59335), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3464[12] ), 
            .O(n59332));
    defparam i45366_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i44803_4_lut (.I0(n59332), .I1(r_SM_Main_c[0]), .I2(n27), 
            .I3(\o_Rx_DV_N_3464[24] ), .O(n59329));
    defparam i44803_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n7849[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47299_4_lut (.I0(\r_SM_Main[2] ), .I1(n59329), .I2(r_SM_Main_2__N_3422[1]), 
            .I3(r_SM_Main[1]), .O(n26549));
    defparam i47299_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(n52133), .I1(r_SM_Main[1]), .I2(r_Rx_Data), 
            .I3(r_SM_Main_c[0]), .O(n55440));
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3464[12] ), 
            .I3(n55440), .O(n55446));
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'h0100;
    SB_LUT4 i44767_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5129), .I2(n22983), 
            .I3(GND_net), .O(n59667));   // verilog/uart_rx.v(119[33:55])
    defparam i44767_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i47308_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3464[24] ), 
            .I2(n27), .I3(n55446), .O(n25247));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i47308_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i3944_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9263), .I3(n19237), 
            .O(n46_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam i3944_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i639_4_lut (.I0(n53214), .I1(n294[19]), .I2(n46_adj_5243), 
            .I3(baudrate[4]), .O(n53216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7589[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45331_2_lut_3_lut (.I0(n22983), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n59296));   // verilog/uart_rx.v(119[33:55])
    defparam i45331_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i41527_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n56417));
    defparam i41527_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1098 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n56164));
    defparam i1_2_lut_4_lut_adj_1098.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1099 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n56162));
    defparam i1_2_lut_4_lut_adj_1099.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7615[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n7641[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1100 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n56124));
    defparam i1_2_lut_4_lut_adj_1100.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1101 (.I0(n62017), .I1(baudrate[17]), .I2(n2596), 
            .I3(n55366), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1101.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45278_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n60178));
    defparam i45278_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45294_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n60194));
    defparam i45294_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47476_2_lut_4_lut (.I0(n62017), .I1(baudrate[17]), .I2(n2596), 
            .I3(n22959), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i47476_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45221_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n60121));
    defparam i45221_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45229_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n60129));
    defparam i45229_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n7667[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45145_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n60045));
    defparam i45145_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i47383_3_lut (.I0(n22983), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n22878));   // verilog/uart_rx.v(119[33:55])
    defparam i47383_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n7693[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45157_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n60057));
    defparam i45157_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45258_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48_adj_5220), 
            .I3(n22990), .O(n1115));
    defparam i45258_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i1_2_lut_4_lut_adj_1102 (.I0(n61975), .I1(baudrate[18]), .I2(n2713), 
            .I3(n55368), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1102.LUT_INIT = 16'h7100;
    SB_LUT4 i47479_2_lut_4_lut (.I0(n61975), .I1(baudrate[18]), .I2(n2713), 
            .I3(n22962), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i47479_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1103 (.I0(n62145), .I1(baudrate[19]), .I2(n2827), 
            .I3(n55370), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1103.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n7719[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n7745[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45108_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n60008));
    defparam i45108_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47497_2_lut_4_lut (.I0(n61912), .I1(baudrate[22]), .I2(n3151), 
            .I3(n22974), .O(n294[1]));
    defparam i47497_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47482_2_lut_4_lut (.I0(n62145), .I1(baudrate[19]), .I2(n2827), 
            .I3(n22965), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i47482_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i45112_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n60012));
    defparam i45112_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n7771[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1104 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55738));
    defparam i1_3_lut_4_lut_adj_1104.LUT_INIT = 16'hfff7;
    SB_LUT4 i44725_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n59625));
    defparam i44725_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n7797[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n7823[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n7849[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n7875[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1105 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55754));
    defparam i1_3_lut_4_lut_adj_1105.LUT_INIT = 16'hff7f;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7563[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1106 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55786));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1106.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1107 (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(n4_adj_5199), .O(n55818));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1107.LUT_INIT = 16'hfffb;
    SB_LUT4 i45204_4_lut (.I0(r_SM_Main_c[0]), .I1(\o_Rx_DV_N_3464[12] ), 
            .I2(n4855), .I3(\o_Rx_DV_N_3464[8] ), .O(n59223));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i45204_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i45307_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3464[12] ), .I2(n52133), 
            .I3(r_SM_Main_c[0]), .O(n59229));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i45307_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i45201_4_lut (.I0(n59223), .I1(\o_Rx_DV_N_3464[24] ), .I2(n29), 
            .I3(n23), .O(n59220));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i45201_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45209_4_lut (.I0(n59229), .I1(\o_Rx_DV_N_3464[24] ), .I2(n29), 
            .I3(n23), .O(n59226));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i45209_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n59226), .I1(n59220), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5154));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7589[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44761_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n59661));
    defparam i44761_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7615[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45060_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n59960));
    defparam i45060_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n7641[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9434), .I3(n19289), 
            .O(n46_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam i4115_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i742_4_lut (.I0(n53216), .I1(n294[18]), .I2(n46_adj_5244), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n7667[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n7693[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n56056));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main_c[0]), .I1(\o_Rx_DV_N_3464[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5245));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3464[12] ), .I2(n23), .I3(n4855), 
            .O(n15_adj_5246));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5246), .I1(\o_Rx_DV_N_3464[8] ), .I2(n14_adj_5245), 
            .I3(n52352), .O(n62842));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45034_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n59934));
    defparam i45034_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n7719[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7537[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7537[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n7745[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n7771[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n7797[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1109 (.I0(n56148), .I1(n56056), .I2(n55860), 
            .I3(baudrate[19]), .O(n55880));
    defparam i1_4_lut_adj_1109.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n7823[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n7849[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5240), .I1(baudrate[4]), 
            .I2(n41_adj_5198), .I3(GND_net), .O(n40_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n7875[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47084_4_lut (.I0(n40_adj_5248), .I1(n36_adj_5247), .I2(n41_adj_5198), 
            .I3(n59508), .O(n61984));   // verilog/uart_rx.v(119[33:55])
    defparam i47084_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n7875[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47085_3_lut (.I0(n61984), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n61985));   // verilog/uart_rx.v(119[33:55])
    defparam i47085_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44886_4_lut (.I0(n33_adj_5192), .I1(n21_adj_5193), .I2(n19_adj_5194), 
            .I3(n17_adj_5191), .O(n59786));
    defparam i44886_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45821_4_lut (.I0(n15_adj_5195), .I1(n13_adj_5197), .I2(n2956), 
            .I3(baudrate[2]), .O(n60721));
    defparam i45821_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_4_lut_adj_1110 (.I0(n55880), .I1(n56106), .I2(n56150), 
            .I3(n56108), .O(n22962));
    defparam i1_4_lut_adj_1110.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1111 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n55314));
    defparam i1_3_lut_4_lut_adj_1111.LUT_INIT = 16'hfffe;
    SB_LUT4 i41606_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n56497));
    defparam i41606_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5008));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44996_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n59896));
    defparam i44996_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5006));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38582_1_lut_4_lut (.I0(n56264), .I1(n56266), .I2(n56104), 
            .I3(n56262), .O(n53438));
    defparam i38582_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i44953_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n59853));
    defparam i44953_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1112 (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), 
            .I2(\r_SM_Main[2] ), .I3(GND_net), .O(n4_adj_5199));
    defparam i1_2_lut_3_lut_adj_1112.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_4_lut_adj_1113 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55722), .O(n55728));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1113.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1114 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55728), .O(n55734));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1114.LUT_INIT = 16'hfffe;
    SB_LUT4 i46968_3_lut (.I0(n61985), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n61868));   // verilog/uart_rx.v(119[33:55])
    defparam i46968_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46347_4_lut (.I0(n21_adj_5193), .I1(n19_adj_5194), .I2(n17_adj_5191), 
            .I3(n60721), .O(n61247));
    defparam i46347_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46343_4_lut (.I0(n27_adj_4985), .I1(n25), .I2(n23_adj_5196), 
            .I3(n61247), .O(n61243));
    defparam i46343_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i44890_4_lut (.I0(n33_adj_5192), .I1(n31_adj_5123), .I2(n29_adj_5088), 
            .I3(n61243), .O(n59790));
    defparam i44890_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46902_3_lut (.I0(n61868), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i46902_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7537[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46523_3_lut (.I0(n10_adj_5249), .I1(baudrate[13]), .I2(n33_adj_5192), 
            .I3(GND_net), .O(n61423));   // verilog/uart_rx.v(119[33:55])
    defparam i46523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38598_1_lut (.I0(n22962), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53454));
    defparam i38598_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46524_3_lut (.I0(n61423), .I1(baudrate[14]), .I2(n35_adj_5090), 
            .I3(GND_net), .O(n61424));   // verilog/uart_rx.v(119[33:55])
    defparam i46524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1115 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55834), .O(n55840));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1115.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1116 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55840), .O(n55846));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1116.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7563[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47423_4_lut_4_lut (.I0(r_SM_Main_2__N_3422[1]), .I1(r_SM_Main[1]), 
            .I2(n6), .I3(n54622), .O(n53350));
    defparam i47423_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55802), .O(n55808));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n29), .I2(n23), 
            .I3(n55808), .O(n55814));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1119 (.I0(n23), .I1(\o_Rx_DV_N_3464[12] ), .I2(n4858), 
            .I3(GND_net), .O(n55390));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_1119.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1120 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n27), .I2(n29), 
            .I3(n55390), .O(\r_SM_Main_2__N_3512[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1120.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1121 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n55316));
    defparam i1_3_lut_4_lut_adj_1121.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1122 (.I0(n23), .I1(\o_Rx_DV_N_3464[12] ), .I2(n4858), 
            .I3(\r_SM_Main[0]_adj_7 ), .O(n55422));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1122.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1123 (.I0(\o_Rx_DV_N_3464[24] ), .I1(n27), .I2(n29), 
            .I3(n55422), .O(n53934));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1123.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5134), .I1(baudrate[17]), 
            .I2(n41_adj_5122), .I3(GND_net), .O(n36_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44913_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n59813));
    defparam i44913_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i44881_4_lut (.I0(n39_adj_5089), .I1(n37), .I2(n35_adj_5090), 
            .I3(n59786), .O(n59781));
    defparam i44881_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47021_4_lut (.I0(n36_adj_5251), .I1(n16_adj_5120), .I2(n41_adj_5122), 
            .I3(n59776), .O(n61921));   // verilog/uart_rx.v(119[33:55])
    defparam i47021_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i41404_2_lut_4_lut (.I0(baudrate[15]), .I1(baudrate[16]), .I2(baudrate[17]), 
            .I3(n22959), .O(n56292));
    defparam i41404_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3935_2_lut_2_lut_4_lut (.I0(baudrate[2]), .I1(n805), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n9263));   // verilog/uart_rx.v(119[33:55])
    defparam i3935_2_lut_2_lut_4_lut.LUT_INIT = 16'h0445;
    SB_LUT4 i2153_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2153_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2146_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2146_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i41405_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[15]), .I1(baudrate[16]), 
            .I2(baudrate[17]), .I3(n22959), .O(n53470));
    defparam i41405_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1124 (.I0(\o_Rx_DV_N_3464[12] ), .I1(n4855), .I2(\o_Rx_DV_N_3464[8] ), 
            .I3(n55818), .O(n55824));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1124.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (\a_new[1] , b_prev, GND_net, ENCODER0_B_N_keep, 
            n1884, ENCODER0_A_N_keep, n1842, n1844, n1846, n1848, 
            n1850, n1852, n1854, n1856, \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            position_31__N_3803, \encoder0_position[18] , \encoder0_position[17] , 
            \encoder0_position[16] , \encoder0_position[15] , \encoder0_position[14] , 
            \encoder0_position[13] , \encoder0_position[12] , \encoder0_position[11] , 
            \encoder0_position[10] , \encoder0_position[9] , \encoder0_position[8] , 
            \encoder0_position[7] , \encoder0_position[6] , \encoder0_position[5] , 
            \encoder0_position[4] , \encoder0_position[3] , \encoder0_position[2] , 
            \encoder0_position[1] , n27057, n1840, \encoder0_position[0] , 
            VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    output b_prev;
    input GND_net;
    input ENCODER0_B_N_keep;
    input n1884;
    input ENCODER0_A_N_keep;
    output n1842;
    output n1844;
    output n1846;
    output n1848;
    output n1850;
    output n1852;
    output n1854;
    output n1856;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output position_31__N_3803;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    input n27057;
    output n1840;
    output \encoder0_position[0] ;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_3811, direction_N_3808;
    wire [31:0]n133;
    
    wire n46167, n46166, n46165, debounce_cnt, n46164, n46163, n46162, 
        n46161, n46160, n46159, n46158, n46157, n46156, n46155, 
        position_31__N_3806, a_prev, n46154, n46153, n46152, n46151, 
        n46150, n46149, n46148, n46147, n46146, n46145, n46144, 
        n46143, n46142, n46141, n46140, n46139, n46138, n46137, 
        n27059, n27058;
    
    SB_LUT4 i47313_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3811));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i47313_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3808));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1884), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1884), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1934_add_4_33_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1842), .I3(n46167), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1934_add_4_32_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1844), .I3(n46166), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_32 (.CI(n46166), .I0(direction_N_3808), 
            .I1(n1844), .CO(n46167));
    SB_LUT4 position_1934_add_4_31_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1846), .I3(n46165), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1884), .D(a_prev_N_3811));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1934_add_4_31 (.CI(n46165), .I0(direction_N_3808), 
            .I1(n1846), .CO(n46166));
    SB_LUT4 position_1934_add_4_30_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1848), .I3(n46164), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_30 (.CI(n46164), .I0(direction_N_3808), 
            .I1(n1848), .CO(n46165));
    SB_LUT4 position_1934_add_4_29_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1850), .I3(n46163), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_29 (.CI(n46163), .I0(direction_N_3808), 
            .I1(n1850), .CO(n46164));
    SB_LUT4 position_1934_add_4_28_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1852), .I3(n46162), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_28 (.CI(n46162), .I0(direction_N_3808), 
            .I1(n1852), .CO(n46163));
    SB_LUT4 position_1934_add_4_27_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1854), .I3(n46161), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_27 (.CI(n46161), .I0(direction_N_3808), 
            .I1(n1854), .CO(n46162));
    SB_LUT4 position_1934_add_4_26_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1856), .I3(n46160), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_26 (.CI(n46160), .I0(direction_N_3808), 
            .I1(n1856), .CO(n46161));
    SB_LUT4 position_1934_add_4_25_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[23] ), .I3(n46159), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_25 (.CI(n46159), .I0(direction_N_3808), 
            .I1(\encoder0_position[23] ), .CO(n46160));
    SB_LUT4 position_1934_add_4_24_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[22] ), .I3(n46158), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_24 (.CI(n46158), .I0(direction_N_3808), 
            .I1(\encoder0_position[22] ), .CO(n46159));
    SB_LUT4 position_1934_add_4_23_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[21] ), .I3(n46157), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_23 (.CI(n46157), .I0(direction_N_3808), 
            .I1(\encoder0_position[21] ), .CO(n46158));
    SB_LUT4 position_1934_add_4_22_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[20] ), .I3(n46156), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_22 (.CI(n46156), .I0(direction_N_3808), 
            .I1(\encoder0_position[20] ), .CO(n46157));
    SB_LUT4 position_1934_add_4_21_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[19] ), .I3(n46155), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3806));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3806), 
            .I3(\a_new[1] ), .O(position_31__N_3803));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_CARRY position_1934_add_4_21 (.CI(n46155), .I0(direction_N_3808), 
            .I1(\encoder0_position[19] ), .CO(n46156));
    SB_LUT4 position_1934_add_4_20_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[18] ), .I3(n46154), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_20 (.CI(n46154), .I0(direction_N_3808), 
            .I1(\encoder0_position[18] ), .CO(n46155));
    SB_LUT4 position_1934_add_4_19_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[17] ), .I3(n46153), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_19 (.CI(n46153), .I0(direction_N_3808), 
            .I1(\encoder0_position[17] ), .CO(n46154));
    SB_LUT4 position_1934_add_4_18_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[16] ), .I3(n46152), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_18 (.CI(n46152), .I0(direction_N_3808), 
            .I1(\encoder0_position[16] ), .CO(n46153));
    SB_LUT4 position_1934_add_4_17_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[15] ), .I3(n46151), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_17 (.CI(n46151), .I0(direction_N_3808), 
            .I1(\encoder0_position[15] ), .CO(n46152));
    SB_LUT4 position_1934_add_4_16_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[14] ), .I3(n46150), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_16 (.CI(n46150), .I0(direction_N_3808), 
            .I1(\encoder0_position[14] ), .CO(n46151));
    SB_LUT4 position_1934_add_4_15_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[13] ), .I3(n46149), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_15 (.CI(n46149), .I0(direction_N_3808), 
            .I1(\encoder0_position[13] ), .CO(n46150));
    SB_LUT4 position_1934_add_4_14_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[12] ), .I3(n46148), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_14 (.CI(n46148), .I0(direction_N_3808), 
            .I1(\encoder0_position[12] ), .CO(n46149));
    SB_LUT4 position_1934_add_4_13_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[11] ), .I3(n46147), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_13 (.CI(n46147), .I0(direction_N_3808), 
            .I1(\encoder0_position[11] ), .CO(n46148));
    SB_LUT4 position_1934_add_4_12_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[10] ), .I3(n46146), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_12 (.CI(n46146), .I0(direction_N_3808), 
            .I1(\encoder0_position[10] ), .CO(n46147));
    SB_LUT4 position_1934_add_4_11_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[9] ), .I3(n46145), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_11 (.CI(n46145), .I0(direction_N_3808), 
            .I1(\encoder0_position[9] ), .CO(n46146));
    SB_LUT4 position_1934_add_4_10_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[8] ), .I3(n46144), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_10 (.CI(n46144), .I0(direction_N_3808), 
            .I1(\encoder0_position[8] ), .CO(n46145));
    SB_LUT4 position_1934_add_4_9_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[7] ), .I3(n46143), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_9 (.CI(n46143), .I0(direction_N_3808), 
            .I1(\encoder0_position[7] ), .CO(n46144));
    SB_LUT4 position_1934_add_4_8_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[6] ), .I3(n46142), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_8 (.CI(n46142), .I0(direction_N_3808), 
            .I1(\encoder0_position[6] ), .CO(n46143));
    SB_LUT4 position_1934_add_4_7_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[5] ), .I3(n46141), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_7 (.CI(n46141), .I0(direction_N_3808), 
            .I1(\encoder0_position[5] ), .CO(n46142));
    SB_LUT4 position_1934_add_4_6_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[4] ), .I3(n46140), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_6 (.CI(n46140), .I0(direction_N_3808), 
            .I1(\encoder0_position[4] ), .CO(n46141));
    SB_LUT4 position_1934_add_4_5_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[3] ), .I3(n46139), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_5 (.CI(n46139), .I0(direction_N_3808), 
            .I1(\encoder0_position[3] ), .CO(n46140));
    SB_LUT4 position_1934_add_4_4_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[2] ), .I3(n46138), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_4 (.CI(n46138), .I0(direction_N_3808), 
            .I1(\encoder0_position[2] ), .CO(n46139));
    SB_LUT4 position_1934_add_4_3_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder0_position[1] ), .I3(n46137), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_3 (.CI(n46137), .I0(direction_N_3808), 
            .I1(\encoder0_position[1] ), .CO(n46138));
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1884), .D(n27059));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1884), .D(n27058));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1840), .C(n1884), .D(n27057));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1934_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1934_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1934_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n46137));
    SB_DFFE position_1934__i0 (.Q(\encoder0_position[0] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1884), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1884), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1934__i1 (.Q(\encoder0_position[1] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i2 (.Q(\encoder0_position[2] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i3 (.Q(\encoder0_position[3] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i4 (.Q(\encoder0_position[4] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i5 (.Q(\encoder0_position[5] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i6 (.Q(\encoder0_position[6] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i7 (.Q(\encoder0_position[7] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i8 (.Q(\encoder0_position[8] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i9 (.Q(\encoder0_position[9] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i10 (.Q(\encoder0_position[10] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i11 (.Q(\encoder0_position[11] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i12 (.Q(\encoder0_position[12] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i13 (.Q(\encoder0_position[13] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i14 (.Q(\encoder0_position[14] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i15 (.Q(\encoder0_position[15] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i16 (.Q(\encoder0_position[16] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i17 (.Q(\encoder0_position[17] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i18 (.Q(\encoder0_position[18] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i19 (.Q(\encoder0_position[19] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i20 (.Q(\encoder0_position[20] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i21 (.Q(\encoder0_position[21] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i22 (.Q(\encoder0_position[22] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i23 (.Q(\encoder0_position[23] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i24 (.Q(n1856), .C(n1884), .E(position_31__N_3803), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i25 (.Q(n1854), .C(n1884), .E(position_31__N_3803), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i26 (.Q(n1852), .C(n1884), .E(position_31__N_3803), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i27 (.Q(n1850), .C(n1884), .E(position_31__N_3803), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i28 (.Q(n1848), .C(n1884), .E(position_31__N_3803), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i29 (.Q(n1846), .C(n1884), .E(position_31__N_3803), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i30 (.Q(n1844), .C(n1884), .E(position_31__N_3803), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1934__i31 (.Q(n1842), .C(n1884), .E(position_31__N_3803), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 i13353_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3811), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n27059));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13352_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3811), .I2(b_new[1]), 
            .I3(b_prev), .O(n27058));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13352_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (clk_out, CS_c, CS_CLK_c, GND_net, n27237, \data[15] , 
            n27236, \data[12] , n27234, \data[11] , n27233, \data[10] , 
            n27232, \data[9] , n27231, \data[8] , n27230, \data[7] , 
            n27228, \data[6] , n27227, \data[5] , n27226, \data[4] , 
            n27224, \data[3] , n27223, \data[2] , n27222, \data[1] , 
            clk16MHz, \state[1] , \state[0] , n27584, \data[0] , n9, 
            n26934, n26932, \current[0] , n25021, \current[15] , n27462, 
            \current[1] , n27461, \current[2] , n27460, \current[3] , 
            n27459, \current[4] , n27458, \current[5] , n27457, \current[6] , 
            n27456, \current[7] , n27455, \current[8] , n27454, \current[9] , 
            n27453, \current[10] , n27452, \current[11] , VCC_net, 
            n15, n4, n22896, n22893, n4_adj_3, n22870, n22880, 
            state_7__N_4293, n6, n6_adj_4, n5, n6_adj_5, n5_adj_6, 
            n37991, n11) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output clk_out;
    output CS_c;
    output CS_CLK_c;
    input GND_net;
    input n27237;
    output \data[15] ;
    input n27236;
    output \data[12] ;
    input n27234;
    output \data[11] ;
    input n27233;
    output \data[10] ;
    input n27232;
    output \data[9] ;
    input n27231;
    output \data[8] ;
    input n27230;
    output \data[7] ;
    input n27228;
    output \data[6] ;
    input n27227;
    output \data[5] ;
    input n27226;
    output \data[4] ;
    input n27224;
    output \data[3] ;
    input n27223;
    output \data[2] ;
    input n27222;
    output \data[1] ;
    input clk16MHz;
    output \state[1] ;
    output \state[0] ;
    input n27584;
    output \data[0] ;
    input n9;
    input n26934;
    input n26932;
    output \current[0] ;
    output n25021;
    output \current[15] ;
    input n27462;
    output \current[1] ;
    input n27461;
    output \current[2] ;
    input n27460;
    output \current[3] ;
    input n27459;
    output \current[4] ;
    input n27458;
    output \current[5] ;
    input n27457;
    output \current[6] ;
    input n27456;
    output \current[7] ;
    input n27455;
    output \current[8] ;
    input n27454;
    output \current[9] ;
    input n27453;
    output \current[10] ;
    input n27452;
    output \current[11] ;
    input VCC_net;
    output n15;
    output n4;
    output n22896;
    output n22893;
    output n4_adj_3;
    output n22870;
    output n22880;
    output state_7__N_4293;
    output n6;
    output n6_adj_4;
    output n5;
    output n6_adj_5;
    output n5_adj_6;
    output n37991;
    output n11;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire clk_slow_N_4206, n26710;
    wire [7:0]n37;
    
    wire n25242;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n9649, n25026, n26186, n20075;
    wire [11:0]n1;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4288;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4207;
    wire [1:0]n1964;
    
    wire n38237;
    wire [7:0]n47;
    
    wire n46105, n46104, n46103, n46102, n46101, n46100, n46099, 
        n59201, n6637, n46242, n46241, n46240, n46239, n46238, 
        n46237, n46236, n46235, n46234, n46233, n46232, n46231, 
        n46230, n6_adj_4977, n6_adj_4978, n55099, n8, n7;
    
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n27237));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n27236));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n27234));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n27233));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n27232));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n27231));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n27230));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n27228));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n27227));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n27226));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n27224));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n27223));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n27222));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4206));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 i13004_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26710));   // verilog/tli4970.v(55[24:39])
    defparam i13004_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n27584));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_1931__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n25242), 
            .D(n37[7]), .R(n26710));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1931__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n25242), 
            .D(n37[6]), .R(n26710));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1931__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n25242), 
            .D(n37[5]), .R(n26710));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1931__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n25242), 
            .D(n37[4]), .R(n26710));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n25026), .D(n9649), 
            .R(n26186));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n26934));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n26932));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1931__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n25242), 
            .D(n20075));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1938_1939__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n1[0]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1940_1941__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n25021), 
            .D(n1964[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n27462));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n27461));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n27460));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n27459));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n27458));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n27457));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n27456));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n27455));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n27454));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n27453));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n27452));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n25026), .D(n38237), 
            .S(n26186));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1931__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n25242), 
            .D(n47[1]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1931__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n25242), 
            .D(n47[2]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1931__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n25242), 
            .D(n47[3]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1938_1939__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n1[1]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n1[2]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n1[3]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n1[4]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n1[5]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n1[6]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n1[7]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n1[8]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n1[9]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n1[10]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1938_1939__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n1[11]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1940_1941__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1940_1941__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 bit_counter_1931_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n46105), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1931_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n46104), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_8 (.CI(n46104), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n46105));
    SB_LUT4 bit_counter_1931_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n46103), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_7 (.CI(n46103), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n46104));
    SB_LUT4 bit_counter_1931_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n46102), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_6 (.CI(n46102), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n46103));
    SB_LUT4 bit_counter_1931_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n46101), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_5 (.CI(n46101), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n46102));
    SB_LUT4 bit_counter_1931_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n46100), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_4 (.CI(n46100), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n46101));
    SB_LUT4 bit_counter_1931_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n46099), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_3 (.CI(n46099), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n46100));
    SB_LUT4 bit_counter_1931_add_4_2_lut (.I0(n6637), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n59201)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1931_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 counter_1940_1941_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n46242), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1931_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n46099));
    SB_LUT4 counter_1940_1941_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n46241), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_3 (.CI(n46241), .I0(GND_net), .I1(counter[1]), 
            .CO(n46242));
    SB_LUT4 counter_1940_1941_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n46241));
    SB_LUT4 delay_counter_1938_1939_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n46240), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1938_1939_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n46239), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_12 (.CI(n46239), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n46240));
    SB_LUT4 delay_counter_1938_1939_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n46238), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_11 (.CI(n46238), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n46239));
    SB_LUT4 delay_counter_1938_1939_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n46237), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_10 (.CI(n46237), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n46238));
    SB_LUT4 delay_counter_1938_1939_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n46236), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_9 (.CI(n46236), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n46237));
    SB_LUT4 delay_counter_1938_1939_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n46235), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_8 (.CI(n46235), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n46236));
    SB_LUT4 delay_counter_1938_1939_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n46234), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_7 (.CI(n46234), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n46235));
    SB_LUT4 delay_counter_1938_1939_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n46233), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_6 (.CI(n46233), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n46234));
    SB_LUT4 delay_counter_1938_1939_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n46232), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_5 (.CI(n46232), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n46233));
    SB_LUT4 delay_counter_1938_1939_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n46231), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_4 (.CI(n46231), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n46232));
    SB_LUT4 delay_counter_1938_1939_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n46230), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_3 (.CI(n46230), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n46231));
    SB_LUT4 delay_counter_1938_1939_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1938_1939_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1938_1939_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n46230));
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4288), .O(n25026));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i12480_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4288), .O(n26186));
    defparam i12480_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_999 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_999.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1000 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n22896));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1000.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1001 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n22893));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1001.LUT_INIT = 16'hffbf;
    SB_LUT4 i2056_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4207));
    defparam i2056_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4207), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4206));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1895_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n6637));   // verilog/tli4970.v(35[10] 68[6])
    defparam i1895_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1002 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4_adj_3));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1002.LUT_INIT = 16'hfffb;
    SB_LUT4 i47329_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n38237));
    defparam i47329_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[1]), 
            .I3(bit_counter[0]), .O(n22870));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1003 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[1]), .I3(bit_counter[0]), .O(n22880));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1003.LUT_INIT = 16'hffbf;
    SB_LUT4 bit_counter_1931_mux_6_i4_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4293), .I3(n37[3]), .O(n47[3]));
    defparam bit_counter_1931_mux_6_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1931_mux_6_i3_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4293), .I3(n37[2]), .O(n47[2]));
    defparam bit_counter_1931_mux_6_i3_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1931_mux_6_i2_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(state_7__N_4293), .I3(n37[1]), .O(n47[1]));
    defparam bit_counter_1931_mux_6_i2_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 equal_342_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_342_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_340_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4));   // verilog/tli4970.v(54[9:26])
    defparam equal_340_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_340_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_340_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_335_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5));   // verilog/tli4970.v(54[9:26])
    defparam equal_335_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2112_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1964[0]));
    defparam i2112_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 equal_333_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_6));   // verilog/tli4970.v(54[9:26])
    defparam equal_333_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4293));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i24403_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n37991));
    defparam i24403_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6608_3_lut (.I0(\state[0] ), .I1(n59201), .I2(\state[1] ), 
            .I3(GND_net), .O(n20075));   // verilog/tli4970.v(55[24:39])
    defparam i6608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_271_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_271_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47293_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n25021));
    defparam i47293_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4977));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_4977), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(delay_counter[2]), .I1(delay_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4978));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1005 (.I0(delay_counter[3]), .I1(delay_counter[1]), 
            .I2(delay_counter[0]), .I3(n6_adj_4978), .O(n55099));
    defparam i4_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(delay_counter[10]), .I1(n55099), .I2(delay_counter[6]), 
            .I3(delay_counter[5]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(delay_counter[9]), .I1(n7), .I2(delay_counter[8]), 
            .I3(n8), .O(delay_counter_15__N_4288));
    defparam i5_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mux_2024_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n9649));
    defparam mux_2024_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i11622_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n25242));
    defparam i11622_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, clk16MHz, \state_7__N_3892[0] , enable_slow_N_4187, 
            data_ready, n26923, ID, n27501, n27500, n27499, n27498, 
            n27497, n27496, n27495, baudrate, n27486, n27485, n27484, 
            n27483, n27482, n27470, n27469, n27468, n27467, n27466, 
            n27465, n27464, n27463, n25014, n25295, n25293, \state[0] , 
            data, \state_7__N_4084[0] , n27252, n27251, sda_enable, 
            sda_out, \counter[0] , n37902, n6352, scl_enable, VCC_net, 
            n27572, n8, n27259, n27257, n27256, n27255, n27253, 
            n22915, scl, \state_7__N_4100[3] , n22875, n6, n22907, 
            n22918) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input \state_7__N_3892[0] ;
    output enable_slow_N_4187;
    output data_ready;
    input n26923;
    output [7:0]ID;
    input n27501;
    input n27500;
    input n27499;
    input n27498;
    input n27497;
    input n27496;
    input n27495;
    output [31:0]baudrate;
    input n27486;
    input n27485;
    input n27484;
    input n27483;
    input n27482;
    input n27470;
    input n27469;
    input n27468;
    input n27467;
    input n27466;
    input n27465;
    input n27464;
    input n27463;
    output n25014;
    output n25295;
    output n25293;
    output \state[0] ;
    output [7:0]data;
    output \state_7__N_4084[0] ;
    input n27252;
    input n27251;
    output sda_enable;
    output sda_out;
    output \counter[0] ;
    output n37902;
    output n6352;
    output scl_enable;
    input VCC_net;
    input n27572;
    input n8;
    input n27259;
    input n27257;
    input n27256;
    input n27255;
    input n27253;
    output n22915;
    output scl;
    input \state_7__N_4100[3] ;
    output n22875;
    output n6;
    output n22907;
    output n22918;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n7, n47599, n25298;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n26714, n27212;
    wire [7:0]state_adj_4971;   // verilog/eeprom.v(27[11:16])
    
    wire n22785, n4, n13, n59382, n51587, ready_prev;
    wire [0:0]n5717;
    
    wire enable;
    wire [15:0]delay_counter_15__N_3930;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    wire [15:0]n5004;
    
    wire n45814, n45813, n45812, n45811, n45810, n38352, n43795, 
        n6612, n45809, n6611, n45808, n6610, n45807, n6609, n45806, 
        n6608, n45805, n45804, n6606, n45803, n45802, rw, n56459, 
        n51707, n35443, n26931, n45801, n45800;
    wire [2:0]n17;
    
    wire n24964, n43799;
    wire [7:0]state_7__N_3859;
    
    wire n54822, n27494, n27493, n27492, n27491, n27490, n27489, 
        n27488, n27487, n27481, n27480, n27479, n27478, n27477, 
        n27476, n27475, n27474, n27473, n27472, n27471, n38297, 
        n50, n66, n9, n43805, n46963, n56329, n28, n26, n27, 
        n25, n47072, n74, n69, n59178, n59180, n4_adj_4970, n59404, 
        n38314;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n51989;
    
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR byte_counter_1937__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n25298), .D(n47599), .R(n26714));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i2 (.Q(state_adj_4971[2]), .C(clk16MHz), .D(n27212));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i33_4_lut (.I0(\state_7__N_3892[0] ), .I1(n22785), .I2(state_adj_4971[1]), 
            .I3(n4), .O(n13));
    defparam i33_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i32_4_lut (.I0(n13), .I1(n59382), .I2(state_adj_4971[0]), 
            .I3(state_adj_4971[2]), .O(n51587));
    defparam i32_4_lut.LUT_INIT = 16'hf0ca;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4187));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5717[0]), .R(state_adj_4971[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1086_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5004[1]), 
            .I3(n45814), .O(delay_counter_15__N_3930[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1086_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5004[1]), 
            .I3(n45813), .O(delay_counter_15__N_3930[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_16 (.CI(n45813), .I0(delay_counter[14]), .I1(n5004[1]), 
            .CO(n45814));
    SB_LUT4 add_1086_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5004[1]), 
            .I3(n45812), .O(delay_counter_15__N_3930[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_15 (.CI(n45812), .I0(delay_counter[13]), .I1(n5004[1]), 
            .CO(n45813));
    SB_LUT4 add_1086_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5004[1]), 
            .I3(n45811), .O(delay_counter_15__N_3930[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_14 (.CI(n45811), .I0(delay_counter[12]), .I1(n5004[1]), 
            .CO(n45812));
    SB_LUT4 add_1086_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5004[1]), 
            .I3(n45810), .O(delay_counter_15__N_3930[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n38352));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i9_2_lut (.I0(state_adj_4971[2]), .I1(n38352), .I2(GND_net), 
            .I3(GND_net), .O(n43795));
    defparam i9_2_lut.LUT_INIT = 16'h7777;
    SB_CARRY add_1086_13 (.CI(n45810), .I0(delay_counter[11]), .I1(n5004[1]), 
            .CO(n45811));
    SB_LUT4 add_1086_12_lut (.I0(n43795), .I1(delay_counter[10]), .I2(n5004[1]), 
            .I3(n45809), .O(n6612)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_12 (.CI(n45809), .I0(delay_counter[10]), .I1(n5004[1]), 
            .CO(n45810));
    SB_LUT4 add_1086_11_lut (.I0(n43795), .I1(delay_counter[9]), .I2(n5004[1]), 
            .I3(n45808), .O(n6611)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_11 (.CI(n45808), .I0(delay_counter[9]), .I1(n5004[1]), 
            .CO(n45809));
    SB_LUT4 add_1086_10_lut (.I0(n43795), .I1(delay_counter[8]), .I2(n5004[1]), 
            .I3(n45807), .O(n6610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_10 (.CI(n45807), .I0(delay_counter[8]), .I1(n5004[1]), 
            .CO(n45808));
    SB_LUT4 add_1086_9_lut (.I0(n43795), .I1(delay_counter[7]), .I2(n5004[1]), 
            .I3(n45806), .O(n6609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_9 (.CI(n45806), .I0(delay_counter[7]), .I1(n5004[1]), 
            .CO(n45807));
    SB_LUT4 add_1086_8_lut (.I0(n43795), .I1(delay_counter[6]), .I2(n5004[1]), 
            .I3(n45805), .O(n6608)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_8 (.CI(n45805), .I0(delay_counter[6]), .I1(n5004[1]), 
            .CO(n45806));
    SB_LUT4 add_1086_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5004[1]), 
            .I3(n45804), .O(delay_counter_15__N_3930[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_7 (.CI(n45804), .I0(delay_counter[5]), .I1(n5004[1]), 
            .CO(n45805));
    SB_LUT4 add_1086_6_lut (.I0(n43795), .I1(delay_counter[4]), .I2(n5004[1]), 
            .I3(n45803), .O(n6606)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1086_6 (.CI(n45803), .I0(delay_counter[4]), .I1(n5004[1]), 
            .CO(n45804));
    SB_LUT4 add_1086_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5004[1]), 
            .I3(n45802), .O(delay_counter_15__N_3930[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut_4_lut (.I0(rw), .I1(state_adj_4971[1]), .I2(state_adj_4971[0]), 
            .I3(n56459), .O(n51707));   // verilog/eeprom.v(27[11:16])
    defparam i11_4_lut_4_lut.LUT_INIT = 16'haace;
    SB_CARRY add_1086_5 (.CI(n45802), .I0(delay_counter[3]), .I1(n5004[1]), 
            .CO(n45803));
    SB_LUT4 i14_4_lut_4_lut (.I0(state_adj_4971[2]), .I1(n38352), .I2(n35443), 
            .I3(data_ready), .O(n26931));   // verilog/eeprom.v(27[11:16])
    defparam i14_4_lut_4_lut.LUT_INIT = 16'hfa08;
    SB_LUT4 add_1086_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5004[1]), 
            .I3(n45801), .O(delay_counter_15__N_3930[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_4 (.CI(n45801), .I0(delay_counter[2]), .I1(n5004[1]), 
            .CO(n45802));
    SB_LUT4 i47283_2_lut (.I0(n22785), .I1(enable_slow_N_4187), .I2(GND_net), 
            .I3(GND_net), .O(n5004[1]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i47283_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_1086_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5004[1]), 
            .I3(n45800), .O(delay_counter_15__N_3930[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_3 (.CI(n45800), .I0(delay_counter[1]), .I1(n5004[1]), 
            .CO(n45801));
    SB_LUT4 add_1086_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5004[1]), 
            .I3(GND_net), .O(delay_counter_15__N_3930[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1086_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1086_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5004[1]), 
            .CO(n45800));
    SB_DFF state_i0 (.Q(state_adj_4971[0]), .C(clk16MHz), .D(n51587));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_1937__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n25298), .D(n17[2]), .R(n26714));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1937__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n25298), .D(n17[1]), .R(n26714));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n24964), .D(delay_counter_15__N_3930[12]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n24964), .D(delay_counter_15__N_3930[13]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n24964), .D(delay_counter_15__N_3930[14]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n24964), .D(delay_counter_15__N_3930[15]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n51707));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n26931));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n26923));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(state_adj_4971[1]), .C(clk16MHz), .E(n54822), 
            .D(state_7__N_3859[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n27501));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n27500));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n27499));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n27498));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n27497));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n27496));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n27495));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n27494));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n27493));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n27492));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n27491));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n27490));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n27489));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n27488));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n27487));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n27486));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n27485));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n27484));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n27483));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n27482));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n27481));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n27480));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n27479));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n27478));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n27477));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n27476));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n27475));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n27474));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n27473));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n27472));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n27471));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n27470));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n27469));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n27468));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n27467));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n27466));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n27465));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n27464));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n27463));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n24964), 
            .D(delay_counter_15__N_3930[1]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n24964), 
            .D(delay_counter_15__N_3930[2]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n24964), 
            .D(delay_counter_15__N_3930[3]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n24964), 
            .D(n6606), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n24964), 
            .D(delay_counter_15__N_3930[5]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n24964), 
            .D(n6608), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n24964), 
            .D(n6609), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n24964), 
            .D(n6610), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n24964), 
            .D(n6611), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n24964), .D(n6612), .S(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n24964), 
            .D(delay_counter_15__N_3930[0]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n24964), .D(delay_counter_15__N_3930[11]), .R(n43799));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i31658_3_lut_4_lut (.I0(n38297), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i31658_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i30301_4_lut_4_lut (.I0(state_adj_4971[2]), .I1(n38352), .I2(state_adj_4971[1]), 
            .I3(state_adj_4971[0]), .O(state_7__N_3859[1]));   // verilog/eeprom.v(27[11:16])
    defparam i30301_4_lut_4_lut.LUT_INIT = 16'ha5f2;
    SB_LUT4 i15_4_lut_4_lut (.I0(state_adj_4971[2]), .I1(n38352), .I2(state_adj_4971[1]), 
            .I3(state_adj_4971[0]), .O(n43799));   // verilog/eeprom.v(27[11:16])
    defparam i15_4_lut_4_lut.LUT_INIT = 16'h0502;
    SB_LUT4 i1_2_lut_3_lut (.I0(state_adj_4971[1]), .I1(state_adj_4971[2]), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n50));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_986 (.I0(state_adj_4971[1]), .I1(state_adj_4971[2]), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n66));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut_adj_986.LUT_INIT = 16'h2020;
    SB_LUT4 i2_3_lut_4_lut (.I0(state_adj_4971[1]), .I1(state_adj_4971[2]), 
            .I2(byte_counter[0]), .I3(n9), .O(n25014));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state_adj_4971[1]), .I1(state_adj_4971[2]), 
            .I2(n43805), .I3(byte_counter[0]), .O(n25295));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i2_3_lut_4_lut_adj_987 (.I0(byte_counter[1]), .I1(n46963), .I2(byte_counter[2]), 
            .I3(n50), .O(n25293));
    defparam i2_3_lut_4_lut_adj_987.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_adj_988 (.I0(byte_counter[1]), .I1(n46963), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n9));
    defparam i1_2_lut_3_lut_adj_988.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_989 (.I0(\state[0] ), .I1(state[3]), 
            .I2(state[1]), .I3(state[2]), .O(n4));
    defparam i1_2_lut_3_lut_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i41439_2_lut_3_lut (.I0(\state[0] ), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n56329));
    defparam i41439_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13788_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[0]), .I3(baudrate[0]), 
            .O(n27494));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13788_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13781_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[7]), .I3(baudrate[7]), 
            .O(n27487));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13781_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13782_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[6]), .I3(baudrate[6]), 
            .O(n27488));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13782_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13783_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[5]), .I3(baudrate[5]), 
            .O(n27489));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13783_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_990 (.I0(enable_slow_N_4187), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n47599));
    defparam i1_2_lut_3_lut_adj_990.LUT_INIT = 16'hd2d2;
    SB_LUT4 i1_4_lut_4_lut (.I0(state_adj_4971[2]), .I1(state_adj_4971[1]), 
            .I2(\state_7__N_3892[0] ), .I3(state_adj_4971[0]), .O(n25298));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h4410;
    SB_LUT4 i13784_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[4]), .I3(baudrate[4]), 
            .O(n27490));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13784_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_4_lut_adj_991 (.I0(state_adj_4971[2]), .I1(state_adj_4971[1]), 
            .I2(\state_7__N_3892[0] ), .I3(state_adj_4971[0]), .O(n26714));   // verilog/eeprom.v(68[25:39])
    defparam i1_4_lut_4_lut_adj_991.LUT_INIT = 16'h0010;
    SB_LUT4 i13785_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[3]), .I3(baudrate[3]), 
            .O(n27491));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13785_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13786_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[2]), .I3(baudrate[2]), 
            .O(n27492));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13786_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13787_3_lut_4_lut (.I0(n9), .I1(n66), .I2(data[1]), .I3(baudrate[1]), 
            .O(n27493));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13787_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n22785));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n22785), .I1(state_adj_4971[0]), .I2(enable_slow_N_4187), 
            .I3(GND_net), .O(n47072));
    defparam i2_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_992 (.I0(byte_counter[0]), .I1(n43805), 
            .I2(state_adj_4971[2]), .I3(state_adj_4971[1]), .O(n74));   // verilog/eeprom.v(68[25:39])
    defparam i1_2_lut_3_lut_4_lut_adj_992.LUT_INIT = 16'hfbff;
    SB_LUT4 mux_1437_Mux_0_i3_3_lut_4_lut (.I0(state_adj_4971[0]), .I1(n22785), 
            .I2(enable_slow_N_4187), .I3(state_adj_4971[1]), .O(n5717[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1437_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h10aa;
    SB_LUT4 i30246_4_lut (.I0(data[7]), .I1(n74), .I2(baudrate[15]), .I3(n25295), 
            .O(n27479));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i30246_4_lut.LUT_INIT = 16'heae0;
    SB_LUT4 i30269_4_lut (.I0(data[6]), .I1(n74), .I2(baudrate[14]), .I3(n25295), 
            .O(n27480));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i30269_4_lut.LUT_INIT = 16'heae0;
    SB_LUT4 i1_2_lut (.I0(state_adj_4971[2]), .I1(state_adj_4971[1]), .I2(GND_net), 
            .I3(GND_net), .O(n69));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i45009_4_lut (.I0(byte_counter[0]), .I1(n69), .I2(data[5]), 
            .I3(n43805), .O(n59178));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i45009_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i45179_2_lut (.I0(n43805), .I1(data[5]), .I2(GND_net), .I3(GND_net), 
            .O(n59180));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i45179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30259_4_lut (.I0(n59180), .I1(n59178), .I2(baudrate[13]), 
            .I3(n50), .O(n27481));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i30259_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i2_3_lut_adj_993 (.I0(byte_counter[2]), .I1(n46963), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n43805));
    defparam i2_3_lut_adj_993.LUT_INIT = 16'h4040;
    SB_LUT4 i13772_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[0]), .I3(baudrate[16]), 
            .O(n27478));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13772_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13765_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[7]), .I3(baudrate[23]), 
            .O(n27471));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13765_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13766_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[6]), .I3(baudrate[22]), 
            .O(n27472));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13766_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13767_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[5]), .I3(baudrate[21]), 
            .O(n27473));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13767_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13768_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[4]), .I3(baudrate[20]), 
            .O(n27474));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13769_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[3]), .I3(baudrate[19]), 
            .O(n27475));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13769_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13770_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[2]), .I3(baudrate[18]), 
            .O(n27476));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13771_3_lut_4_lut (.I0(n43805), .I1(n66), .I2(data[1]), .I3(baudrate[17]), 
            .O(n27477));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i31651_2_lut_3_lut_4_lut (.I0(enable_slow_N_4187), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i31651_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i1_4_lut (.I0(state_adj_4971[2]), .I1(state_adj_4971[0]), .I2(state_adj_4971[1]), 
            .I3(n38297), .O(n27212));
    defparam i1_4_lut.LUT_INIT = 16'ha8e8;
    SB_LUT4 i1_2_lut_adj_994 (.I0(state_adj_4971[0]), .I1(state_adj_4971[1]), 
            .I2(GND_net), .I3(GND_net), .O(n35443));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_995 (.I0(state_adj_4971[2]), .I1(state_adj_4971[1]), 
            .I2(\state_7__N_3892[0] ), .I3(state_adj_4971[0]), .O(n4_adj_4970));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'hbbba;
    SB_LUT4 i45379_4_lut (.I0(n56329), .I1(n22785), .I2(state_adj_4971[1]), 
            .I3(state[3]), .O(n59404));
    defparam i45379_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n59404), .I1(n4_adj_4970), .I2(n38297), .I3(state_adj_4971[0]), 
            .O(n54822));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i2_3_lut_4_lut_adj_996 (.I0(\state[0] ), .I1(state[3]), .I2(state[2]), 
            .I3(state[1]), .O(n38314));
    defparam i2_3_lut_4_lut_adj_996.LUT_INIT = 16'hfffe;
    SB_LUT4 i45330_2_lut_3_lut (.I0(enable_slow_N_4187), .I1(ready_prev), 
            .I2(state_adj_4971[1]), .I3(GND_net), .O(n59382));
    defparam i45330_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i2_3_lut_adj_997 (.I0(state_adj_4971[0]), .I1(ready_prev), .I2(n38314), 
            .I3(GND_net), .O(n46963));
    defparam i2_3_lut_adj_997.LUT_INIT = 16'h0202;
    SB_LUT4 i41568_3_lut (.I0(state_adj_4971[2]), .I1(n47072), .I2(state_adj_4971[1]), 
            .I3(GND_net), .O(n56459));
    defparam i41568_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_998 (.I0(n38314), .I1(saved_addr[0]), .I2(rw), 
            .I3(\state_7__N_4084[0] ), .O(n51989));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_998.LUT_INIT = 16'hd8cc;
    SB_LUT4 i47302_4_lut (.I0(state_adj_4971[0]), .I1(n38352), .I2(state_adj_4971[1]), 
            .I3(state_adj_4971[2]), .O(n24964));
    defparam i47302_4_lut.LUT_INIT = 16'h015a;
    i2c_controller i2c (.n27252(n27252), .data({data}), .n27251(n27251), 
            .sda_enable(sda_enable), .sda_out(sda_out), .GND_net(GND_net), 
            .clk16MHz(clk16MHz), .\counter[0] (\counter[0] ), .\state[2] (state[2]), 
            .\state[3] (state[3]), .n37902(n37902), .n6352(n6352), .\state_7__N_4084[0] (\state_7__N_4084[0] ), 
            .enable_slow_N_4187(enable_slow_N_4187), .scl_enable(scl_enable), 
            .VCC_net(VCC_net), .n27572(n27572), .n8(n8), .\state[0] (\state[0] ), 
            .n51989(n51989), .\saved_addr[0] (saved_addr[0]), .\state[1] (state[1]), 
            .n27259(n27259), .n27257(n27257), .n27256(n27256), .n27255(n27255), 
            .n27253(n27253), .n22915(n22915), .scl(scl), .\state_7__N_4100[3] (\state_7__N_4100[3] ), 
            .enable(enable), .n7(n7), .n22875(n22875), .ready_prev(ready_prev), 
            .n38297(n38297), .n6(n6), .n22907(n22907), .n22918(n22918)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n27252, data, n27251, sda_enable, sda_out, 
            GND_net, clk16MHz, \counter[0] , \state[2] , \state[3] , 
            n37902, n6352, \state_7__N_4084[0] , enable_slow_N_4187, 
            scl_enable, VCC_net, n27572, n8, \state[0] , n51989, 
            \saved_addr[0] , \state[1] , n27259, n27257, n27256, n27255, 
            n27253, n22915, scl, \state_7__N_4100[3] , enable, n7, 
            n22875, ready_prev, n38297, n6, n22907, n22918) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input n27252;
    output [7:0]data;
    input n27251;
    output sda_enable;
    output sda_out;
    input GND_net;
    input clk16MHz;
    output \counter[0] ;
    output \state[2] ;
    output \state[3] ;
    output n37902;
    output n6352;
    output \state_7__N_4084[0] ;
    output enable_slow_N_4187;
    output scl_enable;
    input VCC_net;
    input n27572;
    input n8;
    output \state[0] ;
    input n51989;
    output \saved_addr[0] ;
    output \state[1] ;
    input n27259;
    input n27257;
    input n27256;
    input n27255;
    input n27253;
    output n22915;
    output scl;
    input \state_7__N_4100[3] ;
    input enable;
    input n7;
    output n22875;
    input ready_prev;
    output n38297;
    output n6;
    output n22907;
    output n22918;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire sda_out_adj_4959;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n26560;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n12, n10, n6345, n10_adj_4960, n24935, n11, enable_slow_N_4186, 
        n10_adj_4961, i2c_clk_N_4173, scl_enable_N_4174;
    wire [7:0]n119;
    
    wire n45821, n45820, n45819, n45818, n25072, n45817, n45816, 
        n45815, n46262, n46261, n46260, n46259, n46258, n54417, 
        n25066, n51725, n54305, n25064, n25057, n26413, n5, n38175, 
        n38180, n38375, n55145, n54742, n9, n11_adj_4962, n15, 
        n11_adj_4963;
    wire [1:0]n6416;
    
    wire n6683, n11_adj_4964, n4, n15_adj_4965, n4_adj_4966, n59402, 
        n28, n62178, n53288;
    
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n27252));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n27251));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2417_2_lut (.I0(sda_out_adj_4959), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2417_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter2_1946_1947__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(\counter[0] ), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6345));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_280_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4960));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_280_i10_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i47291_4_lut (.I0(n24935), .I1(n6345), .I2(n11), .I3(n37902), 
            .O(n6352));
    defparam i47291_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i47320_2_lut (.I0(\state_7__N_4084[0] ), .I1(enable_slow_N_4187), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4186));   // verilog/i2c_controller.v(62[6:32])
    defparam i47320_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[4]), .I2(counter2[2]), 
            .I3(counter2[5]), .O(n10_adj_4961));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4961), .I2(counter2[0]), 
            .I3(GND_net), .O(n26560));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4173));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4174));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n45821), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n45820), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n45820), .I0(counter[6]), .I1(VCC_net), 
            .CO(n45821));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n45819), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n45819), .I0(counter[5]), .I1(VCC_net), 
            .CO(n45820));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n45818), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4084[0] ), .C(clk16MHz), .E(n25072), 
            .D(enable_slow_N_4186));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_CARRY sub_39_add_2_6 (.CI(n45818), .I0(counter[4]), .I1(VCC_net), 
            .CO(n45819));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n45817), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n45817), .I0(counter[3]), .I1(VCC_net), 
            .CO(n45818));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n45816), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n45816), .I0(counter[2]), .I1(VCC_net), 
            .CO(n45817));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n45815), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n45815), .I0(counter[1]), .I1(VCC_net), 
            .CO(n45816));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(\counter[0] ), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(\counter[0] ), .I1(GND_net), 
            .CO(n45815));
    SB_LUT4 counter2_1946_1947_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n46262), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n27572));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_1946_1947_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n46261), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1946_1947_add_4_6 (.CI(n46261), .I0(GND_net), .I1(counter2[4]), 
            .CO(n46262));
    SB_LUT4 counter2_1946_1947_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n46260), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1946_1947_add_4_5 (.CI(n46260), .I0(GND_net), .I1(counter2[3]), 
            .CO(n46261));
    SB_LUT4 counter2_1946_1947_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n46259), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1946_1947_add_4_4 (.CI(n46259), .I0(GND_net), .I1(counter2[2]), 
            .CO(n46260));
    SB_LUT4 counter2_1946_1947_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n46258), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1946_1947_add_4_3 (.CI(n46258), .I0(GND_net), .I1(counter2[1]), 
            .CO(n46259));
    SB_LUT4 counter2_1946_1947_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1946_1947_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1946_1947_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n46258));
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n51989));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n25066), 
            .D(n54417), .S(n51725));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4959), .C(i2c_clk), .E(n25064), 
            .D(n54305), .S(n51725));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(\counter[0] ), .C(i2c_clk), .E(n25057), .D(n119[0]), 
            .S(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n25057), .D(n119[1]), 
            .S(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n25057), .D(n119[2]), 
            .S(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n25057), .D(n119[3]), 
            .R(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n25057), .D(n119[4]), 
            .R(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n25057), .D(n119[5]), 
            .R(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n25057), .D(n119[6]), 
            .R(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n25057), .D(n119[7]), 
            .R(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6352), .D(n5), 
            .S(n38175));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6352), .D(n38180), 
            .S(n38375));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6352), .D(n55145), 
            .S(n54742));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1946_1947__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1946_1947__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1946_1947__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1946_1947__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1946_1947__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n26560));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n27259));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n27257));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n27256));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n27255));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n27253));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_279_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_279_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n26560), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4173));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4962));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut (.I0(counter[1]), .I1(counter[2]), .I2(n15), .I3(GND_net), 
            .O(n22915));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i2_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i47339_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(enable_slow_N_4187));   // verilog/i2c_controller.v(44[32:47])
    defparam i47339_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n11));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4963));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6416[1]), 
            .I3(\state[1] ), .O(n54305));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i2_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6683));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i24367_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i24367_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n54417));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'h1110;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4100[3] ), .I1(n11_adj_4963), .I2(n11_adj_4964), 
            .I3(enable), .O(n4));
    defparam i1_4_lut.LUT_INIT = 16'h2a2f;
    SB_LUT4 i47416_2_lut (.I0(\state_7__N_4100[3] ), .I1(n11_adj_4963), 
            .I2(GND_net), .I3(GND_net), .O(n38180));
    defparam i47416_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i12712_2_lut_4_lut (.I0(n25057), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n26413));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12712_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i47411_4_lut (.I0(n6352), .I1(\state[0] ), .I2(n11), .I3(n7), 
            .O(n38175));
    defparam i47411_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i1_4_lut_adj_976 (.I0(n11_adj_4962), .I1(n11_adj_4963), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4100[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_976.LUT_INIT = 16'h5575;
    SB_LUT4 equal_279_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15_adj_4965));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam equal_279_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_977 (.I0(\state[3] ), .I1(n6345), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4966));
    defparam i1_2_lut_adj_977.LUT_INIT = 16'hbbbb;
    SB_LUT4 i45376_4_lut (.I0(n7), .I1(n4_adj_4966), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n59402));
    defparam i45376_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n59402), .I1(n15_adj_4965), .I2(n6683), .I3(\state_7__N_4100[3] ), 
            .O(n25057));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i1_4_lut_adj_978 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut_adj_978.LUT_INIT = 16'h5110;
    SB_LUT4 i47278_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n62178));
    defparam i47278_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_979 (.I0(n11_adj_4964), .I1(n62178), .I2(n28), 
            .I3(n53288), .O(n25064));
    defparam i1_4_lut_adj_979.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1721_Mux_1_i7_4_lut (.I0(counter[1]), .I1(\counter[0] ), 
            .I2(counter[2]), .I3(\saved_addr[0] ), .O(n6416[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1721_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i38439_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n53288));
    defparam i38439_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n7), .I2(\state[3] ), .I3(n11_adj_4964), 
            .O(n51725));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_980 (.I0(n11_adj_4964), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n53288), .O(n25066));
    defparam i1_4_lut_adj_980.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_2_lut_3_lut (.I0(n15), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(n22875));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24707_2_lut (.I0(enable_slow_N_4187), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n38297));
    defparam i24707_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i47408_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6352), 
            .I3(\state[1] ), .O(n54742));   // verilog/i2c_controller.v(130[5:15])
    defparam i47408_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n15));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 equal_1504_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4964));   // verilog/i2c_controller.v(130[5:15])
    defparam equal_1504_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i24609_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n37902));   // verilog/i2c_controller.v(130[5:15])
    defparam i24609_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n24935));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i47410_3_lut_4_lut (.I0(n9), .I1(n10_adj_4960), .I2(n15), 
            .I3(n6352), .O(n38375));   // verilog/i2c_controller.v(139[9:14])
    defparam i47410_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i2_2_lut_3_lut_adj_981 (.I0(n9), .I1(n10_adj_4960), .I2(n11), 
            .I3(GND_net), .O(n6));   // verilog/i2c_controller.v(139[9:14])
    defparam i2_2_lut_3_lut_adj_981.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(\state[0] ), .I1(\state[1] ), .I2(n10_adj_4960), 
            .I3(n4), .O(n55145));   // verilog/i2c_controller.v(109[5:12])
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'hff04;
    SB_LUT4 i1_2_lut_3_lut_adj_983 (.I0(enable), .I1(\state_7__N_4084[0] ), 
            .I2(enable_slow_N_4187), .I3(GND_net), .O(n25072));
    defparam i1_2_lut_3_lut_adj_983.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_3_lut_adj_984 (.I0(n15), .I1(counter[1]), .I2(counter[2]), 
            .I3(GND_net), .O(n22907));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_3_lut_adj_984.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_adj_985 (.I0(n15), .I1(counter[1]), .I2(counter[2]), 
            .I3(GND_net), .O(n22918));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_3_lut_adj_985.LUT_INIT = 16'hfbfb;
    SB_LUT4 i24387_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(scl_enable_N_4174));   // verilog/i2c_controller.v(44[32:47])
    defparam i24387_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[3] , GND_net, \Ki[15] , \PID_CONTROLLER.integral_23__N_3691[7] , 
            \Kp[5] , \Kp[4] , PWMLimit, \Kp[0] , \Kp[1] , control_update, 
            duty, clk16MHz, reset, setpoint, \motor_state[18] , n35, 
            \Kp[6] , n181, IntegralLimit, n155, \Ki[6] , \PID_CONTROLLER.integral_23__N_3691[12] , 
            \Ki[1] , \PID_CONTROLLER.integral_23__N_3691[6] , \Ki[0] , 
            \Kp[2] , \Ki[7] , \Kp[12] , \Kp[7] , \Ki[2] , n11, \Ki[3] , 
            \Ki[8] , \Kp[13] , \Ki[14] , \PID_CONTROLLER.integral_23__N_3691[15] , 
            \PID_CONTROLLER.integral_23__N_3691[14] , n375, \PID_CONTROLLER.integral_23__N_3691[3] , 
            \Ki[9] , \Ki[4] , n214, \PID_CONTROLLER.integral_23__N_3691[16] , 
            \PID_CONTROLLER.integral_23__N_3691[4] , \Kp[8] , \PID_CONTROLLER.integral_23__N_3691[0] , 
            \Ki[12] , \Kp[14] , \Ki[5] , \Kp[15] , deadband, \motor_state[17] , 
            \PID_CONTROLLER.integral_23__N_3691[11] , \Ki[10] , n5, \motor_state[15] , 
            \motor_state[14] , n9, \Ki[11] , \motor_state[12] , n545, 
            n143, n220, \motor_state[11] , \motor_state[10] , VCC_net, 
            n472, \motor_state[9] , \motor_state[8] , \PID_CONTROLLER.integral_23__N_3691[10] , 
            n399, n326, n253, n180, \motor_state[7] , n53, \motor_state[6] , 
            n107, \motor_state[5] , n203, \motor_state[4] , n204, 
            \motor_state[3] , \motor_state[2] , \Kp[11] , \motor_state[1] , 
            \Kp[9] , \motor_state[0] , \PID_CONTROLLER.integral_23__N_3691[1] , 
            \Kp[10] , \PID_CONTROLLER.integral_23__N_3691[13] , \Ki[13] , 
            n26922, \PID_CONTROLLER.integral , n27524, n27523, n27522, 
            n27521, n27520, n27519, n27518, n27517, n27516, n27515, 
            n27514, n27513, n27512, n27511, n27510, n27509, n27508, 
            n27507, n27506, n27505, n27504, n27503, n27502, n23, 
            n53137, \data_in_frame[9][6] , \data_in_frame[11][3] , Kp_23__N_969, 
            n53140, Kp_23__N_645, \data_in_frame[11][4] , \data_in_frame[12][3] , 
            n23958, \data_in_frame[12][5] , n23338, \data_in_frame[12][1] , 
            Kp_23__N_675, n52656, n52455, n52831, n52848, n52925, 
            n22568, n151, n152, n490, n417, n344, n271, n198, 
            n125, \motor_state[23] , n9_adj_1, \motor_state[21] , \PID_CONTROLLER.integral_23__N_3691[23] , 
            \motor_state[20] , \motor_state[19] , n60212, n6, \PID_CONTROLLER.integral_23__N_3691[2] , 
            \PID_CONTROLLER.integral_23__N_3691[5] , \PID_CONTROLLER.integral_23__N_3691[9] , 
            \PID_CONTROLLER.integral_23__N_3691[8] , \PID_CONTROLLER.integral_23__N_3691[18] , 
            \PID_CONTROLLER.integral_23__N_3691[20] , \PID_CONTROLLER.integral_23__N_3691[22] , 
            \PID_CONTROLLER.integral_23__N_3691[19] , \PID_CONTROLLER.integral_23__N_3691[21] , 
            n11_adj_2, n4, n3, \data_in_frame[10][4] , n23375, n23824, 
            n53055, n47989, \data_in_frame[9][5] , \data_in_frame[11][6] , 
            n47452, n16, n52878, Kp_23__N_1724, n30905, n27611) /* synthesis syn_module_defined=1 */ ;
    input \Kp[3] ;
    input GND_net;
    input \Ki[15] ;
    output \PID_CONTROLLER.integral_23__N_3691[7] ;
    input \Kp[5] ;
    input \Kp[4] ;
    input [23:0]PWMLimit;
    input \Kp[0] ;
    input \Kp[1] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input [23:0]setpoint;
    input \motor_state[18] ;
    input n35;
    input \Kp[6] ;
    output n181;
    input [23:0]IntegralLimit;
    output n155;
    input \Ki[6] ;
    output \PID_CONTROLLER.integral_23__N_3691[12] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.integral_23__N_3691[6] ;
    input \Ki[0] ;
    input \Kp[2] ;
    input \Ki[7] ;
    input \Kp[12] ;
    input \Kp[7] ;
    input \Ki[2] ;
    input n11;
    input \Ki[3] ;
    input \Ki[8] ;
    input \Kp[13] ;
    input \Ki[14] ;
    output \PID_CONTROLLER.integral_23__N_3691[15] ;
    output \PID_CONTROLLER.integral_23__N_3691[14] ;
    output n375;
    input \PID_CONTROLLER.integral_23__N_3691[3] ;
    input \Ki[9] ;
    input \Ki[4] ;
    output n214;
    output \PID_CONTROLLER.integral_23__N_3691[16] ;
    output \PID_CONTROLLER.integral_23__N_3691[4] ;
    input \Kp[8] ;
    output \PID_CONTROLLER.integral_23__N_3691[0] ;
    input \Ki[12] ;
    input \Kp[14] ;
    input \Ki[5] ;
    input \Kp[15] ;
    input [23:0]deadband;
    input \motor_state[17] ;
    input \PID_CONTROLLER.integral_23__N_3691[11] ;
    input \Ki[10] ;
    input n5;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input n9;
    input \Ki[11] ;
    input \motor_state[12] ;
    input n545;
    output n143;
    output n220;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input VCC_net;
    input n472;
    input \motor_state[9] ;
    input \motor_state[8] ;
    output \PID_CONTROLLER.integral_23__N_3691[10] ;
    input n399;
    input n326;
    input n253;
    input n180;
    input \motor_state[7] ;
    input n53;
    input \motor_state[6] ;
    input n107;
    input \motor_state[5] ;
    output n203;
    input \motor_state[4] ;
    output n204;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \Kp[11] ;
    input \motor_state[1] ;
    input \Kp[9] ;
    input \motor_state[0] ;
    output \PID_CONTROLLER.integral_23__N_3691[1] ;
    input \Kp[10] ;
    output \PID_CONTROLLER.integral_23__N_3691[13] ;
    input \Ki[13] ;
    input n26922;
    output [23:0]\PID_CONTROLLER.integral ;
    input n27524;
    input n27523;
    input n27522;
    input n27521;
    input n27520;
    input n27519;
    input n27518;
    input n27517;
    input n27516;
    input n27515;
    input n27514;
    input n27513;
    input n27512;
    input n27511;
    input n27510;
    input n27509;
    input n27508;
    input n27507;
    input n27506;
    input n27505;
    input n27504;
    input n27503;
    input n27502;
    input n23;
    input n53137;
    input \data_in_frame[9][6] ;
    input \data_in_frame[11][3] ;
    input Kp_23__N_969;
    input n53140;
    input Kp_23__N_645;
    input \data_in_frame[11][4] ;
    input \data_in_frame[12][3] ;
    input n23958;
    input \data_in_frame[12][5] ;
    input n23338;
    input \data_in_frame[12][1] ;
    input Kp_23__N_675;
    input n52656;
    input n52455;
    input n52831;
    input n52848;
    input n52925;
    output n22568;
    output n151;
    output n152;
    input n490;
    input n417;
    input n344;
    input n271;
    input n198;
    input n125;
    input \motor_state[23] ;
    input n9_adj_1;
    input \motor_state[21] ;
    output \PID_CONTROLLER.integral_23__N_3691[23] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input n60212;
    input n6;
    output \PID_CONTROLLER.integral_23__N_3691[2] ;
    output \PID_CONTROLLER.integral_23__N_3691[5] ;
    output \PID_CONTROLLER.integral_23__N_3691[9] ;
    output \PID_CONTROLLER.integral_23__N_3691[8] ;
    output \PID_CONTROLLER.integral_23__N_3691[18] ;
    output \PID_CONTROLLER.integral_23__N_3691[20] ;
    output \PID_CONTROLLER.integral_23__N_3691[22] ;
    output \PID_CONTROLLER.integral_23__N_3691[19] ;
    output \PID_CONTROLLER.integral_23__N_3691[21] ;
    input n11_adj_2;
    input n4;
    input n3;
    input \data_in_frame[10][4] ;
    output n23375;
    input n23824;
    input n53055;
    input n47989;
    input \data_in_frame[9][5] ;
    input \data_in_frame[11][6] ;
    input n47452;
    output n16;
    input n52878;
    input Kp_23__N_1724;
    input n30905;
    output n27611;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n259, n1117, n393, n46645;
    wire [17:0]n14058;
    
    wire n524, n46646;
    wire [23:0]n356;
    
    wire n62959;
    wire [23:0]n382;
    
    wire n61311, n60843, n332, n55139, n24971, n9611;
    wire [23:0]n49;
    wire [1:0]n18250;
    
    wire n46561;
    wire [5:0]n18034;
    
    wire n487, n46562;
    wire [6:0]n17922;
    
    wire n414, n46560, n45589, n46185;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n46186, n45709;
    wire [23:0]n1_adj_4956;
    
    wire n45710, n46289;
    wire [11:0]n16802;
    
    wire n177, n46290, n45708;
    wire [31:0]n51;
    
    wire n46184, n45590;
    wire [12:0]n16438;
    
    wire n104, n46494;
    wire [21:0]n10158;
    
    wire n877, n46495, n46183, n62942;
    wire [18:0]n13337;
    
    wire n451, n46644, n405, n466;
    wire [23:0]n130;
    wire [23:0]n182;
    wire [23:0]n207;
    
    wire n366, n475, n61631, n92, n23_c, n62937, n439, n59952, 
        n490_c, n56230, n56232, n210, n62924, n56236, n45256, 
        n548, n61299, n62951, n56240;
    wire [3:0]n18202;
    
    wire n6_c, n8, n892, n61875, n62915, n478, n6_adj_4409, n4_c, 
        n54814, n62075, n62912, n539, n165, n27, n15, n13, n60043, 
        n238, n603, n33, n12, n965;
    wire [23:0]n1_adj_4957;
    
    wire n1041, n45707, n116, n47, n189, n10_adj_4413, n38, n229, 
        n554, n262, n512, n621, n676, n35_adj_4414, n30, n302, 
        n311, n122, n83, n14_adj_4417, n585, n9_c, n60088, n60943, 
        n293, n19, n17, n60933, n25, n23_adj_4420, n21, n61917, 
        n31, n29, n61341, n1023, n375_adj_4424, n366_adj_4425, n37, 
        n62002, n439_adj_4426, n195, n1114, n627, n1096, n700, 
        n448, n512_adj_4428, n268, n86, n17_adj_4429, n521, n594, 
        n6_adj_4432, n61575, n43, n16_c, n585_adj_4433, n38360, 
        n8_adj_4437, n46182, n45, n24_adj_4439, n45588, n60061, 
        n61576, n59991, n116_adj_4440, n47_adj_4441, n159, n618, 
        n189_adj_4443, n667, n740, n59989, n61169, counter_31__N_3690, 
        n45706;
    wire [8:0]n17697;
    wire [7:0]n17858;
    
    wire n335, n46374;
    wire [19:0]n12098;
    wire [18:0]n12938;
    
    wire n959, n46435, n46375, n378, n46643;
    wire [10:0]n17114;
    
    wire n910, n46288;
    wire [0:0]n10182;
    wire [21:0]n10689;
    
    wire n46748;
    wire [47:0]n257;
    
    wire n46747, n45587;
    wire [47:0]n306;
    
    wire n804, n46493, n46181, n45705, n45586, n46180, n45704, 
        n837, n46287, n262_adj_4448, n46373, n45703, n305, n46642, 
        n46179, n45585, n232, n46641, n46746, n764, n46286, n46178, 
        n45702, n45584, n341, n60507, n813, n658, n46745, n886, 
        n691, n46285, n46177, n12_adj_4454, n46176, n46744, n45701, 
        n731, n46492, n45583, n46175, n46436, n46434, n46491, 
        n46433, n46559, n46432, n46431, n46372, n46284, n46174, 
        n45700, n46640, n46283, n46173, n46743, n46172, n45699, 
        n45698, n45582, n45697, n45696, n45581, n45695, n59210, 
        n46282, n46171, n46170, n45694, n45693, n46490, n45692, 
        n45580, n46430, n45691, n45690, n45689, n46429, n45579, 
        n46742, n46558, n46489;
    wire [16:0]n14382;
    wire [15:0]n14994;
    
    wire n46371, n46281, n46169, n46168, n46280, n46370, n46428, 
        n4_adj_4461, n46741;
    wire [8:0]n17598;
    wire [7:0]n17778;
    
    wire n46639, n46740, n46638, n46369, n46279, n46557, n46278, 
        n46488, n61563, n46487, n46427, n46739, n61564, n45688, 
        n551, n45687, n45686, n45578, n45685, n46486, n59932, 
        n45684, n46426, n45683, n45577, n46637, n46425, n45682, 
        n62947, n46368, n45681;
    wire [5:0]n18082;
    
    wire n46277, n45680;
    wire [4:0]n18153;
    
    wire n417_c, n46276, n10_adj_4465, n156_adj_4466, n46424, n30_adj_4467, 
        n950, n46738, n45679, n62920, n60819, n59936, n968, n46367, 
        n481, n46636, n344_adj_4469, n46275, n45678, n45677, n45676, 
        n877_adj_4474, n46737, n45576, n4_adj_4475, n624, n45675, 
        n61865, n60519, n45674, n45575, n45673, n45672, n45574, 
        n895, n46366, n271_c, n46274, n694, n220_adj_4481, n46485, 
        n45573, n831, n45572, n658_adj_4482, n822, n46365, n767, 
        n840, n804_adj_4483, n46736;
    wire [13:0]n16242;
    wire [12:0]n16633;
    
    wire n1050, n46556, n977, n46555, n408, n46635, n74, n5_adj_4485, 
        n198_adj_4486, n46273, n335_adj_4487, n147_adj_4488, n46484, 
        n56, n125_adj_4489, n731_adj_4490, n46735, n904, n46554, 
        n749, n46364, n46634;
    wire [9:0]n17378;
    
    wire n46272, n46271, n46734, n46553, n46270;
    wire [20:0]n11174;
    
    wire n46483, n46733, n46363, n46269, n46732, n46633, n62041, 
        n62042, n6_adj_4491, n61565, n61566, n60831, n59910, n24_adj_4492, 
        n8_adj_4493, n62910, n59904, n61171, n60517, n62040, n59916, 
        n61775, n60525, n4_adj_4494, n61573, n61574, n60033, n60029, 
        n61847, n46632, n46362, n46268, n46731;
    wire [16:0]n14705;
    
    wire n46631, n46267, n46730, n46630, n60509, n293_adj_4495, 
        n46729, n220_adj_4497, n46728, n402_adj_4498, n46266, n530, 
        n46361, n46482;
    wire [9:0]n17498;
    
    wire n770, n46423, n758, n46552, n46629, n329, n46265, n457, 
        n46360, n46481, n147_adj_4499, n46727, n1111, n46628, n5_adj_4500, 
        n74_adj_4501, n685, n46551, n256, n46264, n1038, n46627;
    wire [0:0]n9651;
    
    wire n45640, n697, n46422, n612, n46550, n45639, n62108, n62109, 
        n45638, n39, n62061, n110_adj_4503, n41, n59995, n41_adj_4507;
    wire [20:0]n11657;
    
    wire n46726, n46725, n61773, n45637, n45636, n384_adj_4509, 
        n46359, n183_adj_4510, n46263, n46724, n46421, n46420, n46723, 
        n46358, n46480, n45635, n46626, n46357, n45634, n46356, 
        n46549, n60515, n61961, n61963, n46479, n46419, n46625, 
        n46722, n56216, n45633, n47_adj_4511, n46548, n46418, n45632, 
        n45631, n45630, n45629;
    wire [14:0]n15538;
    
    wire n46355, n46721, n45628, n46417, n45627, n46547, n46478, 
        n45626, n46354, n46416, n45625, n45624, n819, n46624, 
        n46720, n320, n46546, n1044, n46353, n46477, n45623, n1099, 
        n46719, n45622, n971, n46352, n45621, n45620, n45619, 
        n247, n46545, n746, n46623, n45445, n186_adj_4514, n46415, 
        n1026, n46718, n45618, n673, n46622, n953, n46717, n600, 
        n46621, n1099_adj_4515, n46476, n174, n46544, n880, n46716, 
        n44_adj_4516, n113_adj_4517, n807, n46715, n898, n46351, 
        n527, n46620, n45617, n45616, n734, n46714, n454, n46619, 
        n45615, n661, n46713, n825, n46350, n588, n46712, n45614, 
        n41_adj_4519, n39_adj_4520, n45_adj_4521, n33_adj_4522, n37_adj_4523, 
        n43_adj_4524, n9_adj_4525, n11_adj_4527, n13_adj_4528, n35_adj_4529, 
        n27_adj_4530, n29_adj_4531, n31_adj_4532, n21_adj_4533, n25_adj_4534, 
        n15_adj_4535, n17_adj_4536, n19_adj_4537, n59426, n60299, 
        n12_adj_4538, n10_adj_4539, n30_adj_4540, n59515, n60376, 
        n60336, n61721, n61413, n62008, n16_adj_4542, n6_adj_4543, 
        n61767, n61768, n8_adj_4544, n24_adj_4545, n45613, n60219;
    wire [17:0]n13698;
    
    wire n46414, n515, n46711, n46413, n32_adj_4546, n101, n442, 
        n46710, n752, n46349, n381, n46618, n369_adj_4547, n46709, 
        n60215, n61165, n679, n46348, n308, n46617, n296_adj_4548, 
        n46708, n61475, n235, n46616, n4_adj_4563, n61587, n162_adj_4564, 
        n46615, n61588;
    wire [11:0]n16970;
    
    wire n980, n46543, n60282, n907, n46542, n1026_adj_4565, n46475, 
        n223, n46707, n46412, n20_adj_4566, n89, n150_adj_4567, 
        n46706, n606, n46347, n45612, n8_adj_4568, n77;
    wire [19:0]n12538;
    
    wire n46705, n46704, n45611, n45610, n533, n46346, n834, n46541, 
        n45609, n22_adj_4569, n24_adj_4570, n60277, n61841, n23_adj_4571, 
        n45608, n460, n46345, n25_adj_4572, n10_adj_4573, n46411;
    wire [15:0]n15282;
    
    wire n46614, n46703, n45607, n46613, n46702, n45606, n953_adj_4574, 
        n46474, n387_adj_4575, n46344, n45605, n45604, n1114_adj_4576, 
        n46612, n761, n46540, n45603, n16_adj_4577, n45602, n46701, 
        n60489, n46700, n62104, n62105, n12_adj_4578, n1041_adj_4579, 
        n46611, n1102, n46699, n314, n46343, n688, n46539, n1029, 
        n46698, n45601, n241, n46342, n956, n46697, n45600, n615, 
        n46538, n883, n46696, n1108, n46410, n45599, n45598, n45597, 
        n1035, n46409, n542, n46537, n810, n46695, n968_adj_4581, 
        n46610, n168, n46341, n737, n46694, n880_adj_4582, n46473, 
        n664, n46693, n895_adj_4583, n46609, n45596, n807_adj_4585, 
        n46472, n962, n46408, n822_adj_4586, n46608, n62068, n26_adj_4587, 
        n95, n45595, n60223, n469, n46536;
    wire [6:0]n17985;
    
    wire n630, n46340, n61769, n591, n46692, n749_adj_4588, n46607, 
        n889, n46407, n557, n46339, n60495, n396_adj_4589, n46535, 
        n518, n46691, n676_adj_4590, n46606, n445, n46690, n734_adj_4591, 
        n46471, n372_adj_4592, n46689, n603_adj_4593, n46605, n299_adj_4594, 
        n46688, n61957, n484, n46338, n816, n46406, n226, n46687, 
        n153_adj_4595, n46686, n39_adj_4596, n530_adj_4597, n46604, 
        n323, n46534, n661_adj_4598, n46470, n457_adj_4599, n46603, 
        n411, n46337, n743, n46405, n41_adj_4600, n11_adj_4601, 
        n80, n338_adj_4602, n46336, n384_adj_4603, n46602, n670, 
        n46404, n588_adj_4604, n46469, n265, n46335, n250, n46533, 
        n770_adj_4605, n46685, n697_adj_4606, n46684, n624_adj_4607, 
        n46683, n192_adj_4608, n46334, n597, n46403, n515_adj_4609, 
        n46468, n524_adj_4610, n46402, n45_adj_4611, n43_adj_4612, 
        n177_adj_4613, n46532, n311_adj_4614, n46601, n551_adj_4615, 
        n46682, n50_adj_4616, n119_adj_4617, n478_adj_4618, n46681, 
        n442_adj_4619, n46467, n35_adj_4620, n104_adj_4621, n405_adj_4622, 
        n46680, n238_adj_4623, n46600;
    wire [13:0]n16018;
    
    wire n1120, n46333, n1047, n46332, n165_adj_4624, n46599, n332_adj_4625, 
        n46679, n55037, n46531, n451_adj_4627, n46401, n259_adj_4628, 
        n46678, n23_adj_4629, n92_adj_4630;
    wire [4:0]n18118;
    
    wire n46530, n630_adj_4632, n46598, n186_adj_4633, n46677, n557_adj_4634, 
        n46597, n484_adj_4635, n46596, n46529, n44_adj_4637, n113_adj_4638, 
        n411_adj_4639, n46595, n46528, n369_adj_4641, n46466, n338_adj_4642, 
        n46594, n46527, n296_adj_4644, n46465, n56_adj_4645, n223_adj_4647, 
        n46464, n27_adj_4648, n46676, n265_adj_4649, n46593, n46675, 
        n46674;
    wire [10:0]n17257;
    
    wire n910_adj_4650, n46526, n974, n46331, n837_adj_4651, n46525, 
        n901, n46330, n378_adj_4652, n46400, n828, n46329, n29_adj_4653, 
        n192_adj_4654, n46592, n764_adj_4655, n46524, n46673, n305_adj_4656, 
        n46399, n50_adj_4657, n119_adj_4658, n232_adj_4659, n46398, 
        n691_adj_4660, n46523, n150_adj_4661, n46463, n46672;
    wire [14:0]n15793;
    
    wire n46591, n618_adj_4662, n46522, n8_adj_4663, n77_adj_4664, 
        n1117_adj_4665, n46590, n545_adj_4666, n46521, n46462, n472_adj_4667, 
        n46520, n46461, n31_adj_4668, n1044_adj_4669, n46589, n399_adj_4670, 
        n46519, n46460, n1105, n46671, n326_adj_4671, n46518, n46459, 
        n755, n46328, n159_adj_4672, n46397, n682, n46327, n46458, 
        n609, n46326, n17_adj_4673, n86_adj_4674, n536, n46325, 
        n463, n46324, n971_adj_4675, n46588, n253_adj_4676, n46517, 
        n46457, n46396, n390_adj_4677, n46323, n46395, n317, n46322, 
        n1102_adj_4678, n46456, n244, n46321, n46394, n171, n46320, 
        n898_adj_4679, n46587, n180_adj_4680, n46516, n1029_adj_4681, 
        n46455, n29_adj_4682, n98, n21_adj_4683, n1111_adj_4684, n46393, 
        n1050_adj_4685, n46319, n977_adj_4686, n46318, n956_adj_4687, 
        n46454, n904_adj_4688, n46317, n1038_adj_4689, n46392, n831_adj_4690, 
        n46316, n38_adj_4691, n107_adj_4692, n883_adj_4693, n46453, 
        n965_adj_4694, n46391, n758_adj_4695, n46315, n1032, n46670, 
        n685_adj_4696, n46314, n892_adj_4697, n46390, n612_adj_4698, 
        n46313, n840_adj_4699, n46515, n810_adj_4700, n46452, n539_adj_4701, 
        n46312, n819_adj_4702, n46389, n466_adj_4703, n46311, n825_adj_4704, 
        n46586, n767_adj_4705, n46514, n694_adj_4706, n46513, n737_adj_4707, 
        n46451, n959_adj_4708, n46669, n752_adj_4709, n46585, n621_adj_4710, 
        n46512, n679_adj_4711, n46584, n548_adj_4712, n46511, n393_adj_4713, 
        n46310, n746_adj_4714, n46388, n23_adj_4715, n25_adj_4716, 
        n475_adj_4717, n46510, n320_adj_4718, n46309, n673_adj_4719, 
        n46387, n247_adj_4720, n46308, n664_adj_4721, n46450, n174_adj_4722, 
        n46307, n600_adj_4723, n46386, n32_adj_4724, n101_adj_4725, 
        n606_adj_4726, n46583, n402_adj_4727, n46509, n560, n46306, 
        n527_adj_4728, n46385, n487_adj_4729, n46305, n414_adj_4730, 
        n46304, n454_adj_4731, n46384, n591_adj_4732, n46449, n341_adj_4733, 
        n46303, n381_adj_4734, n46383, n268_adj_4735, n46302, n886_adj_4736, 
        n46668, n329_adj_4737, n46508, n45594, n195_adj_4738, n46301, 
        n53_adj_4739, n122_adj_4740, n308_adj_4741, n46382, n980_adj_4742, 
        n46300, n518_adj_4743, n46448, n907_adj_4744, n46299, n813_adj_4745, 
        n46667, n533_adj_4746, n46582;
    wire [23:0]n436;
    wire [23:0]n1_adj_4958;
    
    wire n45740, n460_adj_4748, n46581, n235_adj_4749, n46381, n834_adj_4750, 
        n46298, n45739, n256_adj_4752, n46507, n445_adj_4753, n46447, 
        n761_adj_4754, n46297, n45738, n740_adj_4757, n46666, n387_adj_4758, 
        n46580, n162_adj_4759, n46380, n688_adj_4760, n46296, n45737, 
        n615_adj_4762, n46295, n46198, n45593, n45736, n183_adj_4765, 
        n46506, n45735, n372_adj_4768, n46446, n46197, n314_adj_4769, 
        n46579, n45734, n299_adj_4771, n46445, n667_adj_4772, n46665, 
        n45733, n41_adj_4774, n110_adj_4775, n226_adj_4776, n46444, 
        n45732, n241_adj_4779, n46578, n153_adj_4780, n46443, n46196, 
        n45731, n45730, n542_adj_4783, n46294, n46195, n45592, n45729, 
        n20_adj_4786, n89_adj_4787, n46194, n45728, n469_adj_4789, 
        n46293, n46193, n594_adj_4790, n46664, n11_adj_4791, n80_adj_4792, 
        n9_adj_4793, n46505, n45727, n45726, n45591, n168_adj_4797, 
        n46577, n31_adj_4798, n29_adj_4799, n46192, n45725, n11_adj_4801, 
        n396_adj_4802, n46292, n27_adj_4803, n25_adj_4804, n45724, 
        n521_adj_4806, n46663, n45723, n45722, n448_adj_4810, n46662, 
        n26_adj_4811, n95_adj_4812, n46191, n45721, n375_adj_4814, 
        n46661, n1120_adj_4815, n46576, n13_adj_4816, n33_adj_4817, 
        n700_adj_4818, n46379, n45720, n13_adj_4821, n45719, n627_adj_4823, 
        n46378, n45718, n46190, n302_adj_4825, n46660, n15_adj_4826, 
        n1047_adj_4827, n46575, n46504, n229_adj_4828, n46659, n35_adj_4829, 
        n156_adj_4830, n46658, n46503, n46442, n974_adj_4831, n46574, 
        n46441, n323_adj_4832, n46291, n46189, n37_adj_4835, n45717, 
        n23_adj_4837, n46502, n901_adj_4838, n46573, n828_adj_4839, 
        n46572, n14_adj_4840, n83_adj_4841, n755_adj_4842, n46571, 
        n682_adj_4843, n46570, n46501, n46657, n46656, n46500, n37_adj_4844, 
        n250_adj_4845, n46188, n45716, n46655, n15_adj_4847, n46440, 
        n609_adj_4848, n46569, n46439, n554_adj_4849, n46377, n46654, 
        n46499, n536_adj_4850, n46568, n1108_adj_4851, n46653, n45715, 
        n45714, n45713, n46187, n45712, n46438, n46498, n41_adj_4856, 
        n1035_adj_4857, n46652, n17_adj_4858, n463_adj_4859, n46567, 
        n1105_adj_4860, n46437, n45711, n962_adj_4862, n46651, n481_adj_4863, 
        n46376, n19_adj_4864, n35_adj_4865, n19_adj_4867, n9_adj_4868, 
        n21_adj_4869, n13_adj_4870, n889_adj_4871, n46650, n39_adj_4872, 
        n390_adj_4873, n46566, n60165, n816_adj_4874, n46649, n1096_adj_4875, 
        n46497, n408_adj_4876, n60148, n15_adj_4877, n317_adj_4878, 
        n46565, n743_adj_4879, n46648, n244_adj_4880, n46564, n1023_adj_4881, 
        n46496, n1032_adj_4882, n12_adj_4883, n171_adj_4884, n46563, 
        n670_adj_4885, n46647, n29_adj_4886, n98_adj_4887, n950_adj_4888, 
        n560_adj_4889, n10_adj_4890, n17_adj_4891, n4_adj_4892, n61476, 
        n8_adj_4893, n33_adj_4894, n597_adj_4895, n30_adj_4896, n59657, 
        n61029, n61023, n60679, n61933;
    wire [2:0]n18233;
    
    wire n61217, n61379, n45363, n62006, n16_adj_4897, n61583, n61965, 
        n61584, n8_adj_4899, n61193, n45395, n24_adj_4900, n59659, 
        n4_adj_4901, n10_adj_4902, n60099, n61697, n60090, n61167, 
        n60497, n18_adj_4903, n4_adj_4904, n61581, n61582, n60140, 
        n60132, n61845, n60499, n62106, n62107, n16_adj_4905, n62065, 
        n60105, n61771, n36_adj_4906, n61698, n60505, n61959, n59604, 
        n9613, n25210, n25205, n59592, n61978, n61479;
    wire [3:0]n18178;
    
    wire n6_adj_4907, n25200;
    wire [1:0]n18242;
    
    wire n45231;
    wire [2:0]n18218;
    
    wire n56198, n14_adj_4908, n56202, n56200, n45429, n56208, n34138, 
        n4_adj_4909, n8_adj_4910, n12_adj_4911, n6_adj_4912, n25190, 
        n22_adj_4913, n25185, n59720, n61793, n25180, n25175, n61794, 
        n61493, n61458, n62110, n25170, n60539, n25165, n59794, 
        n62150, n25160, n62151, n59834, n25155, n25150, n62147, 
        n25145, n25140, n435, n25135, n25130, n25125, n409, n37_adj_4914, 
        n25120, n41_adj_4915, n39_adj_4916, n25115, n35_adj_4917, 
        n25110, n25105, n29_adj_4918, n31_adj_4919, n25100, n33_adj_4920, 
        n27_adj_4921, n17_adj_4922, n25_adj_4923, n45_adj_4924, n19_adj_4925, 
        n43_adj_4926, n23_adj_4927, n21_adj_4928, n55117, n59900, 
        n6_adj_4929, n20_adj_4930, n26_adj_4931, n12_adj_4932, n55108, 
        n10_adj_4933, n59873, n9_adj_4934, n24_adj_4935, n28_adj_4936, 
        n23_adj_4937, n59856, n12_adj_4939, n10_adj_4940, n30_adj_4941, 
        n60773, n4_adj_4942, n60761, n45272, n61839, n4_adj_4943, 
        n61255, n45313, n61982, n16_adj_4944, n61500, n61501, n8_adj_4947, 
        n24_adj_4948, n59796, n61173, n60527, n4_adj_4949, n61498, 
        n61499, n59841, n61871, n60529, n62050, n62051, n62036, 
        n59802, n61777, n60535, n59976, n60849, n62926, n59968, 
        n60839, n16_adj_4954, n59985, n62934, n59983, n62962;
    
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4550_8 (.CI(n46645), .I0(n14058[5]), .I1(n524), .CO(n46646));
    SB_LUT4 i45943_4_lut (.I0(n356[9]), .I1(n62959), .I2(n382[9]), .I3(n61311), 
            .O(n60843));
    defparam i45943_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24392_4_lut (.I0(PWMLimit[0]), .I1(n55139), .I2(n24971), 
            .I3(n9611), .O(n49[0]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24392_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i31694_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n18250[0]));   // verilog/motorControl.v(50[18:24])
    defparam i31694_4_lut.LUT_INIT = 16'h6ca0;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n49[0]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4843_7 (.CI(n46561), .I0(n18034[4]), .I1(n487), .CO(n46562));
    SB_LUT4 add_4843_6_lut (.I0(GND_net), .I1(n18034[3]), .I2(n414), .I3(n46560), 
            .O(n17922[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n45589), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_20 (.CI(n46185), .I0(GND_net), .I1(counter[18]), 
            .CO(n46186));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n45709), .I0(GND_net), .I1(n1_adj_4956[15]), 
            .CO(n45710));
    SB_CARRY add_4723_3 (.CI(n46289), .I0(n16802[0]), .I1(n177), .CO(n46290));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[14]), 
            .I3(n45708), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n45708), .I0(GND_net), .I1(n1_adj_4956[14]), 
            .CO(n45709));
    SB_LUT4 counter_1935_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n46184), .O(n51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_20 (.CI(n45589), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n45590));
    SB_LUT4 add_4723_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n16438[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_19 (.CI(n46184), .I0(GND_net), .I1(counter[17]), 
            .CO(n46185));
    SB_CARRY mult_17_add_1225_13 (.CI(n46494), .I0(n10158[10]), .I1(n877), 
            .CO(n46495));
    SB_CARRY add_4723_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n46289));
    SB_LUT4 counter_1935_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n46183), .O(n51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i21_rep_124_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n62942));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i21_rep_124_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4550_7_lut (.I0(GND_net), .I1(n14058[4]), .I2(n451), .I3(n46644), 
            .O(n13337[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[7] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46731_4_lut (.I0(n356[11]), .I1(n62942), .I2(n382[11]), .I3(n60843), 
            .O(n61631));
    defparam i46731_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i25_rep_119_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n62937));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i25_rep_119_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45052_4_lut (.I0(n356[13]), .I1(n62937), .I2(n382[13]), .I3(n61631), 
            .O(n59952));
    defparam i45052_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n1[19]), .I3(n1[18]), 
            .O(n56230));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n56230), .I2(n1[20]), .I3(GND_net), 
            .O(n56232));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n1[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i29_rep_106_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n62924));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i29_rep_106_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_945 (.I0(\Kp[1] ), .I1(n210), .I2(n1[22]), .I3(n56232), 
            .O(n56236));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h936c;
    SB_LUT4 i31696_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n45256));   // verilog/motorControl.v(50[18:24])
    defparam i31696_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46399_4_lut (.I0(n356[15]), .I1(n62924), .I2(n382[15]), .I3(n59952), 
            .O(n61299));
    defparam i46399_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i33_rep_133_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n62951));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i33_rep_133_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_946 (.I0(n45256), .I1(\Kp[0] ), .I2(n56236), 
            .I3(n1[23]), .O(n56240));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h695a;
    SB_LUT4 i31898_4_lut (.I0(n18202[2]), .I1(\Kp[4] ), .I2(n6_c), .I3(n1[18]), 
            .O(n8));   // verilog/motorControl.v(50[18:24])
    defparam i31898_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46975_4_lut (.I0(n356[17]), .I1(n62951), .I2(n382[17]), .I3(n61299), 
            .O(n61875));
    defparam i46975_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i37_rep_97_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n62915));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i37_rep_97_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n6_adj_4409), .I1(n8), .I2(n4_c), .I3(n56240), 
            .O(n54814));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i47175_4_lut (.I0(n356[19]), .I1(n62915), .I2(n382[19]), .I3(n61875), 
            .O(n62075));
    defparam i47175_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i41_rep_94_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n62912));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i41_rep_94_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45143_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n60043));
    defparam i45143_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[10]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[11]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[13]), 
            .I3(n45707), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n45707), .I0(GND_net), .I1(n1_adj_4956[13]), 
            .CO(n45708));
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[15] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n207[12]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i13_3_lut (.I0(n207[12]), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[12] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n375), .I1(n356[6]), .I2(n13), 
            .I3(GND_net), .O(n10_adj_4413));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12), .I1(n356[17]), .I2(n35_adj_4414), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[12]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n214));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[4] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4417));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46043_4_lut (.I0(n13), .I1(n11), .I2(n9_c), .I3(n60088), 
            .O(n60943));
    defparam i46043_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[0] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[13]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46033_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n60943), 
            .O(n60933));
    defparam i46033_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[14]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47017_4_lut (.I0(n25), .I1(n23_adj_4420), .I2(n21), .I3(n60933), 
            .O(n61917));
    defparam i47017_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46441_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n61917), 
            .O(n61341));
    defparam i46441_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[15]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[16]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[17]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4424));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4425));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47102_4_lut (.I0(n37), .I1(n35_adj_4414), .I2(n33), .I3(n61341), 
            .O(n62002));
    defparam i47102_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4426));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[6] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1935_add_4_18 (.CI(n46183), .I0(GND_net), .I1(counter[16]), 
            .CO(n46184));
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[14] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4428));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4429));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[18]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[19]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[20]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[21]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46675_3_lut (.I0(n6_adj_4432), .I1(n356[10]), .I2(n21), .I3(GND_net), 
            .O(n61575));   // verilog/motorControl.v(51[12:29])
    defparam i46675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43), 
            .I3(GND_net), .O(n16_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4433));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[22]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[23]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24769_1_lut (.I0(n356[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38360));   // verilog/motorControl.v(50[18:38])
    defparam i24769_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[0]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[1]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[2]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[3]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[4]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[5]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17), 
            .I3(GND_net), .O(n8_adj_4437));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1935_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n46182), .O(n51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_c), .I1(n356[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4439));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n45588), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_19 (.CI(n45588), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n45589));
    SB_LUT4 i45161_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9_c), .O(n60061));
    defparam i45161_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46676_3_lut (.I0(n61575), .I1(n356[11]), .I2(n23_adj_4420), 
            .I3(GND_net), .O(n61576));   // verilog/motorControl.v(51[12:29])
    defparam i46676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45091_4_lut (.I0(n43), .I1(n25), .I2(n23_adj_4420), .I3(n60061), 
            .O(n59991));
    defparam i45091_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4440));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4441));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[6]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4443));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46269_4_lut (.I0(n24_adj_4439), .I1(n8_adj_4437), .I2(n45), 
            .I3(n59989), .O(n61169));   // verilog/motorControl.v(51[12:29])
    defparam i46269_4_lut.LUT_INIT = 16'haaac;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3690));   // verilog/motorControl.v(23[10] 30[6])
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[12]), 
            .I3(n45706), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_7 (.CI(n46644), .I0(n14058[4]), .I1(n451), .CO(n46645));
    SB_LUT4 add_4820_5_lut (.I0(GND_net), .I1(n17858[2]), .I2(n335), .I3(n46374), 
            .O(n17697[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_14_lut (.I0(GND_net), .I1(n12938[11]), .I2(n959), 
            .I3(n46435), .O(n12098[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4820_5 (.CI(n46374), .I0(n17858[2]), .I1(n335), .CO(n46375));
    SB_LUT4 add_4550_6_lut (.I0(GND_net), .I1(n14058[3]), .I2(n378), .I3(n46643), 
            .O(n13337[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4748_13_lut (.I0(GND_net), .I1(n17114[10]), .I2(n910), 
            .I3(n46288), .O(n16802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_17 (.CI(n46182), .I0(GND_net), .I1(counter[15]), 
            .CO(n46183));
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n1[23]), .I1(n10689[21]), .I2(GND_net), 
            .I3(n46748), .O(n10182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n10689[20]), .I2(GND_net), 
            .I3(n46747), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_6 (.CI(n46643), .I0(n14058[3]), .I1(n378), .CO(n46644));
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(n5), 
            .I3(n45587), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n45706), .I0(GND_net), .I1(n1_adj_4956[12]), 
            .CO(n45707));
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n10158[9]), .I2(n804), 
            .I3(n46493), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n46181), .O(n51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_18 (.CI(n45587), .I0(setpoint[16]), .I1(n5), 
            .CO(n45588));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[11]), 
            .I3(n45705), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n45586), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n45705), .I0(GND_net), .I1(n1_adj_4956[11]), 
            .CO(n45706));
    SB_CARRY counter_1935_add_4_16 (.CI(n46181), .I0(GND_net), .I1(counter[14]), 
            .CO(n46182));
    SB_LUT4 counter_1935_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n46180), .O(n51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[10]), 
            .I3(n45704), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n45704), .I0(GND_net), .I1(n1_adj_4956[10]), 
            .CO(n45705));
    SB_LUT4 add_4748_12_lut (.I0(GND_net), .I1(n17114[9]), .I2(n837), 
            .I3(n46287), .O(n16802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4820_4_lut (.I0(GND_net), .I1(n17858[1]), .I2(n262_adj_4448), 
            .I3(n46373), .O(n17697[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_15 (.CI(n46180), .I0(GND_net), .I1(counter[13]), 
            .CO(n46181));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[9]), 
            .I3(n45703), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_12 (.CI(n46287), .I0(n17114[9]), .I1(n837), .CO(n46288));
    SB_CARRY mult_16_add_1225_23 (.CI(n46747), .I0(n10689[20]), .I1(GND_net), 
            .CO(n46748));
    SB_LUT4 add_4550_5_lut (.I0(GND_net), .I1(n14058[2]), .I2(n305), .I3(n46642), 
            .O(n13337[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_17 (.CI(n45586), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n45587));
    SB_CARRY mult_17_add_1225_12 (.CI(n46493), .I0(n10158[9]), .I1(n804), 
            .CO(n46494));
    SB_LUT4 counter_1935_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n46179), .O(n51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n45585), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n45703), .I0(GND_net), .I1(n1_adj_4956[9]), 
            .CO(n45704));
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1935_add_4_14 (.CI(n46179), .I0(GND_net), .I1(counter[12]), 
            .CO(n46180));
    SB_CARRY add_4550_5 (.CI(n46642), .I0(n14058[2]), .I1(n305), .CO(n46643));
    SB_CARRY sub_8_add_2_16 (.CI(n45585), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n45586));
    SB_LUT4 add_4550_4_lut (.I0(GND_net), .I1(n14058[1]), .I2(n232), .I3(n46641), 
            .O(n13337[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n10689[19]), .I2(GND_net), 
            .I3(n46746), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4748_11_lut (.I0(GND_net), .I1(n17114[8]), .I2(n764), 
            .I3(n46286), .O(n16802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n46178), .O(n51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[8]), 
            .I3(n45702), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n45702), .I0(GND_net), .I1(n1_adj_4956[8]), 
            .CO(n45703));
    SB_CARRY add_4550_4 (.CI(n46641), .I0(n14058[1]), .I1(n232), .CO(n46642));
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(n9), 
            .I3(n45584), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_22 (.CI(n46746), .I0(n10689[19]), .I1(GND_net), 
            .CO(n46747));
    SB_CARRY counter_1935_add_4_13 (.CI(n46178), .I0(GND_net), .I1(counter[11]), 
            .CO(n46179));
    SB_LUT4 i45607_3_lut (.I0(n61576), .I1(n356[12]), .I2(n25), .I3(GND_net), 
            .O(n60507));   // verilog/motorControl.v(51[12:29])
    defparam i45607_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4748_11 (.CI(n46286), .I0(n17114[8]), .I1(n764), .CO(n46287));
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n10689[18]), .I2(GND_net), 
            .I3(n46745), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4820_4 (.CI(n46373), .I0(n17858[1]), .I1(n262_adj_4448), 
            .CO(n46374));
    SB_LUT4 add_4748_10_lut (.I0(GND_net), .I1(n17114[7]), .I2(n691), 
            .I3(n46285), .O(n16802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n46177), .O(n51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_12 (.CI(n46177), .I0(GND_net), .I1(counter[10]), 
            .CO(n46178));
    SB_CARRY mult_16_add_1225_21 (.CI(n46745), .I0(n10689[18]), .I1(GND_net), 
            .CO(n46746));
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_4454));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 counter_1935_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n46176), .O(n51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n10689[17]), .I2(GND_net), 
            .I3(n46744), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[7]), 
            .I3(n45701), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_15 (.CI(n45584), .I0(setpoint[13]), .I1(n9), 
            .CO(n45585));
    SB_CARRY add_4748_10 (.CI(n46285), .I0(n17114[7]), .I1(n691), .CO(n46286));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n10158[8]), .I2(n731), 
            .I3(n46492), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n45583), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4843_6 (.CI(n46560), .I0(n18034[3]), .I1(n414), .CO(n46561));
    SB_CARRY unary_minus_20_add_3_9 (.CI(n45701), .I0(GND_net), .I1(n1_adj_4956[7]), 
            .CO(n45702));
    SB_CARRY counter_1935_add_4_11 (.CI(n46176), .I0(GND_net), .I1(counter[9]), 
            .CO(n46177));
    SB_LUT4 counter_1935_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n46175), .O(n51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_11 (.CI(n46492), .I0(n10158[8]), .I1(n731), 
            .CO(n46493));
    SB_CARRY add_4492_14 (.CI(n46435), .I0(n12938[11]), .I1(n959), .CO(n46436));
    SB_LUT4 add_4492_13_lut (.I0(GND_net), .I1(n12938[10]), .I2(n886), 
            .I3(n46434), .O(n12098[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n10158[7]), .I2(n658), 
            .I3(n46491), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_10 (.CI(n46175), .I0(GND_net), .I1(counter[8]), 
            .CO(n46176));
    SB_CARRY add_4492_13 (.CI(n46434), .I0(n12938[10]), .I1(n886), .CO(n46435));
    SB_LUT4 add_4492_12_lut (.I0(GND_net), .I1(n12938[9]), .I2(n813), 
            .I3(n46433), .O(n12098[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_12 (.CI(n46433), .I0(n12938[9]), .I1(n813), .CO(n46434));
    SB_LUT4 add_4843_5_lut (.I0(GND_net), .I1(n18034[2]), .I2(n341), .I3(n46559), 
            .O(n17922[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_10 (.CI(n46491), .I0(n10158[7]), .I1(n658), 
            .CO(n46492));
    SB_LUT4 add_4492_11_lut (.I0(GND_net), .I1(n12938[8]), .I2(n740), 
            .I3(n46432), .O(n12098[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_11 (.CI(n46432), .I0(n12938[8]), .I1(n740), .CO(n46433));
    SB_CARRY sub_8_add_2_14 (.CI(n45583), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n45584));
    SB_LUT4 add_4492_10_lut (.I0(GND_net), .I1(n12938[7]), .I2(n667), 
            .I3(n46431), .O(n12098[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4820_3_lut (.I0(GND_net), .I1(n17858[0]), .I2(n189_adj_4443), 
            .I3(n46372), .O(n17697[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4820_3 (.CI(n46372), .I0(n17858[0]), .I1(n189_adj_4443), 
            .CO(n46373));
    SB_LUT4 add_4748_9_lut (.I0(GND_net), .I1(n17114[6]), .I2(n618), .I3(n46284), 
            .O(n16802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n46174), .O(n51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_9 (.CI(n46284), .I0(n17114[6]), .I1(n618), .CO(n46285));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[6]), 
            .I3(n45700), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4550_3_lut (.I0(GND_net), .I1(n14058[0]), .I2(n159), .I3(n46640), 
            .O(n13337[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4820_2_lut (.I0(GND_net), .I1(n47_adj_4441), .I2(n116_adj_4440), 
            .I3(GND_net), .O(n17697[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_9 (.CI(n46174), .I0(GND_net), .I1(counter[7]), 
            .CO(n46175));
    SB_LUT4 add_4748_8_lut (.I0(GND_net), .I1(n17114[5]), .I2(n545), .I3(n46283), 
            .O(n16802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n45700), .I0(GND_net), .I1(n1_adj_4956[6]), 
            .CO(n45701));
    SB_CARRY add_4820_2 (.CI(GND_net), .I0(n47_adj_4441), .I1(n116_adj_4440), 
            .CO(n46372));
    SB_CARRY mult_16_add_1225_20 (.CI(n46744), .I0(n10689[17]), .I1(GND_net), 
            .CO(n46745));
    SB_LUT4 counter_1935_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n46173), .O(n51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n10689[16]), .I2(GND_net), 
            .I3(n46743), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i12_3_lut (.I0(n143), .I1(n182[11]), .I2(n181), .I3(GND_net), 
            .O(n220));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_19 (.CI(n46743), .I0(n10689[16]), .I1(GND_net), 
            .CO(n46744));
    SB_CARRY counter_1935_add_4_8 (.CI(n46173), .I0(GND_net), .I1(counter[6]), 
            .CO(n46174));
    SB_CARRY add_4748_8 (.CI(n46283), .I0(n17114[5]), .I1(n545), .CO(n46284));
    SB_LUT4 counter_1935_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n46172), .O(n51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[5]), 
            .I3(n45699), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n45699), .I0(GND_net), .I1(n1_adj_4956[5]), 
            .CO(n45700));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[4]), 
            .I3(n45698), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n45698), .I0(GND_net), .I1(n1_adj_4956[4]), 
            .CO(n45699));
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n45582), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[3]), 
            .I3(n45697), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n45697), .I0(GND_net), .I1(n1_adj_4956[3]), 
            .CO(n45698));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[2]), 
            .I3(n45696), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_13 (.CI(n45582), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n45583));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n45696), .I0(GND_net), .I1(n1_adj_4956[2]), 
            .CO(n45697));
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n45581), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[1]), 
            .I3(n45695), .O(n382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n45695), .I0(GND_net), .I1(n1_adj_4956[1]), 
            .CO(n45696));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n38360), .I1(GND_net), .I2(n1_adj_4956[0]), 
            .I3(VCC_net), .O(n59210)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_8_add_2_12 (.CI(n45581), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n45582));
    SB_LUT4 add_4748_7_lut (.I0(GND_net), .I1(n17114[4]), .I2(n472), .I3(n46282), 
            .O(n16802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4956[0]), 
            .CO(n45695));
    SB_CARRY add_4550_3 (.CI(n46640), .I0(n14058[0]), .I1(n159), .CO(n46641));
    SB_CARRY counter_1935_add_4_7 (.CI(n46172), .I0(GND_net), .I1(counter[5]), 
            .CO(n46173));
    SB_CARRY add_4748_7 (.CI(n46282), .I0(n17114[4]), .I1(n472), .CO(n46283));
    SB_LUT4 counter_1935_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n46171), .O(n51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_6 (.CI(n46171), .I0(GND_net), .I1(counter[4]), 
            .CO(n46172));
    SB_CARRY add_4843_5 (.CI(n46559), .I0(n18034[2]), .I1(n341), .CO(n46560));
    SB_LUT4 counter_1935_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n46170), .O(n51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[23]), 
            .I3(n45694), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[22]), 
            .I3(n45693), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n10158[6]), .I2(n585_adj_4433), 
            .I3(n46490), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n45693), .I0(GND_net), .I1(n1_adj_4957[22]), 
            .CO(n45694));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[21]), 
            .I3(n45692), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_10 (.CI(n46431), .I0(n12938[7]), .I1(n667), .CO(n46432));
    SB_CARRY unary_minus_13_add_3_23 (.CI(n45692), .I0(GND_net), .I1(n1_adj_4957[21]), 
            .CO(n45693));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n45580), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_5 (.CI(n46170), .I0(GND_net), .I1(counter[3]), 
            .CO(n46171));
    SB_LUT4 add_4492_9_lut (.I0(GND_net), .I1(n12938[6]), .I2(n594), .I3(n46430), 
            .O(n12098[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[20]), 
            .I3(n45691), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n45691), .I0(GND_net), .I1(n1_adj_4957[20]), 
            .CO(n45692));
    SB_CARRY mult_17_add_1225_9 (.CI(n46490), .I0(n10158[6]), .I1(n585_adj_4433), 
            .CO(n46491));
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[19]), 
            .I3(n45690), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_21 (.CI(n45690), .I0(GND_net), .I1(n1_adj_4957[19]), 
            .CO(n45691));
    SB_CARRY add_4492_9 (.CI(n46430), .I0(n12938[6]), .I1(n594), .CO(n46431));
    SB_CARRY sub_8_add_2_11 (.CI(n45580), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n45581));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[18]), 
            .I3(n45689), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_8_lut (.I0(GND_net), .I1(n12938[5]), .I2(n521), .I3(n46429), 
            .O(n12098[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n45579), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n10689[15]), .I2(GND_net), 
            .I3(n46742), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_18 (.CI(n46742), .I0(n10689[15]), .I1(GND_net), 
            .CO(n46743));
    SB_LUT4 add_4550_2_lut (.I0(GND_net), .I1(n17_adj_4429), .I2(n86), 
            .I3(GND_net), .O(n13337[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4843_4_lut (.I0(GND_net), .I1(n18034[1]), .I2(n268), .I3(n46558), 
            .O(n17922[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n10158[5]), .I2(n512_adj_4428), 
            .I3(n46489), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_8 (.CI(n46429), .I0(n12938[5]), .I1(n521), .CO(n46430));
    SB_LUT4 add_4603_18_lut (.I0(GND_net), .I1(n14994[15]), .I2(GND_net), 
            .I3(n46371), .O(n14382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4748_6_lut (.I0(GND_net), .I1(n17114[3]), .I2(n399), .I3(n46281), 
            .O(n16802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n46169), .O(n51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_4 (.CI(n46169), .I0(GND_net), .I1(counter[2]), 
            .CO(n46170));
    SB_CARRY add_4748_6 (.CI(n46281), .I0(n17114[3]), .I1(n399), .CO(n46282));
    SB_LUT4 counter_1935_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n46168), .O(n51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_3 (.CI(n46168), .I0(GND_net), .I1(counter[1]), 
            .CO(n46169));
    SB_LUT4 add_4748_5_lut (.I0(GND_net), .I1(n17114[2]), .I2(n326), .I3(n46280), 
            .O(n16802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_17_lut (.I0(GND_net), .I1(n14994[14]), .I2(GND_net), 
            .I3(n46370), .O(n14382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_17 (.CI(n46370), .I0(n14994[14]), .I1(GND_net), 
            .CO(n46371));
    SB_CARRY add_4748_5 (.CI(n46280), .I0(n17114[2]), .I1(n326), .CO(n46281));
    SB_CARRY add_4843_4 (.CI(n46558), .I0(n18034[1]), .I1(n268), .CO(n46559));
    SB_LUT4 add_4492_7_lut (.I0(GND_net), .I1(n12938[4]), .I2(n448), .I3(n46428), 
            .O(n12098[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i4_3_lut (.I0(n59210), .I1(n382[1]), .I2(n356[1]), 
            .I3(GND_net), .O(n4_adj_4461));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n10689[14]), .I2(GND_net), 
            .I3(n46741), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_2 (.CI(GND_net), .I0(n17_adj_4429), .I1(n86), .CO(n46640));
    SB_CARRY mult_16_add_1225_17 (.CI(n46741), .I0(n10689[14]), .I1(GND_net), 
            .CO(n46742));
    SB_LUT4 add_4811_10_lut (.I0(GND_net), .I1(n17778[7]), .I2(n700), 
            .I3(n46639), .O(n17598[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n10689[13]), .I2(n1096), 
            .I3(n46740), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_16 (.CI(n46740), .I0(n10689[13]), .I1(n1096), 
            .CO(n46741));
    SB_LUT4 add_4811_9_lut (.I0(GND_net), .I1(n17778[6]), .I2(n627), .I3(n46638), 
            .O(n17598[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_16_lut (.I0(GND_net), .I1(n14994[13]), .I2(n1114), 
            .I3(n46369), .O(n14382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4748_4_lut (.I0(GND_net), .I1(n17114[1]), .I2(n253), .I3(n46279), 
            .O(n16802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_7 (.CI(n46428), .I0(n12938[4]), .I1(n448), .CO(n46429));
    SB_CARRY counter_1935_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n46168));
    SB_CARRY add_4748_4 (.CI(n46279), .I0(n17114[1]), .I1(n253), .CO(n46280));
    SB_CARRY mult_17_add_1225_8 (.CI(n46489), .I0(n10158[5]), .I1(n512_adj_4428), 
            .CO(n46490));
    SB_LUT4 add_4843_3_lut (.I0(GND_net), .I1(n18034[0]), .I2(n195), .I3(n46557), 
            .O(n17922[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4748_3_lut (.I0(GND_net), .I1(n17114[0]), .I2(n180), .I3(n46278), 
            .O(n16802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n10158[4]), .I2(n439_adj_4426), 
            .I3(n46488), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_7 (.CI(n46488), .I0(n10158[4]), .I1(n439_adj_4426), 
            .CO(n46489));
    SB_LUT4 i46663_3_lut (.I0(n4_adj_4461), .I1(n382[13]), .I2(n356[13]), 
            .I3(GND_net), .O(n61563));   // verilog/motorControl.v(51[33:53])
    defparam i46663_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n10158[3]), .I2(n366_adj_4425), 
            .I3(n46487), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n45689), .I0(GND_net), .I1(n1_adj_4957[18]), 
            .CO(n45690));
    SB_CARRY mult_17_add_1225_6 (.CI(n46487), .I0(n10158[3]), .I1(n366_adj_4425), 
            .CO(n46488));
    SB_LUT4 add_4492_6_lut (.I0(GND_net), .I1(n12938[3]), .I2(n375_adj_4424), 
            .I3(n46427), .O(n12098[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_6 (.CI(n46427), .I0(n12938[3]), .I1(n375_adj_4424), 
            .CO(n46428));
    SB_CARRY sub_8_add_2_10 (.CI(n45579), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n45580));
    SB_CARRY add_4603_16 (.CI(n46369), .I0(n14994[13]), .I1(n1114), .CO(n46370));
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n10689[12]), .I2(n1023), 
            .I3(n46739), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46664_3_lut (.I0(n61563), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n61564));   // verilog/motorControl.v(51[33:53])
    defparam i46664_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[17]), 
            .I3(n45688), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_3 (.CI(n46278), .I0(n17114[0]), .I1(n180), .CO(n46279));
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n45688), .I0(GND_net), .I1(n1_adj_4957[17]), 
            .CO(n45689));
    SB_CARRY add_4811_9 (.CI(n46638), .I0(n17778[6]), .I1(n627), .CO(n46639));
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[16]), 
            .I3(n45687), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_18 (.CI(n45687), .I0(GND_net), .I1(n1_adj_4957[16]), 
            .CO(n45688));
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[15]), 
            .I3(n45686), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n45578), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n45686), .I0(GND_net), .I1(n1_adj_4957[15]), 
            .CO(n45687));
    SB_CARRY mult_16_add_1225_15 (.CI(n46739), .I0(n10689[12]), .I1(n1023), 
            .CO(n46740));
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[14]), 
            .I3(n45685), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_9 (.CI(n45578), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n45579));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n10158[2]), .I2(n293), 
            .I3(n46486), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_16 (.CI(n45685), .I0(GND_net), .I1(n1_adj_4957[14]), 
            .CO(n45686));
    SB_LUT4 i45032_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n59932));
    defparam i45032_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[13]), 
            .I3(n45684), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4843_3 (.CI(n46557), .I0(n18034[0]), .I1(n195), .CO(n46558));
    SB_LUT4 add_4843_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n17922[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_5_lut (.I0(GND_net), .I1(n12938[2]), .I2(n302), .I3(n46426), 
            .O(n12098[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n45684), .I0(GND_net), .I1(n1_adj_4957[13]), 
            .CO(n45685));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[12]), 
            .I3(n45683), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n45577), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4811_8_lut (.I0(GND_net), .I1(n17778[5]), .I2(n554), .I3(n46637), 
            .O(n17598[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_5 (.CI(n46426), .I0(n12938[2]), .I1(n302), .CO(n46427));
    SB_LUT4 add_4492_4_lut (.I0(GND_net), .I1(n12938[1]), .I2(n229), .I3(n46425), 
            .O(n12098[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n45683), .I0(GND_net), .I1(n1_adj_4957[12]), 
            .CO(n45684));
    SB_LUT4 add_4748_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n16802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[11]), 
            .I3(n45682), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i35_rep_129_2_lut (.I0(n356[17]), .I1(n382[17]), 
            .I2(GND_net), .I3(GND_net), .O(n62947));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i35_rep_129_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4603_15_lut (.I0(GND_net), .I1(n14994[12]), .I2(n1041), 
            .I3(n46368), .O(n14382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n45682), .I0(GND_net), .I1(n1_adj_4957[11]), 
            .CO(n45683));
    SB_CARRY add_4603_15 (.CI(n46368), .I0(n14994[12]), .I1(n1041), .CO(n46369));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[10]), 
            .I3(n45681), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n46278));
    SB_LUT4 add_4862_7_lut (.I0(GND_net), .I1(n54814), .I2(n490_c), .I3(n46277), 
            .O(n18082[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n45681), .I0(GND_net), .I1(n1_adj_4957[10]), 
            .CO(n45682));
    SB_CARRY add_4492_4 (.CI(n46425), .I0(n12938[1]), .I1(n229), .CO(n46426));
    SB_CARRY sub_8_add_2_8 (.CI(n45577), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n45578));
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[9]), 
            .I3(n45680), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4862_6_lut (.I0(GND_net), .I1(n18153[3]), .I2(n417_c), 
            .I3(n46276), .O(n18082[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4862_6 (.CI(n46276), .I0(n18153[3]), .I1(n417_c), .CO(n46277));
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_4465));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4492_3_lut (.I0(GND_net), .I1(n12938[0]), .I2(n156_adj_4466), 
            .I3(n46424), .O(n12098[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_4454), .I1(n382[17]), .I2(n356[17]), 
            .I3(GND_net), .O(n30_adj_4467));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n45680), .I0(GND_net), .I1(n1_adj_4957[9]), 
            .CO(n45681));
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n10689[11]), .I2(n950), 
            .I3(n46738), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[8]), 
            .I3(n45679), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45036_4_lut (.I0(n356[16]), .I1(n62920), .I2(n382[16]), .I3(n60819), 
            .O(n59936));
    defparam i45036_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_4811_8 (.CI(n46637), .I0(n17778[5]), .I1(n554), .CO(n46638));
    SB_LUT4 add_4603_14_lut (.I0(GND_net), .I1(n14994[11]), .I2(n968), 
            .I3(n46367), .O(n14382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4811_7_lut (.I0(GND_net), .I1(n17778[4]), .I2(n481), .I3(n46636), 
            .O(n17598[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n45679), .I0(GND_net), .I1(n1_adj_4957[8]), 
            .CO(n45680));
    SB_LUT4 add_4862_5_lut (.I0(GND_net), .I1(n18153[2]), .I2(n344_adj_4469), 
            .I3(n46275), .O(n18082[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[7]), 
            .I3(n45678), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n45678), .I0(GND_net), .I1(n1_adj_4957[7]), 
            .CO(n45679));
    SB_CARRY mult_17_add_1225_5 (.CI(n46486), .I0(n10158[2]), .I1(n293), 
            .CO(n46487));
    SB_CARRY add_4603_14 (.CI(n46367), .I0(n14994[11]), .I1(n968), .CO(n46368));
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[7]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_16_add_1225_14 (.CI(n46738), .I0(n10689[11]), .I1(n950), 
            .CO(n46739));
    SB_CARRY add_4862_5 (.CI(n46275), .I0(n18153[2]), .I1(n344_adj_4469), 
            .CO(n46276));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[6]), 
            .I3(n45677), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n45677), .I0(GND_net), .I1(n1_adj_4957[6]), 
            .CO(n45678));
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[5]), 
            .I3(n45676), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n45676), .I0(GND_net), .I1(n1_adj_4957[5]), 
            .CO(n45677));
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n10689[10]), .I2(n877_adj_4474), 
            .I3(n46737), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n45576), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31890_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4475), 
            .I3(n18202[1]), .O(n6_c));   // verilog/motorControl.v(50[18:24])
    defparam i31890_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[4]), 
            .I3(n45675), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46965_4_lut (.I0(n30_adj_4467), .I1(n10_adj_4465), .I2(n62947), 
            .I3(n59932), .O(n61865));   // verilog/motorControl.v(51[33:53])
    defparam i46965_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n45675), .I0(GND_net), .I1(n1_adj_4957[4]), 
            .CO(n45676));
    SB_LUT4 i45619_3_lut (.I0(n61564), .I1(n382[15]), .I2(n356[15]), .I3(GND_net), 
            .O(n60519));   // verilog/motorControl.v(51[33:53])
    defparam i45619_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[3]), 
            .I3(n45674), .O(n203)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_5 (.CI(n45674), .I0(GND_net), .I1(n1_adj_4957[3]), 
            .CO(n45675));
    SB_CARRY sub_8_add_2_7 (.CI(n45576), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n45577));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n45575), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[2]), 
            .I3(n45673), .O(n204)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n45673), .I0(GND_net), .I1(n1_adj_4957[2]), 
            .CO(n45674));
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[1]), 
            .I3(n45672), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n45672), .I0(GND_net), .I1(n1_adj_4957[1]), 
            .CO(n45673));
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4957[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_6 (.CI(n45575), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n45576));
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4957[0]), 
            .CO(n45672));
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(\motor_state[3] ), 
            .I3(n45574), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_5 (.CI(n45574), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n45575));
    SB_LUT4 add_4603_13_lut (.I0(GND_net), .I1(n14994[10]), .I2(n895), 
            .I3(n46366), .O(n14382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4862_4_lut (.I0(GND_net), .I1(n18153[1]), .I2(n271_c), 
            .I3(n46274), .O(n18082[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n10158[1]), .I2(n220_adj_4481), 
            .I3(n46485), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(\motor_state[2] ), 
            .I3(n45573), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n45573), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n45574));
    SB_CARRY add_4603_13 (.CI(n46366), .I0(n14994[10]), .I1(n895), .CO(n46367));
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(\motor_state[1] ), 
            .I3(n45572), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4482));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4603_12_lut (.I0(GND_net), .I1(n14994[9]), .I2(n822), 
            .I3(n46365), .O(n14382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_3 (.CI(n45572), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n45573));
    SB_CARRY add_4843_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n46557));
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(\motor_state[0] ), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4811_7 (.CI(n46636), .I0(n17778[4]), .I1(n481), .CO(n46637));
    SB_CARRY mult_16_add_1225_13 (.CI(n46737), .I0(n10689[10]), .I1(n877_adj_4474), 
            .CO(n46738));
    SB_CARRY add_4862_4 (.CI(n46274), .I0(n18153[1]), .I1(n271_c), .CO(n46275));
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n45572));
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n10689[9]), .I2(n804_adj_4483), 
            .I3(n46736), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_12 (.CI(n46736), .I0(n10689[9]), .I1(n804_adj_4483), 
            .CO(n46737));
    SB_LUT4 add_4710_15_lut (.I0(GND_net), .I1(n16633[12]), .I2(n1050), 
            .I3(n46556), .O(n16242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4710_14_lut (.I0(GND_net), .I1(n16633[11]), .I2(n977), 
            .I3(n46555), .O(n16242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4811_6_lut (.I0(GND_net), .I1(n17778[3]), .I2(n408), .I3(n46635), 
            .O(n17598[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[1] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_4 (.CI(n46485), .I0(n10158[1]), .I1(n220_adj_4481), 
            .CO(n46486));
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4485));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4862_3_lut (.I0(GND_net), .I1(n18153[0]), .I2(n198_adj_4486), 
            .I3(n46273), .O(n18082[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4862_3 (.CI(n46273), .I0(n18153[0]), .I1(n198_adj_4486), 
            .CO(n46274));
    SB_CARRY add_4492_3 (.CI(n46424), .I0(n12938[0]), .I1(n156_adj_4466), 
            .CO(n46425));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n10158[0]), .I2(n147_adj_4488), 
            .I3(n46484), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_14 (.CI(n46555), .I0(n16633[11]), .I1(n977), .CO(n46556));
    SB_CARRY add_4603_12 (.CI(n46365), .I0(n14994[9]), .I1(n822), .CO(n46366));
    SB_LUT4 add_4862_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_4489), 
            .I3(GND_net), .O(n18082[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4862_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4811_6 (.CI(n46635), .I0(n17778[3]), .I1(n408), .CO(n46636));
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n10689[8]), .I2(n731_adj_4490), 
            .I3(n46735), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4710_13_lut (.I0(GND_net), .I1(n16633[10]), .I2(n904), 
            .I3(n46554), .O(n16242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_11_lut (.I0(GND_net), .I1(n14994[8]), .I2(n749), 
            .I3(n46364), .O(n14382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n46735), .I0(n10689[8]), .I1(n731_adj_4490), 
            .CO(n46736));
    SB_CARRY mult_17_add_1225_3 (.CI(n46484), .I0(n10158[0]), .I1(n147_adj_4488), 
            .CO(n46485));
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4811_5_lut (.I0(GND_net), .I1(n17778[2]), .I2(n335_adj_4487), 
            .I3(n46634), .O(n17598[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4862_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_4489), .CO(n46273));
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4485), .I2(n74), 
            .I3(GND_net), .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_12_lut (.I0(GND_net), .I1(n17378[9]), .I2(n840), 
            .I3(n46272), .O(n17114[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_11_lut (.I0(GND_net), .I1(n17378[8]), .I2(n767), 
            .I3(n46271), .O(n17114[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n10689[7]), .I2(n658_adj_4482), 
            .I3(n46734), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4710_13 (.CI(n46554), .I0(n16633[10]), .I1(n904), .CO(n46555));
    SB_CARRY mult_16_add_1225_10 (.CI(n46734), .I0(n10689[7]), .I1(n658_adj_4482), 
            .CO(n46735));
    SB_CARRY add_4771_11 (.CI(n46271), .I0(n17378[8]), .I1(n767), .CO(n46272));
    SB_CARRY add_4603_11 (.CI(n46364), .I0(n14994[8]), .I1(n749), .CO(n46365));
    SB_LUT4 add_4710_12_lut (.I0(GND_net), .I1(n16633[9]), .I2(n831), 
            .I3(n46553), .O(n16242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4490));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4771_10_lut (.I0(GND_net), .I1(n17378[7]), .I2(n694), 
            .I3(n46270), .O(n17114[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4489));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4488));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_4485), .I1(n74), 
            .CO(n46484));
    SB_CARRY add_4811_5 (.CI(n46634), .I0(n17778[2]), .I1(n335_adj_4487), 
            .CO(n46635));
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4486));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4406_23_lut (.I0(GND_net), .I1(n11174[20]), .I2(GND_net), 
            .I3(n46483), .O(n10158[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n10689[6]), .I2(n585), 
            .I3(n46733), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_9 (.CI(n46733), .I0(n10689[6]), .I1(n585), 
            .CO(n46734));
    SB_LUT4 add_4492_2_lut (.I0(GND_net), .I1(n14_adj_4417), .I2(n83), 
            .I3(GND_net), .O(n12098[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_2 (.CI(GND_net), .I0(n14_adj_4417), .I1(n83), .CO(n46424));
    SB_LUT4 add_4603_10_lut (.I0(GND_net), .I1(n14994[7]), .I2(n676), 
            .I3(n46363), .O(n14382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n18202[1]), 
            .I3(n4_adj_4475), .O(n18153[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_CARRY add_4771_10 (.CI(n46270), .I0(n17378[7]), .I1(n694), .CO(n46271));
    SB_LUT4 add_4771_9_lut (.I0(GND_net), .I1(n17378[6]), .I2(n621), .I3(n46269), 
            .O(n17114[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n10689[5]), .I2(n512), 
            .I3(n46732), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4811_4_lut (.I0(GND_net), .I1(n17778[1]), .I2(n262), .I3(n46633), 
            .O(n17598[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47141_4_lut (.I0(n60519), .I1(n61865), .I2(n62947), .I3(n59936), 
            .O(n62041));   // verilog/motorControl.v(51[33:53])
    defparam i47141_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47142_3_lut (.I0(n62041), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n62042));   // verilog/motorControl.v(51[33:53])
    defparam i47142_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_4491));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46665_3_lut (.I0(n6_adj_4491), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n61565));   // verilog/motorControl.v(51[33:53])
    defparam i46665_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46666_3_lut (.I0(n61565), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n61566));   // verilog/motorControl.v(51[33:53])
    defparam i46666_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45010_4_lut (.I0(n356[21]), .I1(n62937), .I2(n382[21]), .I3(n60831), 
            .O(n59910));
    defparam i45010_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i46271_4_lut (.I0(n24_adj_4492), .I1(n8_adj_4493), .I2(n62910), 
            .I3(n59904), .O(n61171));   // verilog/motorControl.v(51[33:53])
    defparam i46271_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[14]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45617_3_lut (.I0(n61566), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n60517));   // verilog/motorControl.v(51[33:53])
    defparam i45617_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[10] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47140_3_lut (.I0(n62042), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n62040));   // verilog/motorControl.v(51[33:53])
    defparam i47140_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45016_4_lut (.I0(n356[21]), .I1(n62912), .I2(n382[21]), .I3(n62075), 
            .O(n59916));
    defparam i45016_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[15]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_21_i45_rep_92_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n62910));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i45_rep_92_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46875_4_lut (.I0(n60517), .I1(n61171), .I2(n62910), .I3(n59910), 
            .O(n61775));   // verilog/motorControl.v(51[33:53])
    defparam i46875_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45625_3_lut (.I0(n62040), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n60525));   // verilog/motorControl.v(51[33:53])
    defparam i45625_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(deadband[0]), .I1(n356[1]), .I2(deadband[1]), 
            .I3(n356[0]), .O(n4_adj_4494));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46673_3_lut (.I0(n4_adj_4494), .I1(n356[13]), .I2(n27), .I3(GND_net), 
            .O(n61573));   // verilog/motorControl.v(51[12:29])
    defparam i46673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46674_3_lut (.I0(n61573), .I1(n356[14]), .I2(n29), .I3(GND_net), 
            .O(n61574));   // verilog/motorControl.v(51[12:29])
    defparam i46674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45133_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n60043), 
            .O(n60033));
    defparam i45133_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46947_4_lut (.I0(n30), .I1(n10_adj_4413), .I2(n35_adj_4414), 
            .I3(n60029), .O(n61847));   // verilog/motorControl.v(51[12:29])
    defparam i46947_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4811_4 (.CI(n46633), .I0(n17778[1]), .I1(n262), .CO(n46634));
    SB_CARRY add_4603_10 (.CI(n46363), .I0(n14994[7]), .I1(n676), .CO(n46364));
    SB_LUT4 add_4811_3_lut (.I0(GND_net), .I1(n17778[0]), .I2(n189), .I3(n46632), 
            .O(n17598[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4811_3 (.CI(n46632), .I0(n17778[0]), .I1(n189), .CO(n46633));
    SB_CARRY add_4771_9 (.CI(n46269), .I0(n17378[6]), .I1(n621), .CO(n46270));
    SB_CARRY mult_16_add_1225_8 (.CI(n46732), .I0(n10689[5]), .I1(n512), 
            .CO(n46733));
    SB_LUT4 add_4811_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n17598[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4811_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4483));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4603_9_lut (.I0(GND_net), .I1(n14994[6]), .I2(n603), .I3(n46362), 
            .O(n14382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_8_lut (.I0(GND_net), .I1(n17378[5]), .I2(n548), .I3(n46268), 
            .O(n17114[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n10689[4]), .I2(n439), 
            .I3(n46731), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4771_8 (.CI(n46268), .I0(n17378[5]), .I1(n548), .CO(n46269));
    SB_CARRY add_4710_12 (.CI(n46553), .I0(n16633[9]), .I1(n831), .CO(n46554));
    SB_CARRY add_4811_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n46632));
    SB_LUT4 add_4586_19_lut (.I0(GND_net), .I1(n14705[16]), .I2(GND_net), 
            .I3(n46631), .O(n14058[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4771_7_lut (.I0(GND_net), .I1(n17378[4]), .I2(n475), .I3(n46267), 
            .O(n17114[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_7 (.CI(n46731), .I0(n10689[4]), .I1(n439), 
            .CO(n46732));
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n10689[3]), .I2(n366), 
            .I3(n46730), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_9 (.CI(n46362), .I0(n14994[6]), .I1(n603), .CO(n46363));
    SB_CARRY mult_16_add_1225_6 (.CI(n46730), .I0(n10689[3]), .I1(n366), 
            .CO(n46731));
    SB_LUT4 add_4586_18_lut (.I0(GND_net), .I1(n14705[15]), .I2(GND_net), 
            .I3(n46630), .O(n14058[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_18 (.CI(n46630), .I0(n14705[15]), .I1(GND_net), 
            .CO(n46631));
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4481));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45609_3_lut (.I0(n61574), .I1(n356[15]), .I2(n31), .I3(GND_net), 
            .O(n60509));   // verilog/motorControl.v(51[12:29])
    defparam i45609_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4771_7 (.CI(n46267), .I0(n17378[4]), .I1(n475), .CO(n46268));
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n10689[2]), .I2(n293_adj_4495), 
            .I3(n46729), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_5 (.CI(n46729), .I0(n10689[2]), .I1(n293_adj_4495), 
            .CO(n46730));
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n10689[1]), .I2(n220_adj_4497), 
            .I3(n46728), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_6_lut (.I0(GND_net), .I1(n17378[3]), .I2(n402_adj_4498), 
            .I3(n46266), .O(n17114[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_8_lut (.I0(GND_net), .I1(n14994[5]), .I2(n530), .I3(n46361), 
            .O(n14382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4406_22_lut (.I0(GND_net), .I1(n11174[19]), .I2(GND_net), 
            .I3(n46482), .O(n10158[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_11_lut (.I0(GND_net), .I1(n17697[8]), .I2(n770), 
            .I3(n46423), .O(n17498[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_8 (.CI(n46361), .I0(n14994[5]), .I1(n530), .CO(n46362));
    SB_CARRY add_4771_6 (.CI(n46266), .I0(n17378[3]), .I1(n402_adj_4498), 
            .CO(n46267));
    SB_LUT4 add_4710_11_lut (.I0(GND_net), .I1(n16633[8]), .I2(n758), 
            .I3(n46552), .O(n16242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_17_lut (.I0(GND_net), .I1(n14705[14]), .I2(GND_net), 
            .I3(n46629), .O(n14058[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_5_lut (.I0(GND_net), .I1(n17378[2]), .I2(n329), .I3(n46265), 
            .O(n17114[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_11 (.CI(n46552), .I0(n16633[8]), .I1(n758), .CO(n46553));
    SB_CARRY add_4586_17 (.CI(n46629), .I0(n14705[14]), .I1(GND_net), 
            .CO(n46630));
    SB_CARRY add_4406_22 (.CI(n46482), .I0(n11174[19]), .I1(GND_net), 
            .CO(n46483));
    SB_LUT4 add_4603_7_lut (.I0(GND_net), .I1(n14994[4]), .I2(n457), .I3(n46360), 
            .O(n14382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4771_5 (.CI(n46265), .I0(n17378[2]), .I1(n329), .CO(n46266));
    SB_CARRY mult_16_add_1225_4 (.CI(n46728), .I0(n10689[1]), .I1(n220_adj_4497), 
            .CO(n46729));
    SB_LUT4 add_4406_21_lut (.I0(GND_net), .I1(n11174[18]), .I2(GND_net), 
            .I3(n46481), .O(n10158[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n10689[0]), .I2(n147_adj_4499), 
            .I3(n46727), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_16_lut (.I0(GND_net), .I1(n14705[13]), .I2(n1111), 
            .I3(n46628), .O(n14058[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n46727), .I0(n10689[0]), .I1(n147_adj_4499), 
            .CO(n46728));
    SB_CARRY add_4586_16 (.CI(n46628), .I0(n14705[13]), .I1(n1111), .CO(n46629));
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4500), .I2(n74_adj_4501), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4710_10_lut (.I0(GND_net), .I1(n16633[7]), .I2(n685), 
            .I3(n46551), .O(n16242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_4_lut (.I0(GND_net), .I1(n17378[1]), .I2(n256), .I3(n46264), 
            .O(n17114[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_15_lut (.I0(GND_net), .I1(n14705[12]), .I2(n1038), 
            .I3(n46627), .O(n14058[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_10 (.CI(n46551), .I0(n16633[7]), .I1(n685), .CO(n46552));
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n10182[0]), .I2(n9651[0]), 
            .I3(n45640), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_10_lut (.I0(GND_net), .I1(n17697[7]), .I2(n697), 
            .I3(n46422), .O(n17498[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_7 (.CI(n46360), .I0(n14994[4]), .I1(n457), .CO(n46361));
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[0]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4710_9_lut (.I0(GND_net), .I1(n16633[6]), .I2(n612), .I3(n46550), 
            .O(n16242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[1]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4802_10 (.CI(n46422), .I0(n17697[7]), .I1(n697), .CO(n46423));
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5_adj_4500), .I1(n74_adj_4501), 
            .CO(n46727));
    SB_CARRY add_4771_4 (.CI(n46264), .I0(n17378[1]), .I1(n256), .CO(n46265));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n45639), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_24 (.CI(n45639), .I0(n257[22]), .I1(n306[22]), .CO(n45640));
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[2]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47208_4_lut (.I0(n60509), .I1(n61847), .I2(n35_adj_4414), 
            .I3(n60033), .O(n62108));   // verilog/motorControl.v(51[12:29])
    defparam i47208_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47209_3_lut (.I0(n62108), .I1(n356[18]), .I2(n37), .I3(GND_net), 
            .O(n62109));   // verilog/motorControl.v(51[12:29])
    defparam i47209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n45638), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[3]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[4]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n49[23]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 i47161_3_lut (.I0(n62109), .I1(n356[19]), .I2(n39), .I3(GND_net), 
            .O(n62061));   // verilog/motorControl.v(51[12:29])
    defparam i47161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4474));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[13] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[5]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4503));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i75_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n49[22]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[6]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n49[21]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n49[20]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n49[19]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n49[18]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n49[17]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n49[16]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n49[15]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n49[14]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n49[13]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n49[12]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n49[11]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n49[10]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n49[9]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n49[8]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n49[7]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n49[6]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 i45095_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n62002), 
            .O(n59995));
    defparam i45095_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4507));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4429_23_lut (.I0(GND_net), .I1(n11657[20]), .I2(GND_net), 
            .I3(n46726), .O(n10689[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_22_lut (.I0(GND_net), .I1(n11657[19]), .I2(GND_net), 
            .I3(n46725), .O(n10689[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[7]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4469));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46873_4_lut (.I0(n60507), .I1(n61169), .I2(n45), .I3(n59991), 
            .O(n61773));   // verilog/motorControl.v(51[12:29])
    defparam i46873_4_lut.LUT_INIT = 16'hccca;
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n49[5]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n49[4]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n49[3]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n49[2]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n49[1]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_23 (.CI(n45638), .I0(n257[21]), .I1(n306[21]), .CO(n45639));
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[8]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4466));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n18202[2]), .I1(n6_c), .I2(\Kp[4] ), 
            .I3(n1[18]), .O(n18153[3]));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h9666;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4957[9]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4586_15 (.CI(n46627), .I0(n14705[12]), .I1(n1038), .CO(n46628));
    SB_CARRY add_4429_22 (.CI(n46725), .I0(n11657[19]), .I1(GND_net), 
            .CO(n46726));
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n45637), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_22 (.CI(n45637), .I0(n257[20]), .I1(n306[20]), .CO(n45638));
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n45636), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_6_lut (.I0(GND_net), .I1(n14994[3]), .I2(n384_adj_4509), 
            .I3(n46359), .O(n14382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4771_3_lut (.I0(GND_net), .I1(n17378[0]), .I2(n183_adj_4510), 
            .I3(n46263), .O(n17114[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_21_lut (.I0(GND_net), .I1(n11657[18]), .I2(GND_net), 
            .I3(n46724), .O(n10689[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_21 (.CI(n46724), .I0(n11657[18]), .I1(GND_net), 
            .CO(n46725));
    SB_CARRY add_4771_3 (.CI(n46263), .I0(n17378[0]), .I1(n183_adj_4510), 
            .CO(n46264));
    SB_LUT4 add_4771_2_lut (.I0(GND_net), .I1(n41_adj_4507), .I2(n110_adj_4503), 
            .I3(GND_net), .O(n17114[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_21 (.CI(n46481), .I0(n11174[18]), .I1(GND_net), 
            .CO(n46482));
    SB_CARRY add_4771_2 (.CI(GND_net), .I0(n41_adj_4507), .I1(n110_adj_4503), 
            .CO(n46263));
    SB_CARRY add_4603_6 (.CI(n46359), .I0(n14994[3]), .I1(n384_adj_4509), 
            .CO(n46360));
    SB_LUT4 add_4802_9_lut (.I0(GND_net), .I1(n17697[6]), .I2(n624), .I3(n46421), 
            .O(n17498[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4802_9 (.CI(n46421), .I0(n17697[6]), .I1(n624), .CO(n46422));
    SB_LUT4 add_4802_8_lut (.I0(GND_net), .I1(n17697[5]), .I2(n551), .I3(n46420), 
            .O(n17498[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_20_lut (.I0(GND_net), .I1(n11657[17]), .I2(GND_net), 
            .I3(n46723), .O(n10689[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_5_lut (.I0(GND_net), .I1(n14994[2]), .I2(n311), .I3(n46358), 
            .O(n14382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_21 (.CI(n45636), .I0(n257[19]), .I1(n306[19]), .CO(n45637));
    SB_LUT4 add_4406_20_lut (.I0(GND_net), .I1(n11174[17]), .I2(GND_net), 
            .I3(n46480), .O(n10158[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n45635), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4802_8 (.CI(n46420), .I0(n17697[5]), .I1(n551), .CO(n46421));
    SB_CARRY add_4603_5 (.CI(n46358), .I0(n14994[2]), .I1(n311), .CO(n46359));
    SB_LUT4 add_4586_14_lut (.I0(GND_net), .I1(n14705[11]), .I2(n965), 
            .I3(n46626), .O(n14058[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_9 (.CI(n46550), .I0(n16633[6]), .I1(n612), .CO(n46551));
    SB_LUT4 add_4603_4_lut (.I0(GND_net), .I1(n14994[1]), .I2(n238), .I3(n46357), 
            .O(n14382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_4 (.CI(n46357), .I0(n14994[1]), .I1(n238), .CO(n46358));
    SB_CARRY add_18_20 (.CI(n45635), .I0(n257[18]), .I1(n306[18]), .CO(n45636));
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n45634), .O(n356[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_3_lut (.I0(GND_net), .I1(n14994[0]), .I2(n165), .I3(n46356), 
            .O(n14382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4710_8_lut (.I0(GND_net), .I1(n16633[5]), .I2(n539), .I3(n46549), 
            .O(n16242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_14 (.CI(n46626), .I0(n14705[11]), .I1(n965), .CO(n46627));
    SB_CARRY add_4406_20 (.CI(n46480), .I0(n11174[17]), .I1(GND_net), 
            .CO(n46481));
    SB_LUT4 i45615_3_lut (.I0(n62061), .I1(n356[20]), .I2(n41), .I3(GND_net), 
            .O(n60515));   // verilog/motorControl.v(51[12:29])
    defparam i45615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47061_4_lut (.I0(n60515), .I1(n61773), .I2(n45), .I3(n59995), 
            .O(n61961));   // verilog/motorControl.v(51[12:29])
    defparam i47061_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47063_4_lut (.I0(n60525), .I1(n61775), .I2(n62910), .I3(n59916), 
            .O(n61963));   // verilog/motorControl.v(51[33:53])
    defparam i47063_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4406_19_lut (.I0(GND_net), .I1(n11174[16]), .I2(GND_net), 
            .I3(n46479), .O(n10158[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_7_lut (.I0(GND_net), .I1(n17697[4]), .I2(n478), .I3(n46419), 
            .O(n17498[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_8 (.CI(n46549), .I0(n16633[5]), .I1(n539), .CO(n46550));
    SB_CARRY add_4603_3 (.CI(n46356), .I0(n14994[0]), .I1(n165), .CO(n46357));
    SB_CARRY add_4429_20 (.CI(n46723), .I0(n11657[17]), .I1(GND_net), 
            .CO(n46724));
    SB_LUT4 add_4586_13_lut (.I0(GND_net), .I1(n14705[10]), .I2(n892), 
            .I3(n46625), .O(n14058[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_19_lut (.I0(GND_net), .I1(n11657[16]), .I2(GND_net), 
            .I3(n46722), .O(n10689[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_19 (.CI(n46722), .I0(n11657[16]), .I1(GND_net), 
            .CO(n46723));
    SB_LUT4 i1_4_lut_adj_949 (.I0(n61961), .I1(control_update), .I2(deadband[23]), 
            .I3(n356[23]), .O(n56216));
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h4c04;
    SB_CARRY add_4406_19 (.CI(n46479), .I0(n11174[16]), .I1(GND_net), 
            .CO(n46480));
    SB_CARRY add_4802_7 (.CI(n46419), .I0(n17697[4]), .I1(n478), .CO(n46420));
    SB_LUT4 add_4603_2_lut (.I0(GND_net), .I1(n23_c), .I2(n92), .I3(GND_net), 
            .O(n14382[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n45634), .I0(n257[17]), .I1(n306[17]), .CO(n45635));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n45633), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n56216), .I1(n61963), .I2(n356[23]), 
            .I3(n47_adj_4511), .O(n55139));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h0a22;
    SB_LUT4 add_4710_7_lut (.I0(GND_net), .I1(n16633[4]), .I2(n466), .I3(n46548), 
            .O(n16242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_6_lut (.I0(GND_net), .I1(n17697[3]), .I2(n405), .I3(n46418), 
            .O(n17498[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_18 (.CI(n45633), .I0(n257[16]), .I1(n306[16]), .CO(n45634));
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n45632), .O(n356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_17 (.CI(n45632), .I0(n257[15]), .I1(n306[15]), .CO(n45633));
    SB_CARRY add_4603_2 (.CI(GND_net), .I0(n23_c), .I1(n92), .CO(n46356));
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n45631), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n45631), .I0(n257[14]), .I1(n306[14]), .CO(n45632));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n45630), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4802_6 (.CI(n46418), .I0(n17697[3]), .I1(n405), .CO(n46419));
    SB_CARRY add_18_15 (.CI(n45630), .I0(n257[13]), .I1(n306[13]), .CO(n45631));
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n45629), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_17_lut (.I0(GND_net), .I1(n15538[14]), .I2(GND_net), 
            .I3(n46355), .O(n14994[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_14 (.CI(n45629), .I0(n257[12]), .I1(n306[12]), .CO(n45630));
    SB_LUT4 add_4429_18_lut (.I0(GND_net), .I1(n11657[15]), .I2(GND_net), 
            .I3(n46721), .O(n10689[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n45628), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_5_lut (.I0(GND_net), .I1(n17697[2]), .I2(n332), .I3(n46417), 
            .O(n17498[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_13 (.CI(n45628), .I0(n257[11]), .I1(n306[11]), .CO(n45629));
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n45627), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_7 (.CI(n46548), .I0(n16633[4]), .I1(n466), .CO(n46549));
    SB_CARRY add_4802_5 (.CI(n46417), .I0(n17697[2]), .I1(n332), .CO(n46418));
    SB_LUT4 add_4710_6_lut (.I0(GND_net), .I1(n16633[3]), .I2(n393), .I3(n46547), 
            .O(n16242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4406_18_lut (.I0(GND_net), .I1(n11174[15]), .I2(GND_net), 
            .I3(n46478), .O(n10158[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_13 (.CI(n46625), .I0(n14705[10]), .I1(n892), .CO(n46626));
    SB_CARRY add_18_12 (.CI(n45627), .I0(n257[10]), .I1(n306[10]), .CO(n45628));
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n45626), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_16_lut (.I0(GND_net), .I1(n15538[13]), .I2(n1117), 
            .I3(n46354), .O(n14994[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4802_4_lut (.I0(GND_net), .I1(n17697[1]), .I2(n259), .I3(n46416), 
            .O(n17498[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_11 (.CI(n45626), .I0(n257[9]), .I1(n306[9]), .CO(n45627));
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n45625), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_16 (.CI(n46354), .I0(n15538[13]), .I1(n1117), .CO(n46355));
    SB_CARRY add_4429_18 (.CI(n46721), .I0(n11657[15]), .I1(GND_net), 
            .CO(n46722));
    SB_CARRY add_4710_6 (.CI(n46547), .I0(n16633[3]), .I1(n393), .CO(n46548));
    SB_CARRY add_18_10 (.CI(n45625), .I0(n257[8]), .I1(n306[8]), .CO(n45626));
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n45624), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_9 (.CI(n45624), .I0(n257[7]), .I1(n306[7]), .CO(n45625));
    SB_LUT4 add_4586_12_lut (.I0(GND_net), .I1(n14705[9]), .I2(n819), 
            .I3(n46624), .O(n14058[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_17_lut (.I0(GND_net), .I1(n11657[14]), .I2(GND_net), 
            .I3(n46720), .O(n10689[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4510));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n26922), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4406_18 (.CI(n46478), .I0(n11174[15]), .I1(GND_net), 
            .CO(n46479));
    SB_CARRY add_4429_17 (.CI(n46720), .I0(n11657[14]), .I1(GND_net), 
            .CO(n46721));
    SB_LUT4 add_4710_5_lut (.I0(GND_net), .I1(n16633[2]), .I2(n320), .I3(n46546), 
            .O(n16242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[8]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n27524), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n27523), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_4636_15_lut (.I0(GND_net), .I1(n15538[12]), .I2(n1044), 
            .I3(n46353), .O(n14994[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4406_17_lut (.I0(GND_net), .I1(n11174[14]), .I2(GND_net), 
            .I3(n46477), .O(n10158[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n45623), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_8 (.CI(n45623), .I0(n257[6]), .I1(n306[6]), .CO(n45624));
    SB_LUT4 add_4429_16_lut (.I0(GND_net), .I1(n11657[13]), .I2(n1099), 
            .I3(n46719), .O(n10689[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4509));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n27522), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n27521), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n27520), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFSR counter_1935__i0 (.Q(counter[0]), .C(clk16MHz), .D(n51[0]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n27519), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n27518), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n27517), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n27516), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n27515), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n27514), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4429_16 (.CI(n46719), .I0(n11657[13]), .I1(n1099), .CO(n46720));
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n27513), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4636_15 (.CI(n46353), .I0(n15538[12]), .I1(n1044), .CO(n46354));
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n45622), 
            .O(n375)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_7 (.CI(n45622), .I0(n257[5]), .I1(n306[5]), .CO(n45623));
    SB_CARRY add_4586_12 (.CI(n46624), .I0(n14705[9]), .I1(n819), .CO(n46625));
    SB_LUT4 add_4636_14_lut (.I0(GND_net), .I1(n15538[11]), .I2(n971), 
            .I3(n46352), .O(n14994[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n45621), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_6 (.CI(n45621), .I0(n257[4]), .I1(n306[4]), .CO(n45622));
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n45620), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4802_4 (.CI(n46416), .I0(n17697[1]), .I1(n259), .CO(n46417));
    SB_CARRY add_18_5 (.CI(n45620), .I0(n257[3]), .I1(n306[3]), .CO(n45621));
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n45619), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n27512), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_18_4 (.CI(n45619), .I0(n257[2]), .I1(n306[2]), .CO(n45620));
    SB_CARRY add_4710_5 (.CI(n46546), .I0(n16633[2]), .I1(n320), .CO(n46547));
    SB_LUT4 add_4710_4_lut (.I0(GND_net), .I1(n16633[1]), .I2(n247), .I3(n46545), 
            .O(n16242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_11_lut (.I0(GND_net), .I1(n14705[8]), .I2(n746), 
            .I3(n46623), .O(n14058[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n27511), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 i1_3_lut_4_lut_adj_951 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n18202[0]), 
            .I3(n45445), .O(n18153[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_951.LUT_INIT = 16'h8778;
    SB_LUT4 add_4802_3_lut (.I0(GND_net), .I1(n17697[0]), .I2(n186_adj_4514), 
            .I3(n46415), .O(n17498[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_15_lut (.I0(GND_net), .I1(n11657[12]), .I2(n1026), 
            .I3(n46718), .O(n10689[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n27510), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4429_15 (.CI(n46718), .I0(n11657[12]), .I1(n1026), .CO(n46719));
    SB_CARRY add_4586_11 (.CI(n46623), .I0(n14705[8]), .I1(n746), .CO(n46624));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n45618), 
            .O(n356[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n27509), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_4586_10_lut (.I0(GND_net), .I1(n14705[7]), .I2(n673), 
            .I3(n46622), .O(n14058[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_17 (.CI(n46477), .I0(n11174[14]), .I1(GND_net), 
            .CO(n46478));
    SB_LUT4 add_4429_14_lut (.I0(GND_net), .I1(n11657[11]), .I2(n953), 
            .I3(n46717), .O(n10689[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_10 (.CI(n46622), .I0(n14705[7]), .I1(n673), .CO(n46623));
    SB_LUT4 add_4586_9_lut (.I0(GND_net), .I1(n14705[6]), .I2(n600), .I3(n46621), 
            .O(n14058[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_4 (.CI(n46545), .I0(n16633[1]), .I1(n247), .CO(n46546));
    SB_LUT4 add_4406_16_lut (.I0(GND_net), .I1(n11174[13]), .I2(n1099_adj_4515), 
            .I3(n46476), .O(n10158[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_9 (.CI(n46621), .I0(n14705[6]), .I1(n600), .CO(n46622));
    SB_CARRY add_4802_3 (.CI(n46415), .I0(n17697[0]), .I1(n186_adj_4514), 
            .CO(n46416));
    SB_CARRY add_4636_14 (.CI(n46352), .I0(n15538[11]), .I1(n971), .CO(n46353));
    SB_LUT4 add_4710_3_lut (.I0(GND_net), .I1(n16633[0]), .I2(n174), .I3(n46544), 
            .O(n16242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n27508), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4429_14 (.CI(n46717), .I0(n11657[11]), .I1(n953), .CO(n46718));
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n27507), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_4429_13_lut (.I0(GND_net), .I1(n11657[10]), .I2(n880), 
            .I3(n46716), .O(n10689[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n27506), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_4710_3 (.CI(n46544), .I0(n16633[0]), .I1(n174), .CO(n46545));
    SB_CARRY add_4429_13 (.CI(n46716), .I0(n11657[10]), .I1(n880), .CO(n46717));
    SB_LUT4 add_4802_2_lut (.I0(GND_net), .I1(n44_adj_4516), .I2(n113_adj_4517), 
            .I3(GND_net), .O(n17498[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4802_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_3 (.CI(n45618), .I0(n257[1]), .I1(n306[1]), .CO(n45619));
    SB_LUT4 add_4429_12_lut (.I0(GND_net), .I1(n11657[9]), .I2(n807), 
            .I3(n46715), .O(n10689[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_13_lut (.I0(GND_net), .I1(n15538[10]), .I2(n898), 
            .I3(n46351), .O(n14994[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_8_lut (.I0(GND_net), .I1(n14705[5]), .I2(n527), .I3(n46620), 
            .O(n14058[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_13 (.CI(n46351), .I0(n15538[10]), .I1(n898), .CO(n46352));
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_12 (.CI(n46715), .I0(n11657[9]), .I1(n807), .CO(n46716));
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n45618));
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n1[23]), .I3(n45617), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n1[22]), .I3(n45616), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_11_lut (.I0(GND_net), .I1(n11657[8]), .I2(n734), 
            .I3(n46714), .O(n10689[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_8 (.CI(n46620), .I0(n14705[5]), .I1(n527), .CO(n46621));
    SB_CARRY add_4429_11 (.CI(n46714), .I0(n11657[8]), .I1(n734), .CO(n46715));
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n27505), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n27504), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n27503), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_4586_7_lut (.I0(GND_net), .I1(n14705[4]), .I2(n454), .I3(n46619), 
            .O(n14058[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_24 (.CI(n45616), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n1[22]), .CO(n45617));
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n27502), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n1[21]), .I3(n45615), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_10_lut (.I0(GND_net), .I1(n11657[7]), .I2(n661), 
            .I3(n46713), .O(n10689[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_10 (.CI(n46713), .I0(n11657[7]), .I1(n661), .CO(n46714));
    SB_CARRY add_9_23 (.CI(n45615), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n1[21]), .CO(n45616));
    SB_CARRY add_4802_2 (.CI(GND_net), .I0(n44_adj_4516), .I1(n113_adj_4517), 
            .CO(n46415));
    SB_LUT4 add_4636_12_lut (.I0(GND_net), .I1(n15538[9]), .I2(n825), 
            .I3(n46350), .O(n14994[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_9_lut (.I0(GND_net), .I1(n11657[6]), .I2(n588), .I3(n46712), 
            .O(n10689[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n1[20]), .I3(n45614), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4519));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4520));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4521));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4522));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4523));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4524));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4525));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4527));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4528));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4529));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4530));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4531));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4532));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4533));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4534));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4535));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4536));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4537));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44526_4_lut (.I0(n21_adj_4533), .I1(n19_adj_4537), .I2(n17_adj_4536), 
            .I3(n9_adj_4525), .O(n59426));
    defparam i44526_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45399_4_lut (.I0(n27_adj_4530), .I1(n15_adj_4535), .I2(n13_adj_4528), 
            .I3(n11_adj_4527), .O(n60299));
    defparam i45399_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_4522), 
            .I3(GND_net), .O(n12_adj_4538));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_4528), 
            .I3(GND_net), .O(n10_adj_4539));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_4538), .I1(n130[17]), .I2(n35_adj_4529), 
            .I3(GND_net), .O(n30_adj_4540));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45476_4_lut (.I0(n13_adj_4528), .I1(n11_adj_4527), .I2(n9_adj_4525), 
            .I3(n59515), .O(n60376));
    defparam i45476_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i45436_4_lut (.I0(n19_adj_4537), .I1(n17_adj_4536), .I2(n15_adj_4535), 
            .I3(n60376), .O(n60336));
    defparam i45436_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46821_4_lut (.I0(n25_adj_4534), .I1(n23), .I2(n21_adj_4533), 
            .I3(n60336), .O(n61721));
    defparam i46821_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46513_4_lut (.I0(n31_adj_4532), .I1(n29_adj_4531), .I2(n27_adj_4530), 
            .I3(n61721), .O(n61413));
    defparam i46513_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47108_4_lut (.I0(n37_adj_4523), .I1(n35_adj_4529), .I2(n33_adj_4522), 
            .I3(n61413), .O(n62008));
    defparam i47108_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_adj_4524), 
            .I3(GND_net), .O(n16_adj_4542));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46867_3_lut (.I0(n6_adj_4543), .I1(n130[10]), .I2(n21_adj_4533), 
            .I3(GND_net), .O(n61767));   // verilog/motorControl.v(45[12:34])
    defparam i46867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46868_3_lut (.I0(n61767), .I1(n143), .I2(n23), .I3(GND_net), 
            .O(n61768));   // verilog/motorControl.v(45[12:34])
    defparam i46868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_4536), 
            .I3(GND_net), .O(n8_adj_4544));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_4542), .I1(n130[22]), .I2(n45_adj_4521), 
            .I3(GND_net), .O(n24_adj_4545));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4636_12 (.CI(n46350), .I0(n15538[9]), .I1(n825), .CO(n46351));
    SB_CARRY add_9_22 (.CI(n45614), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n1[20]), .CO(n45615));
    SB_CARRY add_4429_9 (.CI(n46712), .I0(n11657[6]), .I1(n588), .CO(n46713));
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n1[19]), .I3(n45613), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45319_4_lut (.I0(n43_adj_4524), .I1(n25_adj_4534), .I2(n23), 
            .I3(n59426), .O(n60219));
    defparam i45319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4531_20_lut (.I0(GND_net), .I1(n13698[17]), .I2(GND_net), 
            .I3(n46414), .O(n12938[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_8_lut (.I0(GND_net), .I1(n11657[5]), .I2(n515), .I3(n46711), 
            .O(n10689[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_8 (.CI(n46711), .I0(n11657[5]), .I1(n515), .CO(n46712));
    SB_CARRY add_4406_16 (.CI(n46476), .I0(n11174[13]), .I1(n1099_adj_4515), 
            .CO(n46477));
    SB_LUT4 add_4531_19_lut (.I0(GND_net), .I1(n13698[16]), .I2(GND_net), 
            .I3(n46413), .O(n12938[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4710_2_lut (.I0(GND_net), .I1(n32_adj_4546), .I2(n101), 
            .I3(GND_net), .O(n16242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4710_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_7_lut (.I0(GND_net), .I1(n11657[4]), .I2(n442), .I3(n46710), 
            .O(n10689[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_7 (.CI(n46619), .I0(n14705[4]), .I1(n454), .CO(n46620));
    SB_LUT4 add_4636_11_lut (.I0(GND_net), .I1(n15538[8]), .I2(n752), 
            .I3(n46349), .O(n14994[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_7 (.CI(n46710), .I0(n11657[4]), .I1(n442), .CO(n46711));
    SB_LUT4 add_4586_6_lut (.I0(GND_net), .I1(n14705[3]), .I2(n381), .I3(n46618), 
            .O(n14058[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_6_lut (.I0(GND_net), .I1(n11657[3]), .I2(n369_adj_4547), 
            .I3(n46709), .O(n10689[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_11 (.CI(n46349), .I0(n15538[8]), .I1(n752), .CO(n46350));
    SB_CARRY add_4586_6 (.CI(n46618), .I0(n14705[3]), .I1(n381), .CO(n46619));
    SB_LUT4 i46265_4_lut (.I0(n24_adj_4545), .I1(n8_adj_4544), .I2(n45_adj_4521), 
            .I3(n60215), .O(n61165));   // verilog/motorControl.v(45[12:34])
    defparam i46265_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4636_10_lut (.I0(GND_net), .I1(n15538[7]), .I2(n679), 
            .I3(n46348), .O(n14994[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_5_lut (.I0(GND_net), .I1(n14705[2]), .I2(n308), .I3(n46617), 
            .O(n14058[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4710_2 (.CI(GND_net), .I0(n32_adj_4546), .I1(n101), .CO(n46544));
    SB_CARRY add_4429_6 (.CI(n46709), .I0(n11657[3]), .I1(n369_adj_4547), 
            .CO(n46710));
    SB_CARRY add_4586_5 (.CI(n46617), .I0(n14705[2]), .I1(n308), .CO(n46618));
    SB_LUT4 add_4429_5_lut (.I0(GND_net), .I1(n11657[2]), .I2(n296_adj_4548), 
            .I3(n46708), .O(n10689[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1935__i1 (.Q(counter[1]), .C(clk16MHz), .D(n51[1]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 i46575_3_lut (.I0(n61768), .I1(n130[12]), .I2(n25_adj_4534), 
            .I3(GND_net), .O(n61475));   // verilog/motorControl.v(45[12:34])
    defparam i46575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4586_4_lut (.I0(GND_net), .I1(n14705[1]), .I2(n235), .I3(n46616), 
            .O(n14058[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1935__i2 (.Q(counter[2]), .C(clk16MHz), .D(n51[2]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i3 (.Q(counter[3]), .C(clk16MHz), .D(n51[3]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i4 (.Q(counter[4]), .C(clk16MHz), .D(n51[4]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i5 (.Q(counter[5]), .C(clk16MHz), .D(n51[5]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i6 (.Q(counter[6]), .C(clk16MHz), .D(n51[6]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i7 (.Q(counter[7]), .C(clk16MHz), .D(n51[7]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i8 (.Q(counter[8]), .C(clk16MHz), .D(n51[8]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i9 (.Q(counter[9]), .C(clk16MHz), .D(n51[9]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i10 (.Q(counter[10]), .C(clk16MHz), .D(n51[10]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i11 (.Q(counter[11]), .C(clk16MHz), .D(n51[11]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i12 (.Q(counter[12]), .C(clk16MHz), .D(n51[12]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i13 (.Q(counter[13]), .C(clk16MHz), .D(n51[13]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i14 (.Q(counter[14]), .C(clk16MHz), .D(n51[14]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i15 (.Q(counter[15]), .C(clk16MHz), .D(n51[15]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i16 (.Q(counter[16]), .C(clk16MHz), .D(n51[16]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i17 (.Q(counter[17]), .C(clk16MHz), .D(n51[17]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i18 (.Q(counter[18]), .C(clk16MHz), .D(n51[18]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i19 (.Q(counter[19]), .C(clk16MHz), .D(n51[19]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i20 (.Q(counter[20]), .C(clk16MHz), .D(n51[20]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i21 (.Q(counter[21]), .C(clk16MHz), .D(n51[21]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i22 (.Q(counter[22]), .C(clk16MHz), .D(n51[22]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i23 (.Q(counter[23]), .C(clk16MHz), .D(n51[23]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i24 (.Q(counter[24]), .C(clk16MHz), .D(n51[24]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i25 (.Q(counter[25]), .C(clk16MHz), .D(n51[25]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i26 (.Q(counter[26]), .C(clk16MHz), .D(n51[26]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i27 (.Q(counter[27]), .C(clk16MHz), .D(n51[27]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i28 (.Q(counter[28]), .C(clk16MHz), .D(n51[28]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i29 (.Q(counter[29]), .C(clk16MHz), .D(n51[29]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i30 (.Q(counter[30]), .C(clk16MHz), .D(n51[30]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1935__i31 (.Q(counter[31]), .C(clk16MHz), .D(n51[31]), 
            .R(counter_31__N_3690));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4563));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i46687_3_lut (.I0(n4_adj_4563), .I1(n130[13]), .I2(n27_adj_4530), 
            .I3(GND_net), .O(n61587));   // verilog/motorControl.v(45[12:34])
    defparam i46687_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4586_4 (.CI(n46616), .I0(n14705[1]), .I1(n235), .CO(n46617));
    SB_CARRY add_4429_5 (.CI(n46708), .I0(n11657[2]), .I1(n296_adj_4548), 
            .CO(n46709));
    SB_LUT4 add_4586_3_lut (.I0(GND_net), .I1(n14705[0]), .I2(n162_adj_4564), 
            .I3(n46615), .O(n14058[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46688_3_lut (.I0(n61587), .I1(n130[14]), .I2(n29_adj_4531), 
            .I3(GND_net), .O(n61588));   // verilog/motorControl.v(45[12:34])
    defparam i46688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4736_14_lut (.I0(GND_net), .I1(n16970[11]), .I2(n980), 
            .I3(n46543), .O(n16633[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45382_4_lut (.I0(n33_adj_4522), .I1(n31_adj_4532), .I2(n29_adj_4531), 
            .I3(n60299), .O(n60282));
    defparam i45382_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_9_21 (.CI(n45613), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n1[19]), .CO(n45614));
    SB_CARRY add_4636_10 (.CI(n46348), .I0(n15538[7]), .I1(n679), .CO(n46349));
    SB_LUT4 add_4736_13_lut (.I0(GND_net), .I1(n16970[10]), .I2(n907), 
            .I3(n46542), .O(n16633[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_3 (.CI(n46615), .I0(n14705[0]), .I1(n162_adj_4564), 
            .CO(n46616));
    SB_LUT4 add_4406_15_lut (.I0(GND_net), .I1(n11174[12]), .I2(n1026_adj_4565), 
            .I3(n46475), .O(n10158[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_19 (.CI(n46413), .I0(n13698[16]), .I1(GND_net), 
            .CO(n46414));
    SB_LUT4 add_4429_4_lut (.I0(GND_net), .I1(n11657[1]), .I2(n223), .I3(n46707), 
            .O(n10689[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_18_lut (.I0(GND_net), .I1(n13698[15]), .I2(GND_net), 
            .I3(n46412), .O(n12938[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_4 (.CI(n46707), .I0(n11657[1]), .I1(n223), .CO(n46708));
    SB_LUT4 add_4586_2_lut (.I0(GND_net), .I1(n20_adj_4566), .I2(n89), 
            .I3(GND_net), .O(n14058[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_3_lut (.I0(GND_net), .I1(n11657[0]), .I2(n150_adj_4567), 
            .I3(n46706), .O(n10689[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_9_lut (.I0(GND_net), .I1(n15538[6]), .I2(n606), .I3(n46347), 
            .O(n14994[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_9 (.CI(n46347), .I0(n15538[6]), .I1(n606), .CO(n46348));
    SB_CARRY add_4429_3 (.CI(n46706), .I0(n11657[0]), .I1(n150_adj_4567), 
            .CO(n46707));
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n1[18]), .I3(n45612), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_2_lut (.I0(GND_net), .I1(n8_adj_4568), .I2(n77), 
            .I3(GND_net), .O(n10689[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_2 (.CI(GND_net), .I0(n8_adj_4568), .I1(n77), .CO(n46706));
    SB_LUT4 add_4472_22_lut (.I0(GND_net), .I1(n12538[19]), .I2(GND_net), 
            .I3(n46705), .O(n11657[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_2 (.CI(GND_net), .I0(n20_adj_4566), .I1(n89), .CO(n46615));
    SB_LUT4 add_4472_21_lut (.I0(GND_net), .I1(n12538[18]), .I2(GND_net), 
            .I3(n46704), .O(n11657[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_13 (.CI(n46542), .I0(n16970[10]), .I1(n907), .CO(n46543));
    SB_CARRY add_9_20 (.CI(n45612), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n1[18]), .CO(n45613));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n1[17]), .I3(n45611), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n45611), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n1[17]), .CO(n45612));
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n1[16]), .I3(n45610), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_8_lut (.I0(GND_net), .I1(n15538[5]), .I2(n533), .I3(n46346), 
            .O(n14994[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4736_12_lut (.I0(GND_net), .I1(n16970[9]), .I2(n834), 
            .I3(n46541), .O(n16633[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_18 (.CI(n45610), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n1[16]), .CO(n45611));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n1[15]), .I3(n45609), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n53137), .I1(\data_in_frame[9][6] ), .I2(\data_in_frame[11][3] ), 
            .I3(Kp_23__N_969), .O(n22_adj_4569));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n53140), .I1(Kp_23__N_645), .I2(\data_in_frame[11][4] ), 
            .I3(\data_in_frame[12][3] ), .O(n24_adj_4570));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4636_8 (.CI(n46346), .I0(n15538[5]), .I1(n533), .CO(n46347));
    SB_LUT4 i46941_4_lut (.I0(n30_adj_4540), .I1(n10_adj_4539), .I2(n35_adj_4529), 
            .I3(n60277), .O(n61841));   // verilog/motorControl.v(45[12:34])
    defparam i46941_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i9_4_lut (.I0(n23958), .I1(\data_in_frame[12][5] ), .I2(n23338), 
            .I3(\data_in_frame[12][1] ), .O(n23_adj_4571));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_9_17 (.CI(n45609), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n1[15]), .CO(n45610));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n1[14]), .I3(n45608), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_16 (.CI(n45608), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n1[14]), .CO(n45609));
    SB_LUT4 add_4636_7_lut (.I0(GND_net), .I1(n15538[4]), .I2(n460), .I3(n46345), 
            .O(n14994[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_952 (.I0(Kp_23__N_675), .I1(n25_adj_4572), .I2(n23_adj_4571), 
            .I3(n24_adj_4570), .O(n10_adj_4573));
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_CARRY add_4531_18 (.CI(n46412), .I0(n13698[15]), .I1(GND_net), 
            .CO(n46413));
    SB_CARRY add_4472_21 (.CI(n46704), .I0(n12538[18]), .I1(GND_net), 
            .CO(n46705));
    SB_LUT4 add_4531_17_lut (.I0(GND_net), .I1(n13698[14]), .I2(GND_net), 
            .I3(n46411), .O(n12938[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_15 (.CI(n46475), .I0(n11174[12]), .I1(n1026_adj_4565), 
            .CO(n46476));
    SB_LUT4 add_4620_18_lut (.I0(GND_net), .I1(n15282[15]), .I2(GND_net), 
            .I3(n46614), .O(n14705[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_20_lut (.I0(GND_net), .I1(n12538[17]), .I2(GND_net), 
            .I3(n46703), .O(n11657[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n1[13]), .I3(n45607), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_17_lut (.I0(GND_net), .I1(n15282[14]), .I2(GND_net), 
            .I3(n46613), .O(n14705[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_20 (.CI(n46703), .I0(n12538[17]), .I1(GND_net), 
            .CO(n46704));
    SB_LUT4 add_4472_19_lut (.I0(GND_net), .I1(n12538[16]), .I2(GND_net), 
            .I3(n46702), .O(n11657[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_17 (.CI(n46613), .I0(n15282[14]), .I1(GND_net), 
            .CO(n46614));
    SB_CARRY add_9_15 (.CI(n45607), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n1[13]), .CO(n45608));
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n1[12]), .I3(n45606), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_7 (.CI(n46345), .I0(n15538[4]), .I1(n460), .CO(n46346));
    SB_LUT4 add_4406_14_lut (.I0(GND_net), .I1(n11174[11]), .I2(n953_adj_4574), 
            .I3(n46474), .O(n10158[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_19 (.CI(n46702), .I0(n12538[16]), .I1(GND_net), 
            .CO(n46703));
    SB_CARRY add_4736_12 (.CI(n46541), .I0(n16970[9]), .I1(n834), .CO(n46542));
    SB_LUT4 add_4636_6_lut (.I0(GND_net), .I1(n15538[3]), .I2(n387_adj_4575), 
            .I3(n46344), .O(n14994[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_14 (.CI(n45606), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n1[12]), .CO(n45607));
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n1[11]), .I3(n45605), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n45605), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n1[11]), .CO(n45606));
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n1[10]), .I3(n45604), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_12 (.CI(n45604), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n1[10]), .CO(n45605));
    SB_LUT4 add_4620_16_lut (.I0(GND_net), .I1(n15282[13]), .I2(n1114_adj_4576), 
            .I3(n46612), .O(n14705[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_6 (.CI(n46344), .I0(n15538[3]), .I1(n387_adj_4575), 
            .CO(n46345));
    SB_LUT4 add_4736_11_lut (.I0(GND_net), .I1(n16970[8]), .I2(n761), 
            .I3(n46540), .O(n16633[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n1[9]), .I3(n45603), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(n52656), .I1(n52455), .I2(n52831), .I3(n10_adj_4573), 
            .O(n16_adj_4577));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_9_11 (.CI(n45603), .I0(\PID_CONTROLLER.integral [9]), .I1(n1[9]), 
            .CO(n45604));
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n1[8]), .I3(n45602), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_18_lut (.I0(GND_net), .I1(n12538[15]), .I2(GND_net), 
            .I3(n46701), .O(n11657[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45589_3_lut (.I0(n61588), .I1(n130[15]), .I2(n31_adj_4532), 
            .I3(GND_net), .O(n60489));   // verilog/motorControl.v(45[12:34])
    defparam i45589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4472_18 (.CI(n46701), .I0(n12538[15]), .I1(GND_net), 
            .CO(n46702));
    SB_LUT4 add_4472_17_lut (.I0(GND_net), .I1(n12538[14]), .I2(GND_net), 
            .I3(n46700), .O(n11657[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47204_4_lut (.I0(n60489), .I1(n61841), .I2(n35_adj_4529), 
            .I3(n60282), .O(n62104));   // verilog/motorControl.v(45[12:34])
    defparam i47204_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47205_3_lut (.I0(n62104), .I1(n130[18]), .I2(n37_adj_4523), 
            .I3(GND_net), .O(n62105));   // verilog/motorControl.v(45[12:34])
    defparam i47205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_953 (.I0(n52848), .I1(n16_adj_4577), .I2(n12_adj_4578), 
            .I3(n52925), .O(n22568));
    defparam i8_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_CARRY add_4472_17 (.CI(n46700), .I0(n12538[14]), .I1(GND_net), 
            .CO(n46701));
    SB_CARRY add_4620_16 (.CI(n46612), .I0(n15282[13]), .I1(n1114_adj_4576), 
            .CO(n46613));
    SB_LUT4 add_4620_15_lut (.I0(GND_net), .I1(n15282[12]), .I2(n1041_adj_4579), 
            .I3(n46611), .O(n14705[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_11 (.CI(n46540), .I0(n16970[8]), .I1(n761), .CO(n46541));
    SB_CARRY add_4406_14 (.CI(n46474), .I0(n11174[11]), .I1(n953_adj_4574), 
            .CO(n46475));
    SB_CARRY add_4531_17 (.CI(n46411), .I0(n13698[14]), .I1(GND_net), 
            .CO(n46412));
    SB_LUT4 add_4472_16_lut (.I0(GND_net), .I1(n12538[13]), .I2(n1102), 
            .I3(n46699), .O(n11657[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4636_5_lut (.I0(GND_net), .I1(n15538[2]), .I2(n314), .I3(n46343), 
            .O(n14994[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4736_10_lut (.I0(GND_net), .I1(n16970[7]), .I2(n688), 
            .I3(n46539), .O(n16633[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_10 (.CI(n45602), .I0(\PID_CONTROLLER.integral [8]), .I1(n1[8]), 
            .CO(n45603));
    SB_CARRY add_4472_16 (.CI(n46699), .I0(n12538[13]), .I1(n1102), .CO(n46700));
    SB_LUT4 add_4472_15_lut (.I0(GND_net), .I1(n12538[12]), .I2(n1029), 
            .I3(n46698), .O(n11657[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_5 (.CI(n46343), .I0(n15538[2]), .I1(n314), .CO(n46344));
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n1[7]), .I3(n45601), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_15 (.CI(n46698), .I0(n12538[12]), .I1(n1029), .CO(n46699));
    SB_LUT4 add_4636_4_lut (.I0(GND_net), .I1(n15538[1]), .I2(n241), .I3(n46342), 
            .O(n14994[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_10 (.CI(n46539), .I0(n16970[7]), .I1(n688), .CO(n46540));
    SB_LUT4 add_4472_14_lut (.I0(GND_net), .I1(n12538[11]), .I2(n956), 
            .I3(n46697), .O(n11657[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n45601), .I0(\PID_CONTROLLER.integral [7]), .I1(n1[7]), 
            .CO(n45602));
    SB_CARRY add_4472_14 (.CI(n46697), .I0(n12538[11]), .I1(n956), .CO(n46698));
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n1[6]), .I3(n45600), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4736_9_lut (.I0(GND_net), .I1(n16970[6]), .I2(n615), .I3(n46538), 
            .O(n16633[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_8 (.CI(n45600), .I0(\PID_CONTROLLER.integral [6]), .I1(n1[6]), 
            .CO(n45601));
    SB_LUT4 add_4472_13_lut (.I0(GND_net), .I1(n12538[10]), .I2(n883), 
            .I3(n46696), .O(n11657[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_16_lut (.I0(GND_net), .I1(n13698[13]), .I2(n1108), 
            .I3(n46410), .O(n12938[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n1[5]), .I3(n45599), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_7 (.CI(n45599), .I0(\PID_CONTROLLER.integral [5]), .I1(n1[5]), 
            .CO(n45600));
    SB_CARRY add_4636_4 (.CI(n46342), .I0(n15538[1]), .I1(n241), .CO(n46343));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n1[4]), .I3(n45598), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n45598), .I0(\PID_CONTROLLER.integral [4]), .I1(n1[4]), 
            .CO(n45599));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n1[3]), .I3(n45597), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_16 (.CI(n46410), .I0(n13698[13]), .I1(n1108), .CO(n46411));
    SB_CARRY add_4620_15 (.CI(n46611), .I0(n15282[12]), .I1(n1041_adj_4579), 
            .CO(n46612));
    SB_CARRY add_4736_9 (.CI(n46538), .I0(n16970[6]), .I1(n615), .CO(n46539));
    SB_LUT4 add_4531_15_lut (.I0(GND_net), .I1(n13698[12]), .I2(n1035), 
            .I3(n46409), .O(n12938[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_13 (.CI(n46696), .I0(n12538[10]), .I1(n883), .CO(n46697));
    SB_CARRY add_9_5 (.CI(n45597), .I0(\PID_CONTROLLER.integral [3]), .I1(n1[3]), 
            .CO(n45598));
    SB_LUT4 add_4736_8_lut (.I0(GND_net), .I1(n16970[5]), .I2(n542), .I3(n46537), 
            .O(n16633[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_12_lut (.I0(GND_net), .I1(n12538[9]), .I2(n810), 
            .I3(n46695), .O(n11657[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_14_lut (.I0(GND_net), .I1(n15282[11]), .I2(n968_adj_4581), 
            .I3(n46610), .O(n14705[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_12 (.CI(n46695), .I0(n12538[9]), .I1(n810), .CO(n46696));
    SB_LUT4 add_4636_3_lut (.I0(GND_net), .I1(n15538[0]), .I2(n168), .I3(n46341), 
            .O(n14994[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_11_lut (.I0(GND_net), .I1(n12538[8]), .I2(n737), 
            .I3(n46694), .O(n11657[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_11 (.CI(n46694), .I0(n12538[8]), .I1(n737), .CO(n46695));
    SB_CARRY add_4620_14 (.CI(n46610), .I0(n15282[11]), .I1(n968_adj_4581), 
            .CO(n46611));
    SB_LUT4 add_4406_13_lut (.I0(GND_net), .I1(n11174[10]), .I2(n880_adj_4582), 
            .I3(n46473), .O(n10158[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_15 (.CI(n46409), .I0(n13698[12]), .I1(n1035), .CO(n46410));
    SB_LUT4 add_4472_10_lut (.I0(GND_net), .I1(n12538[7]), .I2(n664), 
            .I3(n46693), .O(n11657[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_13_lut (.I0(GND_net), .I1(n15282[10]), .I2(n895_adj_4583), 
            .I3(n46609), .O(n14705[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n1[2]), .I3(n45596), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4636_3 (.CI(n46341), .I0(n15538[0]), .I1(n168), .CO(n46342));
    SB_CARRY add_4406_13 (.CI(n46473), .I0(n11174[10]), .I1(n880_adj_4582), 
            .CO(n46474));
    SB_LUT4 add_4406_12_lut (.I0(GND_net), .I1(n11174[9]), .I2(n807_adj_4585), 
            .I3(n46472), .O(n10158[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_10 (.CI(n46693), .I0(n12538[7]), .I1(n664), .CO(n46694));
    SB_CARRY add_4620_13 (.CI(n46609), .I0(n15282[10]), .I1(n895_adj_4583), 
            .CO(n46610));
    SB_LUT4 add_4531_14_lut (.I0(GND_net), .I1(n13698[11]), .I2(n962), 
            .I3(n46408), .O(n12938[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_12_lut (.I0(GND_net), .I1(n15282[9]), .I2(n822_adj_4586), 
            .I3(n46608), .O(n14705[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47168_3_lut (.I0(n62105), .I1(n130[19]), .I2(n39_adj_4520), 
            .I3(GND_net), .O(n62068));   // verilog/motorControl.v(45[12:34])
    defparam i47168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4636_2_lut (.I0(GND_net), .I1(n26_adj_4587), .I2(n95), 
            .I3(GND_net), .O(n14994[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4636_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_4 (.CI(n45596), .I0(\PID_CONTROLLER.integral [2]), .I1(n1[2]), 
            .CO(n45597));
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n1[1]), .I3(n45595), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_3 (.CI(n45595), .I0(\PID_CONTROLLER.integral [1]), .I1(n1[1]), 
            .CO(n45596));
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n1[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45323_4_lut (.I0(n43_adj_4524), .I1(n41_adj_4519), .I2(n39_adj_4520), 
            .I3(n62008), .O(n60223));
    defparam i45323_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4736_8 (.CI(n46537), .I0(n16970[5]), .I1(n542), .CO(n46538));
    SB_CARRY add_4636_2 (.CI(GND_net), .I0(n26_adj_4587), .I1(n95), .CO(n46341));
    SB_CARRY add_4531_14 (.CI(n46408), .I0(n13698[11]), .I1(n962), .CO(n46409));
    SB_LUT4 add_4736_7_lut (.I0(GND_net), .I1(n16970[4]), .I2(n469), .I3(n46536), 
            .O(n16633[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4836_9_lut (.I0(GND_net), .I1(n17985[6]), .I2(n630), .I3(n46340), 
            .O(n17858[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n1[0]), 
            .CO(n45595));
    SB_LUT4 i46869_4_lut (.I0(n61475), .I1(n61165), .I2(n45_adj_4521), 
            .I3(n60219), .O(n61769));   // verilog/motorControl.v(45[12:34])
    defparam i46869_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4472_9_lut (.I0(GND_net), .I1(n12538[6]), .I2(n591), .I3(n46692), 
            .O(n11657[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_12 (.CI(n46608), .I0(n15282[9]), .I1(n822_adj_4586), 
            .CO(n46609));
    SB_CARRY add_4736_7 (.CI(n46536), .I0(n16970[4]), .I1(n469), .CO(n46537));
    SB_LUT4 add_4620_11_lut (.I0(GND_net), .I1(n15282[8]), .I2(n749_adj_4588), 
            .I3(n46607), .O(n14705[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_9 (.CI(n46692), .I0(n12538[6]), .I1(n591), .CO(n46693));
    SB_LUT4 add_4531_13_lut (.I0(GND_net), .I1(n13698[10]), .I2(n889), 
            .I3(n46407), .O(n12938[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4836_8_lut (.I0(GND_net), .I1(n17985[5]), .I2(n557), .I3(n46339), 
            .O(n17858[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_13 (.CI(n46407), .I0(n13698[10]), .I1(n889), .CO(n46408));
    SB_CARRY add_4620_11 (.CI(n46607), .I0(n15282[8]), .I1(n749_adj_4588), 
            .CO(n46608));
    SB_CARRY add_4406_12 (.CI(n46472), .I0(n11174[9]), .I1(n807_adj_4585), 
            .CO(n46473));
    SB_LUT4 i45595_3_lut (.I0(n62068), .I1(n130[20]), .I2(n41_adj_4519), 
            .I3(GND_net), .O(n60495));   // verilog/motorControl.v(45[12:34])
    defparam i45595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4736_6_lut (.I0(GND_net), .I1(n16970[3]), .I2(n396_adj_4589), 
            .I3(n46535), .O(n16633[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_8_lut (.I0(GND_net), .I1(n12538[5]), .I2(n518), .I3(n46691), 
            .O(n11657[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_8 (.CI(n46691), .I0(n12538[5]), .I1(n518), .CO(n46692));
    SB_LUT4 add_4620_10_lut (.I0(GND_net), .I1(n15282[7]), .I2(n676_adj_4590), 
            .I3(n46606), .O(n14705[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_10 (.CI(n46606), .I0(n15282[7]), .I1(n676_adj_4590), 
            .CO(n46607));
    SB_LUT4 add_4472_7_lut (.I0(GND_net), .I1(n12538[4]), .I2(n445), .I3(n46690), 
            .O(n11657[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_7 (.CI(n46690), .I0(n12538[4]), .I1(n445), .CO(n46691));
    SB_LUT4 add_4406_11_lut (.I0(GND_net), .I1(n11174[8]), .I2(n734_adj_4591), 
            .I3(n46471), .O(n10158[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_6_lut (.I0(GND_net), .I1(n12538[3]), .I2(n372_adj_4592), 
            .I3(n46689), .O(n11657[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_9_lut (.I0(GND_net), .I1(n15282[6]), .I2(n603_adj_4593), 
            .I3(n46605), .O(n14705[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_11 (.CI(n46471), .I0(n11174[8]), .I1(n734_adj_4591), 
            .CO(n46472));
    SB_CARRY add_4472_6 (.CI(n46689), .I0(n12538[3]), .I1(n372_adj_4592), 
            .CO(n46690));
    SB_CARRY add_4836_8 (.CI(n46339), .I0(n17985[5]), .I1(n557), .CO(n46340));
    SB_LUT4 add_4472_5_lut (.I0(GND_net), .I1(n12538[2]), .I2(n299_adj_4594), 
            .I3(n46688), .O(n11657[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47057_4_lut (.I0(n60495), .I1(n61769), .I2(n45_adj_4521), 
            .I3(n60223), .O(n61957));   // verilog/motorControl.v(45[12:34])
    defparam i47057_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4836_7_lut (.I0(GND_net), .I1(n17985[4]), .I2(n484), .I3(n46338), 
            .O(n17858[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47058_3_lut (.I0(n61957), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(45[12:34])
    defparam i47058_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4472_5 (.CI(n46688), .I0(n12538[2]), .I1(n299_adj_4594), 
            .CO(n46689));
    SB_CARRY add_4620_9 (.CI(n46605), .I0(n15282[6]), .I1(n603_adj_4593), 
            .CO(n46606));
    SB_CARRY add_4736_6 (.CI(n46535), .I0(n16970[3]), .I1(n396_adj_4589), 
            .CO(n46536));
    SB_LUT4 add_4531_12_lut (.I0(GND_net), .I1(n13698[9]), .I2(n816), 
            .I3(n46406), .O(n12938[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4472_4_lut (.I0(GND_net), .I1(n12538[1]), .I2(n226), .I3(n46687), 
            .O(n11657[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4836_7 (.CI(n46338), .I0(n17985[4]), .I1(n484), .CO(n46339));
    SB_CARRY add_4472_4 (.CI(n46687), .I0(n12538[1]), .I1(n226), .CO(n46688));
    SB_LUT4 add_4472_3_lut (.I0(GND_net), .I1(n12538[0]), .I2(n153_adj_4595), 
            .I3(n46686), .O(n11657[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4596));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4620_8_lut (.I0(GND_net), .I1(n15282[5]), .I2(n530_adj_4597), 
            .I3(n46604), .O(n14705[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4736_5_lut (.I0(GND_net), .I1(n16970[2]), .I2(n323), .I3(n46534), 
            .O(n16633[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_5 (.CI(n46534), .I0(n16970[2]), .I1(n323), .CO(n46535));
    SB_CARRY add_4620_8 (.CI(n46604), .I0(n15282[5]), .I1(n530_adj_4597), 
            .CO(n46605));
    SB_LUT4 add_4406_10_lut (.I0(GND_net), .I1(n11174[7]), .I2(n661_adj_4598), 
            .I3(n46470), .O(n10158[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4472_3 (.CI(n46686), .I0(n12538[0]), .I1(n153_adj_4595), 
            .CO(n46687));
    SB_LUT4 add_4620_7_lut (.I0(GND_net), .I1(n15282[4]), .I2(n457_adj_4599), 
            .I3(n46603), .O(n14705[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_12 (.CI(n46406), .I0(n13698[9]), .I1(n816), .CO(n46407));
    SB_LUT4 add_4836_6_lut (.I0(GND_net), .I1(n17985[3]), .I2(n411), .I3(n46337), 
            .O(n17858[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_7 (.CI(n46603), .I0(n15282[4]), .I1(n457_adj_4599), 
            .CO(n46604));
    SB_LUT4 add_4531_11_lut (.I0(GND_net), .I1(n13698[8]), .I2(n743), 
            .I3(n46405), .O(n12938[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4836_6 (.CI(n46337), .I0(n17985[3]), .I1(n411), .CO(n46338));
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4600));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4531_11 (.CI(n46405), .I0(n13698[8]), .I1(n743), .CO(n46406));
    SB_LUT4 add_4472_2_lut (.I0(GND_net), .I1(n11_adj_4601), .I2(n80), 
            .I3(GND_net), .O(n11657[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4472_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4836_5_lut (.I0(GND_net), .I1(n17985[2]), .I2(n338_adj_4602), 
            .I3(n46336), .O(n17858[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_6_lut (.I0(GND_net), .I1(n15282[3]), .I2(n384_adj_4603), 
            .I3(n46602), .O(n14705[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_10 (.CI(n46470), .I0(n11174[7]), .I1(n661_adj_4598), 
            .CO(n46471));
    SB_LUT4 add_4531_10_lut (.I0(GND_net), .I1(n13698[7]), .I2(n670), 
            .I3(n46404), .O(n12938[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4836_5 (.CI(n46336), .I0(n17985[2]), .I1(n338_adj_4602), 
            .CO(n46337));
    SB_CARRY add_4472_2 (.CI(GND_net), .I0(n11_adj_4601), .I1(n80), .CO(n46686));
    SB_LUT4 add_4406_9_lut (.I0(GND_net), .I1(n11174[6]), .I2(n588_adj_4604), 
            .I3(n46469), .O(n10158[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4836_4_lut (.I0(GND_net), .I1(n17985[1]), .I2(n265), .I3(n46335), 
            .O(n17858[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4736_4_lut (.I0(GND_net), .I1(n16970[1]), .I2(n250), .I3(n46533), 
            .O(n16633[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_10 (.CI(n46404), .I0(n13698[7]), .I1(n670), .CO(n46405));
    SB_CARRY add_4836_4 (.CI(n46335), .I0(n17985[1]), .I1(n265), .CO(n46336));
    SB_LUT4 add_4792_11_lut (.I0(GND_net), .I1(n17598[8]), .I2(n770_adj_4605), 
            .I3(n46685), .O(n17378[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_9 (.CI(n46469), .I0(n11174[6]), .I1(n588_adj_4604), 
            .CO(n46470));
    SB_LUT4 add_4792_10_lut (.I0(GND_net), .I1(n17598[7]), .I2(n697_adj_4606), 
            .I3(n46684), .O(n17378[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4792_10 (.CI(n46684), .I0(n17598[7]), .I1(n697_adj_4606), 
            .CO(n46685));
    SB_LUT4 add_4792_9_lut (.I0(GND_net), .I1(n17598[6]), .I2(n624_adj_4607), 
            .I3(n46683), .O(n17378[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4836_3_lut (.I0(GND_net), .I1(n17985[0]), .I2(n192_adj_4608), 
            .I3(n46334), .O(n17858[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_9_lut (.I0(GND_net), .I1(n13698[6]), .I2(n597), .I3(n46403), 
            .O(n12938[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_4 (.CI(n46533), .I0(n16970[1]), .I1(n250), .CO(n46534));
    SB_LUT4 add_4406_8_lut (.I0(GND_net), .I1(n11174[5]), .I2(n515_adj_4609), 
            .I3(n46468), .O(n10158[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_9 (.CI(n46403), .I0(n13698[6]), .I1(n597), .CO(n46404));
    SB_CARRY add_4836_3 (.CI(n46334), .I0(n17985[0]), .I1(n192_adj_4608), 
            .CO(n46335));
    SB_CARRY add_4792_9 (.CI(n46683), .I0(n17598[6]), .I1(n624_adj_4607), 
            .CO(n46684));
    SB_CARRY add_4620_6 (.CI(n46602), .I0(n15282[3]), .I1(n384_adj_4603), 
            .CO(n46603));
    SB_LUT4 add_4531_8_lut (.I0(GND_net), .I1(n13698[5]), .I2(n524_adj_4610), 
            .I3(n46402), .O(n12938[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4611));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4612));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4736_3_lut (.I0(GND_net), .I1(n16970[0]), .I2(n177_adj_4613), 
            .I3(n46532), .O(n16633[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_5_lut (.I0(GND_net), .I1(n15282[2]), .I2(n311_adj_4614), 
            .I3(n46601), .O(n14705[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4736_3 (.CI(n46532), .I0(n16970[0]), .I1(n177_adj_4613), 
            .CO(n46533));
    SB_LUT4 add_4792_8_lut (.I0(GND_net), .I1(n17598[5]), .I2(n551_adj_4615), 
            .I3(n46682), .O(n17378[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_5 (.CI(n46601), .I0(n15282[2]), .I1(n311_adj_4614), 
            .CO(n46602));
    SB_CARRY add_4792_8 (.CI(n46682), .I0(n17598[5]), .I1(n551_adj_4615), 
            .CO(n46683));
    SB_LUT4 add_4836_2_lut (.I0(GND_net), .I1(n50_adj_4616), .I2(n119_adj_4617), 
            .I3(GND_net), .O(n17858[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4836_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4792_7_lut (.I0(GND_net), .I1(n17598[4]), .I2(n478_adj_4618), 
            .I3(n46681), .O(n17378[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4792_7 (.CI(n46681), .I0(n17598[4]), .I1(n478_adj_4618), 
            .CO(n46682));
    SB_CARRY add_4406_8 (.CI(n46468), .I0(n11174[5]), .I1(n515_adj_4609), 
            .CO(n46469));
    SB_LUT4 add_4406_7_lut (.I0(GND_net), .I1(n11174[4]), .I2(n442_adj_4619), 
            .I3(n46467), .O(n10158[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4836_2 (.CI(GND_net), .I0(n50_adj_4616), .I1(n119_adj_4617), 
            .CO(n46334));
    SB_LUT4 add_4736_2_lut (.I0(GND_net), .I1(n35_adj_4620), .I2(n104_adj_4621), 
            .I3(GND_net), .O(n16633[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4736_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4792_6_lut (.I0(GND_net), .I1(n17598[3]), .I2(n405_adj_4622), 
            .I3(n46680), .O(n17378[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4792_6 (.CI(n46680), .I0(n17598[3]), .I1(n405_adj_4622), 
            .CO(n46681));
    SB_CARRY add_4736_2 (.CI(GND_net), .I0(n35_adj_4620), .I1(n104_adj_4621), 
            .CO(n46532));
    SB_CARRY add_4531_8 (.CI(n46402), .I0(n13698[5]), .I1(n524_adj_4610), 
            .CO(n46403));
    SB_LUT4 add_4620_4_lut (.I0(GND_net), .I1(n15282[1]), .I2(n238_adj_4623), 
            .I3(n46600), .O(n14705[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_16_lut (.I0(GND_net), .I1(n16018[13]), .I2(n1120), 
            .I3(n46333), .O(n15538[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_4 (.CI(n46600), .I0(n15282[1]), .I1(n238_adj_4623), 
            .CO(n46601));
    SB_LUT4 add_4667_15_lut (.I0(GND_net), .I1(n16018[12]), .I2(n1047), 
            .I3(n46332), .O(n15538[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4620_3_lut (.I0(GND_net), .I1(n15282[0]), .I2(n165_adj_4624), 
            .I3(n46599), .O(n14705[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4792_5_lut (.I0(GND_net), .I1(n17598[2]), .I2(n332_adj_4625), 
            .I3(n46679), .O(n17378[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4856_7_lut (.I0(GND_net), .I1(n55037), .I2(n490), .I3(n46531), 
            .O(n18034[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4792_5 (.CI(n46679), .I0(n17598[2]), .I1(n332_adj_4625), 
            .CO(n46680));
    SB_LUT4 add_4531_7_lut (.I0(GND_net), .I1(n13698[4]), .I2(n451_adj_4627), 
            .I3(n46401), .O(n12938[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4792_4_lut (.I0(GND_net), .I1(n17598[1]), .I2(n259_adj_4628), 
            .I3(n46678), .O(n17378[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4620_3 (.CI(n46599), .I0(n15282[0]), .I1(n165_adj_4624), 
            .CO(n46600));
    SB_LUT4 add_4620_2_lut (.I0(GND_net), .I1(n23_adj_4629), .I2(n92_adj_4630), 
            .I3(GND_net), .O(n14705[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4620_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4792_4 (.CI(n46678), .I0(n17598[1]), .I1(n259_adj_4628), 
            .CO(n46679));
    SB_CARRY add_4620_2 (.CI(GND_net), .I0(n23_adj_4629), .I1(n92_adj_4630), 
            .CO(n46599));
    SB_LUT4 add_4856_6_lut (.I0(GND_net), .I1(n18118[3]), .I2(n417), .I3(n46530), 
            .O(n18034[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4828_9_lut (.I0(GND_net), .I1(n17922[6]), .I2(n630_adj_4632), 
            .I3(n46598), .O(n17778[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4856_6 (.CI(n46530), .I0(n18118[3]), .I1(n417), .CO(n46531));
    SB_LUT4 add_4792_3_lut (.I0(GND_net), .I1(n17598[0]), .I2(n186_adj_4633), 
            .I3(n46677), .O(n17378[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4828_8_lut (.I0(GND_net), .I1(n17922[5]), .I2(n557_adj_4634), 
            .I3(n46597), .O(n17778[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4828_8 (.CI(n46597), .I0(n17922[5]), .I1(n557_adj_4634), 
            .CO(n46598));
    SB_CARRY add_4792_3 (.CI(n46677), .I0(n17598[0]), .I1(n186_adj_4633), 
            .CO(n46678));
    SB_LUT4 add_4828_7_lut (.I0(GND_net), .I1(n17922[4]), .I2(n484_adj_4635), 
            .I3(n46596), .O(n17778[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4856_5_lut (.I0(GND_net), .I1(n18118[2]), .I2(n344), .I3(n46529), 
            .O(n18034[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4828_7 (.CI(n46596), .I0(n17922[4]), .I1(n484_adj_4635), 
            .CO(n46597));
    SB_CARRY add_4856_5 (.CI(n46529), .I0(n18118[2]), .I1(n344), .CO(n46530));
    SB_LUT4 add_4792_2_lut (.I0(GND_net), .I1(n44_adj_4637), .I2(n113_adj_4638), 
            .I3(GND_net), .O(n17378[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4792_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4828_6_lut (.I0(GND_net), .I1(n17922[3]), .I2(n411_adj_4639), 
            .I3(n46595), .O(n17778[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4856_4_lut (.I0(GND_net), .I1(n18118[1]), .I2(n271), .I3(n46528), 
            .O(n18034[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_7 (.CI(n46467), .I0(n11174[4]), .I1(n442_adj_4619), 
            .CO(n46468));
    SB_CARRY add_4828_6 (.CI(n46595), .I0(n17922[3]), .I1(n411_adj_4639), 
            .CO(n46596));
    SB_CARRY add_4856_4 (.CI(n46528), .I0(n18118[1]), .I1(n271), .CO(n46529));
    SB_LUT4 add_4406_6_lut (.I0(GND_net), .I1(n11174[3]), .I2(n369_adj_4641), 
            .I3(n46466), .O(n10158[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_6 (.CI(n46466), .I0(n11174[3]), .I1(n369_adj_4641), 
            .CO(n46467));
    SB_CARRY add_4792_2 (.CI(GND_net), .I0(n44_adj_4637), .I1(n113_adj_4638), 
            .CO(n46677));
    SB_LUT4 add_4828_5_lut (.I0(GND_net), .I1(n17922[2]), .I2(n338_adj_4642), 
            .I3(n46594), .O(n17778[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4856_3_lut (.I0(GND_net), .I1(n18118[0]), .I2(n198), .I3(n46527), 
            .O(n18034[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4406_5_lut (.I0(GND_net), .I1(n11174[2]), .I2(n296_adj_4644), 
            .I3(n46465), .O(n10158[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_5 (.CI(n46465), .I0(n11174[2]), .I1(n296_adj_4644), 
            .CO(n46466));
    SB_CARRY add_4856_3 (.CI(n46527), .I0(n18118[0]), .I1(n198), .CO(n46528));
    SB_CARRY add_4828_5 (.CI(n46594), .I0(n17922[2]), .I1(n338_adj_4642), 
            .CO(n46595));
    SB_LUT4 add_4856_2_lut (.I0(GND_net), .I1(n56_adj_4645), .I2(n125), 
            .I3(GND_net), .O(n18034[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4856_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4406_4_lut (.I0(GND_net), .I1(n11174[1]), .I2(n223_adj_4647), 
            .I3(n46464), .O(n10158[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4856_2 (.CI(GND_net), .I0(n56_adj_4645), .I1(n125), .CO(n46527));
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4648));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4512_21_lut (.I0(GND_net), .I1(n13337[18]), .I2(GND_net), 
            .I3(n46676), .O(n12538[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4828_4_lut (.I0(GND_net), .I1(n17922[1]), .I2(n265_adj_4649), 
            .I3(n46593), .O(n17778[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_20_lut (.I0(GND_net), .I1(n13337[17]), .I2(GND_net), 
            .I3(n46675), .O(n12538[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_20 (.CI(n46675), .I0(n13337[17]), .I1(GND_net), 
            .CO(n46676));
    SB_LUT4 add_4512_19_lut (.I0(GND_net), .I1(n13337[16]), .I2(GND_net), 
            .I3(n46674), .O(n12538[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_13_lut (.I0(GND_net), .I1(n17257[10]), .I2(n910_adj_4650), 
            .I3(n46526), .O(n16970[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_15 (.CI(n46332), .I0(n16018[12]), .I1(n1047), .CO(n46333));
    SB_LUT4 add_4667_14_lut (.I0(GND_net), .I1(n16018[11]), .I2(n974), 
            .I3(n46331), .O(n15538[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_14 (.CI(n46331), .I0(n16018[11]), .I1(n974), .CO(n46332));
    SB_CARRY add_4531_7 (.CI(n46401), .I0(n13698[4]), .I1(n451_adj_4627), 
            .CO(n46402));
    SB_LUT4 add_4760_12_lut (.I0(GND_net), .I1(n17257[9]), .I2(n837_adj_4651), 
            .I3(n46525), .O(n16970[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4828_4 (.CI(n46593), .I0(n17922[1]), .I1(n265_adj_4649), 
            .CO(n46594));
    SB_CARRY add_4760_12 (.CI(n46525), .I0(n17257[9]), .I1(n837_adj_4651), 
            .CO(n46526));
    SB_LUT4 add_4667_13_lut (.I0(GND_net), .I1(n16018[10]), .I2(n901), 
            .I3(n46330), .O(n15538[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_6_lut (.I0(GND_net), .I1(n13698[3]), .I2(n378_adj_4652), 
            .I3(n46400), .O(n12938[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_13 (.CI(n46330), .I0(n16018[10]), .I1(n901), .CO(n46331));
    SB_LUT4 add_4667_12_lut (.I0(GND_net), .I1(n16018[9]), .I2(n828), 
            .I3(n46329), .O(n15538[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_6 (.CI(n46400), .I0(n13698[3]), .I1(n378_adj_4652), 
            .CO(n46401));
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4653));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4828_3_lut (.I0(GND_net), .I1(n17922[0]), .I2(n192_adj_4654), 
            .I3(n46592), .O(n17778[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_19 (.CI(n46674), .I0(n13337[16]), .I1(GND_net), 
            .CO(n46675));
    SB_LUT4 add_4760_11_lut (.I0(GND_net), .I1(n17257[8]), .I2(n764_adj_4655), 
            .I3(n46524), .O(n16970[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4828_3 (.CI(n46592), .I0(n17922[0]), .I1(n192_adj_4654), 
            .CO(n46593));
    SB_LUT4 add_4512_18_lut (.I0(GND_net), .I1(n13337[15]), .I2(GND_net), 
            .I3(n46673), .O(n12538[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_5_lut (.I0(GND_net), .I1(n13698[2]), .I2(n305_adj_4656), 
            .I3(n46399), .O(n12938[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4760_11 (.CI(n46524), .I0(n17257[8]), .I1(n764_adj_4655), 
            .CO(n46525));
    SB_LUT4 add_4828_2_lut (.I0(GND_net), .I1(n50_adj_4657), .I2(n119_adj_4658), 
            .I3(GND_net), .O(n17778[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4828_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_5 (.CI(n46399), .I0(n13698[2]), .I1(n305_adj_4656), 
            .CO(n46400));
    SB_LUT4 add_4531_4_lut (.I0(GND_net), .I1(n13698[1]), .I2(n232_adj_4659), 
            .I3(n46398), .O(n12938[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_10_lut (.I0(GND_net), .I1(n17257[7]), .I2(n691_adj_4660), 
            .I3(n46523), .O(n16970[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4828_2 (.CI(GND_net), .I0(n50_adj_4657), .I1(n119_adj_4658), 
            .CO(n46592));
    SB_CARRY add_4512_18 (.CI(n46673), .I0(n13337[15]), .I1(GND_net), 
            .CO(n46674));
    SB_CARRY add_4760_10 (.CI(n46523), .I0(n17257[7]), .I1(n691_adj_4660), 
            .CO(n46524));
    SB_CARRY add_4406_4 (.CI(n46464), .I0(n11174[1]), .I1(n223_adj_4647), 
            .CO(n46465));
    SB_CARRY add_4667_12 (.CI(n46329), .I0(n16018[9]), .I1(n828), .CO(n46330));
    SB_LUT4 add_4406_3_lut (.I0(GND_net), .I1(n11174[0]), .I2(n150_adj_4661), 
            .I3(n46463), .O(n10158[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_17_lut (.I0(GND_net), .I1(n13337[14]), .I2(GND_net), 
            .I3(n46672), .O(n12538[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_17_lut (.I0(GND_net), .I1(n15793[14]), .I2(GND_net), 
            .I3(n46591), .O(n15282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_9_lut (.I0(GND_net), .I1(n17257[6]), .I2(n618_adj_4662), 
            .I3(n46522), .O(n16970[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_3 (.CI(n46463), .I0(n11174[0]), .I1(n150_adj_4661), 
            .CO(n46464));
    SB_CARRY add_4760_9 (.CI(n46522), .I0(n17257[6]), .I1(n618_adj_4662), 
            .CO(n46523));
    SB_LUT4 add_4406_2_lut (.I0(GND_net), .I1(n8_adj_4663), .I2(n77_adj_4664), 
            .I3(GND_net), .O(n10158[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4406_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_16_lut (.I0(GND_net), .I1(n15793[13]), .I2(n1117_adj_4665), 
            .I3(n46590), .O(n15282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_8_lut (.I0(GND_net), .I1(n17257[5]), .I2(n545_adj_4666), 
            .I3(n46521), .O(n16970[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4406_2 (.CI(GND_net), .I0(n8_adj_4663), .I1(n77_adj_4664), 
            .CO(n46463));
    SB_CARRY add_4760_8 (.CI(n46521), .I0(n17257[5]), .I1(n545_adj_4666), 
            .CO(n46522));
    SB_LUT4 add_4451_22_lut (.I0(GND_net), .I1(n12098[19]), .I2(GND_net), 
            .I3(n46462), .O(n11174[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_17 (.CI(n46672), .I0(n13337[14]), .I1(GND_net), 
            .CO(n46673));
    SB_CARRY add_4652_16 (.CI(n46590), .I0(n15793[13]), .I1(n1117_adj_4665), 
            .CO(n46591));
    SB_LUT4 add_4760_7_lut (.I0(GND_net), .I1(n17257[4]), .I2(n472_adj_4667), 
            .I3(n46520), .O(n16970[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_21_lut (.I0(GND_net), .I1(n12098[18]), .I2(GND_net), 
            .I3(n46461), .O(n11174[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4760_7 (.CI(n46520), .I0(n17257[4]), .I1(n472_adj_4667), 
            .CO(n46521));
    SB_CARRY add_4451_21 (.CI(n46461), .I0(n12098[18]), .I1(GND_net), 
            .CO(n46462));
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4668));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4652_15_lut (.I0(GND_net), .I1(n15793[12]), .I2(n1044_adj_4669), 
            .I3(n46589), .O(n15282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_6_lut (.I0(GND_net), .I1(n17257[3]), .I2(n399_adj_4670), 
            .I3(n46519), .O(n16970[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_20_lut (.I0(GND_net), .I1(n12098[17]), .I2(GND_net), 
            .I3(n46460), .O(n11174[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4760_6 (.CI(n46519), .I0(n17257[3]), .I1(n399_adj_4670), 
            .CO(n46520));
    SB_CARRY add_4451_20 (.CI(n46460), .I0(n12098[17]), .I1(GND_net), 
            .CO(n46461));
    SB_LUT4 add_4512_16_lut (.I0(GND_net), .I1(n13337[13]), .I2(n1105), 
            .I3(n46671), .O(n12538[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_15 (.CI(n46589), .I0(n15793[12]), .I1(n1044_adj_4669), 
            .CO(n46590));
    SB_LUT4 add_4760_5_lut (.I0(GND_net), .I1(n17257[2]), .I2(n326_adj_4671), 
            .I3(n46518), .O(n16970[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_19_lut (.I0(GND_net), .I1(n12098[16]), .I2(GND_net), 
            .I3(n46459), .O(n11174[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_19 (.CI(n46459), .I0(n12098[16]), .I1(GND_net), 
            .CO(n46460));
    SB_CARRY add_4531_4 (.CI(n46398), .I0(n13698[1]), .I1(n232_adj_4659), 
            .CO(n46399));
    SB_LUT4 add_4667_11_lut (.I0(GND_net), .I1(n16018[8]), .I2(n755), 
            .I3(n46328), .O(n15538[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_11 (.CI(n46328), .I0(n16018[8]), .I1(n755), .CO(n46329));
    SB_LUT4 add_4531_3_lut (.I0(GND_net), .I1(n13698[0]), .I2(n159_adj_4672), 
            .I3(n46397), .O(n12938[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_10_lut (.I0(GND_net), .I1(n16018[7]), .I2(n682), 
            .I3(n46327), .O(n15538[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_10 (.CI(n46327), .I0(n16018[7]), .I1(n682), .CO(n46328));
    SB_CARRY add_4760_5 (.CI(n46518), .I0(n17257[2]), .I1(n326_adj_4671), 
            .CO(n46519));
    SB_LUT4 add_4451_18_lut (.I0(GND_net), .I1(n12098[15]), .I2(GND_net), 
            .I3(n46458), .O(n11174[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_18 (.CI(n46458), .I0(n12098[15]), .I1(GND_net), 
            .CO(n46459));
    SB_CARRY add_4531_3 (.CI(n46397), .I0(n13698[0]), .I1(n159_adj_4672), 
            .CO(n46398));
    SB_LUT4 add_4667_9_lut (.I0(GND_net), .I1(n16018[6]), .I2(n609), .I3(n46326), 
            .O(n15538[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4531_2_lut (.I0(GND_net), .I1(n17_adj_4673), .I2(n86_adj_4674), 
            .I3(GND_net), .O(n12938[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4531_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_9 (.CI(n46326), .I0(n16018[6]), .I1(n609), .CO(n46327));
    SB_LUT4 add_4667_8_lut (.I0(GND_net), .I1(n16018[5]), .I2(n536), .I3(n46325), 
            .O(n15538[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4531_2 (.CI(GND_net), .I0(n17_adj_4673), .I1(n86_adj_4674), 
            .CO(n46397));
    SB_CARRY add_4667_8 (.CI(n46325), .I0(n16018[5]), .I1(n536), .CO(n46326));
    SB_LUT4 add_4667_7_lut (.I0(GND_net), .I1(n16018[4]), .I2(n463), .I3(n46324), 
            .O(n15538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_14_lut (.I0(GND_net), .I1(n15793[11]), .I2(n971_adj_4675), 
            .I3(n46588), .O(n15282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_7 (.CI(n46324), .I0(n16018[4]), .I1(n463), .CO(n46325));
    SB_CARRY add_4652_14 (.CI(n46588), .I0(n15793[11]), .I1(n971_adj_4675), 
            .CO(n46589));
    SB_LUT4 add_4760_4_lut (.I0(GND_net), .I1(n17257[1]), .I2(n253_adj_4676), 
            .I3(n46517), .O(n16970[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_17_lut (.I0(GND_net), .I1(n12098[14]), .I2(GND_net), 
            .I3(n46457), .O(n11174[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_17 (.CI(n46457), .I0(n12098[14]), .I1(GND_net), 
            .CO(n46458));
    SB_LUT4 add_4568_19_lut (.I0(GND_net), .I1(n14382[16]), .I2(GND_net), 
            .I3(n46396), .O(n13698[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_6_lut (.I0(GND_net), .I1(n16018[3]), .I2(n390_adj_4677), 
            .I3(n46323), .O(n15538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_6 (.CI(n46323), .I0(n16018[3]), .I1(n390_adj_4677), 
            .CO(n46324));
    SB_LUT4 add_4568_18_lut (.I0(GND_net), .I1(n14382[15]), .I2(GND_net), 
            .I3(n46395), .O(n13698[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_5_lut (.I0(GND_net), .I1(n16018[2]), .I2(n317), .I3(n46322), 
            .O(n15538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_5 (.CI(n46322), .I0(n16018[2]), .I1(n317), .CO(n46323));
    SB_CARRY add_4760_4 (.CI(n46517), .I0(n17257[1]), .I1(n253_adj_4676), 
            .CO(n46518));
    SB_LUT4 add_4451_16_lut (.I0(GND_net), .I1(n12098[13]), .I2(n1102_adj_4678), 
            .I3(n46456), .O(n11174[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_16 (.CI(n46456), .I0(n12098[13]), .I1(n1102_adj_4678), 
            .CO(n46457));
    SB_CARRY add_4568_18 (.CI(n46395), .I0(n14382[15]), .I1(GND_net), 
            .CO(n46396));
    SB_LUT4 add_4667_4_lut (.I0(GND_net), .I1(n16018[1]), .I2(n244), .I3(n46321), 
            .O(n15538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_4 (.CI(n46321), .I0(n16018[1]), .I1(n244), .CO(n46322));
    SB_LUT4 add_4568_17_lut (.I0(GND_net), .I1(n14382[14]), .I2(GND_net), 
            .I3(n46394), .O(n13698[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4667_3_lut (.I0(GND_net), .I1(n16018[0]), .I2(n171), .I3(n46320), 
            .O(n15538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4667_3 (.CI(n46320), .I0(n16018[0]), .I1(n171), .CO(n46321));
    SB_CARRY add_4512_16 (.CI(n46671), .I0(n13337[13]), .I1(n1105), .CO(n46672));
    SB_LUT4 add_4652_13_lut (.I0(GND_net), .I1(n15793[10]), .I2(n898_adj_4679), 
            .I3(n46587), .O(n15282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4760_3_lut (.I0(GND_net), .I1(n17257[0]), .I2(n180_adj_4680), 
            .I3(n46516), .O(n16970[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_15_lut (.I0(GND_net), .I1(n12098[12]), .I2(n1029_adj_4681), 
            .I3(n46455), .O(n11174[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_15 (.CI(n46455), .I0(n12098[12]), .I1(n1029_adj_4681), 
            .CO(n46456));
    SB_CARRY add_4568_17 (.CI(n46394), .I0(n14382[14]), .I1(GND_net), 
            .CO(n46395));
    SB_LUT4 add_4667_2_lut (.I0(GND_net), .I1(n29_adj_4682), .I2(n98), 
            .I3(GND_net), .O(n15538[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4667_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4683));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4667_2 (.CI(GND_net), .I0(n29_adj_4682), .I1(n98), .CO(n46320));
    SB_LUT4 add_4568_16_lut (.I0(GND_net), .I1(n14382[13]), .I2(n1111_adj_4684), 
            .I3(n46393), .O(n13698[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_15_lut (.I0(GND_net), .I1(n16438[12]), .I2(n1050_adj_4685), 
            .I3(n46319), .O(n16018[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_14_lut (.I0(GND_net), .I1(n16438[11]), .I2(n977_adj_4686), 
            .I3(n46318), .O(n16018[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4760_3 (.CI(n46516), .I0(n17257[0]), .I1(n180_adj_4680), 
            .CO(n46517));
    SB_LUT4 add_4451_14_lut (.I0(GND_net), .I1(n12098[11]), .I2(n956_adj_4687), 
            .I3(n46454), .O(n11174[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_16 (.CI(n46393), .I0(n14382[13]), .I1(n1111_adj_4684), 
            .CO(n46394));
    SB_CARRY add_4696_14 (.CI(n46318), .I0(n16438[11]), .I1(n977_adj_4686), 
            .CO(n46319));
    SB_LUT4 add_4696_13_lut (.I0(GND_net), .I1(n16438[10]), .I2(n904_adj_4688), 
            .I3(n46317), .O(n16018[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4568_15_lut (.I0(GND_net), .I1(n14382[12]), .I2(n1038_adj_4689), 
            .I3(n46392), .O(n13698[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_13 (.CI(n46317), .I0(n16438[10]), .I1(n904_adj_4688), 
            .CO(n46318));
    SB_LUT4 add_4696_12_lut (.I0(GND_net), .I1(n16438[9]), .I2(n831_adj_4690), 
            .I3(n46316), .O(n16018[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_13 (.CI(n46587), .I0(n15793[10]), .I1(n898_adj_4679), 
            .CO(n46588));
    SB_LUT4 add_4760_2_lut (.I0(GND_net), .I1(n38_adj_4691), .I2(n107_adj_4692), 
            .I3(GND_net), .O(n16970[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4760_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_14 (.CI(n46454), .I0(n12098[11]), .I1(n956_adj_4687), 
            .CO(n46455));
    SB_LUT4 add_4451_13_lut (.I0(GND_net), .I1(n12098[10]), .I2(n883_adj_4693), 
            .I3(n46453), .O(n11174[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_15 (.CI(n46392), .I0(n14382[12]), .I1(n1038_adj_4689), 
            .CO(n46393));
    SB_LUT4 add_4568_14_lut (.I0(GND_net), .I1(n14382[11]), .I2(n965_adj_4694), 
            .I3(n46391), .O(n13698[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_12 (.CI(n46316), .I0(n16438[9]), .I1(n831_adj_4690), 
            .CO(n46317));
    SB_LUT4 add_4696_11_lut (.I0(GND_net), .I1(n16438[8]), .I2(n758_adj_4695), 
            .I3(n46315), .O(n16018[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_15_lut (.I0(GND_net), .I1(n13337[12]), .I2(n1032), 
            .I3(n46670), .O(n12538[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_11 (.CI(n46315), .I0(n16438[8]), .I1(n758_adj_4695), 
            .CO(n46316));
    SB_LUT4 add_4696_10_lut (.I0(GND_net), .I1(n16438[7]), .I2(n685_adj_4696), 
            .I3(n46314), .O(n16018[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_14 (.CI(n46391), .I0(n14382[11]), .I1(n965_adj_4694), 
            .CO(n46392));
    SB_CARRY add_4696_10 (.CI(n46314), .I0(n16438[7]), .I1(n685_adj_4696), 
            .CO(n46315));
    SB_CARRY add_4760_2 (.CI(GND_net), .I0(n38_adj_4691), .I1(n107_adj_4692), 
            .CO(n46516));
    SB_CARRY add_4451_13 (.CI(n46453), .I0(n12098[10]), .I1(n883_adj_4693), 
            .CO(n46454));
    SB_LUT4 add_4568_13_lut (.I0(GND_net), .I1(n14382[10]), .I2(n892_adj_4697), 
            .I3(n46390), .O(n13698[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_9_lut (.I0(GND_net), .I1(n16438[6]), .I2(n612_adj_4698), 
            .I3(n46313), .O(n16018[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_9 (.CI(n46313), .I0(n16438[6]), .I1(n612_adj_4698), 
            .CO(n46314));
    SB_LUT4 add_4782_12_lut (.I0(GND_net), .I1(n17498[9]), .I2(n840_adj_4699), 
            .I3(n46515), .O(n17257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_12_lut (.I0(GND_net), .I1(n12098[9]), .I2(n810_adj_4700), 
            .I3(n46452), .O(n11174[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_13 (.CI(n46390), .I0(n14382[10]), .I1(n892_adj_4697), 
            .CO(n46391));
    SB_LUT4 add_4696_8_lut (.I0(GND_net), .I1(n16438[5]), .I2(n539_adj_4701), 
            .I3(n46312), .O(n16018[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_8 (.CI(n46312), .I0(n16438[5]), .I1(n539_adj_4701), 
            .CO(n46313));
    SB_LUT4 add_4568_12_lut (.I0(GND_net), .I1(n14382[9]), .I2(n819_adj_4702), 
            .I3(n46389), .O(n13698[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_7_lut (.I0(GND_net), .I1(n16438[4]), .I2(n466_adj_4703), 
            .I3(n46311), .O(n16018[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_7 (.CI(n46311), .I0(n16438[4]), .I1(n466_adj_4703), 
            .CO(n46312));
    SB_CARRY add_4512_15 (.CI(n46670), .I0(n13337[12]), .I1(n1032), .CO(n46671));
    SB_LUT4 add_4652_12_lut (.I0(GND_net), .I1(n15793[9]), .I2(n825_adj_4704), 
            .I3(n46586), .O(n15282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_11_lut (.I0(GND_net), .I1(n17498[8]), .I2(n767_adj_4705), 
            .I3(n46514), .O(n17257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_12 (.CI(n46452), .I0(n12098[9]), .I1(n810_adj_4700), 
            .CO(n46453));
    SB_CARRY add_4782_11 (.CI(n46514), .I0(n17498[8]), .I1(n767_adj_4705), 
            .CO(n46515));
    SB_CARRY add_4652_12 (.CI(n46586), .I0(n15793[9]), .I1(n825_adj_4704), 
            .CO(n46587));
    SB_LUT4 add_4782_10_lut (.I0(GND_net), .I1(n17498[7]), .I2(n694_adj_4706), 
            .I3(n46513), .O(n17257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_11_lut (.I0(GND_net), .I1(n12098[8]), .I2(n737_adj_4707), 
            .I3(n46451), .O(n11174[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_10 (.CI(n46513), .I0(n17498[7]), .I1(n694_adj_4706), 
            .CO(n46514));
    SB_LUT4 add_4512_14_lut (.I0(GND_net), .I1(n13337[11]), .I2(n959_adj_4708), 
            .I3(n46669), .O(n12538[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_11_lut (.I0(GND_net), .I1(n15793[8]), .I2(n752_adj_4709), 
            .I3(n46585), .O(n15282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_11 (.CI(n46585), .I0(n15793[8]), .I1(n752_adj_4709), 
            .CO(n46586));
    SB_LUT4 add_4782_9_lut (.I0(GND_net), .I1(n17498[6]), .I2(n621_adj_4710), 
            .I3(n46512), .O(n17257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_9 (.CI(n46512), .I0(n17498[6]), .I1(n621_adj_4710), 
            .CO(n46513));
    SB_LUT4 add_4652_10_lut (.I0(GND_net), .I1(n15793[7]), .I2(n679_adj_4711), 
            .I3(n46584), .O(n15282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_8_lut (.I0(GND_net), .I1(n17498[5]), .I2(n548_adj_4712), 
            .I3(n46511), .O(n17257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_12 (.CI(n46389), .I0(n14382[9]), .I1(n819_adj_4702), 
            .CO(n46390));
    SB_LUT4 add_4696_6_lut (.I0(GND_net), .I1(n16438[3]), .I2(n393_adj_4713), 
            .I3(n46310), .O(n16018[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_8 (.CI(n46511), .I0(n17498[5]), .I1(n548_adj_4712), 
            .CO(n46512));
    SB_LUT4 add_4568_11_lut (.I0(GND_net), .I1(n14382[8]), .I2(n746_adj_4714), 
            .I3(n46388), .O(n13698[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_6 (.CI(n46310), .I0(n16438[3]), .I1(n393_adj_4713), 
            .CO(n46311));
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n143), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4715));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4716));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4512_14 (.CI(n46669), .I0(n13337[11]), .I1(n959_adj_4708), 
            .CO(n46670));
    SB_CARRY add_4652_10 (.CI(n46584), .I0(n15793[7]), .I1(n679_adj_4711), 
            .CO(n46585));
    SB_LUT4 add_4782_7_lut (.I0(GND_net), .I1(n17498[4]), .I2(n475_adj_4717), 
            .I3(n46510), .O(n17257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_11 (.CI(n46451), .I0(n12098[8]), .I1(n737_adj_4707), 
            .CO(n46452));
    SB_CARRY add_4568_11 (.CI(n46388), .I0(n14382[8]), .I1(n746_adj_4714), 
            .CO(n46389));
    SB_LUT4 add_4696_5_lut (.I0(GND_net), .I1(n16438[2]), .I2(n320_adj_4718), 
            .I3(n46309), .O(n16018[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_5 (.CI(n46309), .I0(n16438[2]), .I1(n320_adj_4718), 
            .CO(n46310));
    SB_LUT4 add_4568_10_lut (.I0(GND_net), .I1(n14382[7]), .I2(n673_adj_4719), 
            .I3(n46387), .O(n13698[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_4_lut (.I0(GND_net), .I1(n16438[1]), .I2(n247_adj_4720), 
            .I3(n46308), .O(n16018[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_4 (.CI(n46308), .I0(n16438[1]), .I1(n247_adj_4720), 
            .CO(n46309));
    SB_CARRY add_4782_7 (.CI(n46510), .I0(n17498[4]), .I1(n475_adj_4717), 
            .CO(n46511));
    SB_LUT4 add_4451_10_lut (.I0(GND_net), .I1(n12098[7]), .I2(n664_adj_4721), 
            .I3(n46450), .O(n11174[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_10 (.CI(n46387), .I0(n14382[7]), .I1(n673_adj_4719), 
            .CO(n46388));
    SB_LUT4 add_4696_3_lut (.I0(GND_net), .I1(n16438[0]), .I2(n174_adj_4722), 
            .I3(n46307), .O(n16018[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_3 (.CI(n46307), .I0(n16438[0]), .I1(n174_adj_4722), 
            .CO(n46308));
    SB_LUT4 add_4568_9_lut (.I0(GND_net), .I1(n14382[6]), .I2(n600_adj_4723), 
            .I3(n46386), .O(n13698[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4696_2_lut (.I0(GND_net), .I1(n32_adj_4724), .I2(n101_adj_4725), 
            .I3(GND_net), .O(n16018[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4696_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4696_2 (.CI(GND_net), .I0(n32_adj_4724), .I1(n101_adj_4725), 
            .CO(n46307));
    SB_LUT4 add_4652_9_lut (.I0(GND_net), .I1(n15793[6]), .I2(n606_adj_4726), 
            .I3(n46583), .O(n15282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4782_6_lut (.I0(GND_net), .I1(n17498[3]), .I2(n402_adj_4727), 
            .I3(n46509), .O(n17257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_9 (.CI(n46386), .I0(n14382[6]), .I1(n600_adj_4723), 
            .CO(n46387));
    SB_LUT4 add_4850_8_lut (.I0(GND_net), .I1(n18082[5]), .I2(n560), .I3(n46306), 
            .O(n17985[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_10 (.CI(n46450), .I0(n12098[7]), .I1(n664_adj_4721), 
            .CO(n46451));
    SB_LUT4 add_4568_8_lut (.I0(GND_net), .I1(n14382[5]), .I2(n527_adj_4728), 
            .I3(n46385), .O(n13698[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_7_lut (.I0(GND_net), .I1(n18082[4]), .I2(n487_adj_4729), 
            .I3(n46305), .O(n17985[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_7 (.CI(n46305), .I0(n18082[4]), .I1(n487_adj_4729), 
            .CO(n46306));
    SB_CARRY add_4568_8 (.CI(n46385), .I0(n14382[5]), .I1(n527_adj_4728), 
            .CO(n46386));
    SB_LUT4 add_4850_6_lut (.I0(GND_net), .I1(n18082[3]), .I2(n414_adj_4730), 
            .I3(n46304), .O(n17985[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_6 (.CI(n46304), .I0(n18082[3]), .I1(n414_adj_4730), 
            .CO(n46305));
    SB_CARRY add_4782_6 (.CI(n46509), .I0(n17498[3]), .I1(n402_adj_4727), 
            .CO(n46510));
    SB_LUT4 add_4568_7_lut (.I0(GND_net), .I1(n14382[4]), .I2(n454_adj_4731), 
            .I3(n46384), .O(n13698[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_9_lut (.I0(GND_net), .I1(n12098[6]), .I2(n591_adj_4732), 
            .I3(n46449), .O(n11174[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_7 (.CI(n46384), .I0(n14382[4]), .I1(n454_adj_4731), 
            .CO(n46385));
    SB_LUT4 add_4850_5_lut (.I0(GND_net), .I1(n18082[2]), .I2(n341_adj_4733), 
            .I3(n46303), .O(n17985[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_5 (.CI(n46303), .I0(n18082[2]), .I1(n341_adj_4733), 
            .CO(n46304));
    SB_LUT4 add_4568_6_lut (.I0(GND_net), .I1(n14382[3]), .I2(n381_adj_4734), 
            .I3(n46383), .O(n13698[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_4_lut (.I0(GND_net), .I1(n18082[1]), .I2(n268_adj_4735), 
            .I3(n46302), .O(n17985[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_4 (.CI(n46302), .I0(n18082[1]), .I1(n268_adj_4735), 
            .CO(n46303));
    SB_LUT4 add_4512_13_lut (.I0(GND_net), .I1(n13337[10]), .I2(n886_adj_4736), 
            .I3(n46668), .O(n12538[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_9 (.CI(n46583), .I0(n15793[6]), .I1(n606_adj_4726), 
            .CO(n46584));
    SB_LUT4 add_4782_5_lut (.I0(GND_net), .I1(n17498[2]), .I2(n329_adj_4737), 
            .I3(n46508), .O(n17257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_9 (.CI(n46449), .I0(n12098[6]), .I1(n591_adj_4732), 
            .CO(n46450));
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n45594), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_3_lut (.I0(GND_net), .I1(n18082[0]), .I2(n195_adj_4738), 
            .I3(n46301), .O(n17985[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_6 (.CI(n46383), .I0(n14382[3]), .I1(n381_adj_4734), 
            .CO(n46384));
    SB_CARRY add_4850_3 (.CI(n46301), .I0(n18082[0]), .I1(n195_adj_4738), 
            .CO(n46302));
    SB_LUT4 add_4850_2_lut (.I0(GND_net), .I1(n53_adj_4739), .I2(n122_adj_4740), 
            .I3(GND_net), .O(n17985[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4568_5_lut (.I0(GND_net), .I1(n14382[2]), .I2(n308_adj_4741), 
            .I3(n46382), .O(n13698[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_2 (.CI(GND_net), .I0(n53_adj_4739), .I1(n122_adj_4740), 
            .CO(n46301));
    SB_LUT4 add_4723_14_lut (.I0(GND_net), .I1(n16802[11]), .I2(n980_adj_4742), 
            .I3(n46300), .O(n16438[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_5 (.CI(n46508), .I0(n17498[2]), .I1(n329_adj_4737), 
            .CO(n46509));
    SB_LUT4 add_4451_8_lut (.I0(GND_net), .I1(n12098[5]), .I2(n518_adj_4743), 
            .I3(n46448), .O(n11174[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_5 (.CI(n46382), .I0(n14382[2]), .I1(n308_adj_4741), 
            .CO(n46383));
    SB_LUT4 add_4723_13_lut (.I0(GND_net), .I1(n16802[10]), .I2(n907_adj_4744), 
            .I3(n46299), .O(n16438[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_13 (.CI(n46299), .I0(n16802[10]), .I1(n907_adj_4744), 
            .CO(n46300));
    SB_CARRY add_4512_13 (.CI(n46668), .I0(n13337[10]), .I1(n886_adj_4736), 
            .CO(n46669));
    SB_LUT4 add_4512_12_lut (.I0(GND_net), .I1(n13337[9]), .I2(n813_adj_4745), 
            .I3(n46667), .O(n12538[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_8_lut (.I0(GND_net), .I1(n15793[5]), .I2(n533_adj_4746), 
            .I3(n46582), .O(n15282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_8 (.CI(n46582), .I0(n15793[5]), .I1(n533_adj_4746), 
            .CO(n46583));
    SB_CARRY add_4512_12 (.CI(n46667), .I0(n13337[9]), .I1(n813_adj_4745), 
            .CO(n46668));
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[23]), 
            .I3(n45740), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_7_lut (.I0(GND_net), .I1(n15793[4]), .I2(n460_adj_4748), 
            .I3(n46581), .O(n15282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4568_4_lut (.I0(GND_net), .I1(n14382[1]), .I2(n235_adj_4749), 
            .I3(n46381), .O(n13698[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4723_12_lut (.I0(GND_net), .I1(n16802[9]), .I2(n834_adj_4750), 
            .I3(n46298), .O(n16438[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_12 (.CI(n46298), .I0(n16802[9]), .I1(n834_adj_4750), 
            .CO(n46299));
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[22]), 
            .I3(n45739), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n45739), .I0(GND_net), .I1(n1_adj_4958[22]), 
            .CO(n45740));
    SB_CARRY add_4451_8 (.CI(n46448), .I0(n12098[5]), .I1(n518_adj_4743), 
            .CO(n46449));
    SB_CARRY add_4652_7 (.CI(n46581), .I0(n15793[4]), .I1(n460_adj_4748), 
            .CO(n46582));
    SB_LUT4 add_4782_4_lut (.I0(GND_net), .I1(n17498[1]), .I2(n256_adj_4752), 
            .I3(n46507), .O(n17257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_7_lut (.I0(GND_net), .I1(n12098[4]), .I2(n445_adj_4753), 
            .I3(n46447), .O(n11174[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4568_4 (.CI(n46381), .I0(n14382[1]), .I1(n235_adj_4749), 
            .CO(n46382));
    SB_LUT4 add_4723_11_lut (.I0(GND_net), .I1(n16802[8]), .I2(n761_adj_4754), 
            .I3(n46297), .O(n16438[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[21]), 
            .I3(n45738), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_11_lut (.I0(GND_net), .I1(n13337[8]), .I2(n740_adj_4757), 
            .I3(n46666), .O(n12538[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_23 (.CI(n45738), .I0(GND_net), .I1(n1_adj_4958[21]), 
            .CO(n45739));
    SB_LUT4 add_4652_6_lut (.I0(GND_net), .I1(n15793[3]), .I2(n387_adj_4758), 
            .I3(n46580), .O(n15282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_11 (.CI(n46297), .I0(n16802[8]), .I1(n761_adj_4754), 
            .CO(n46298));
    SB_LUT4 add_4568_3_lut (.I0(GND_net), .I1(n14382[0]), .I2(n162_adj_4759), 
            .I3(n46380), .O(n13698[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4723_10_lut (.I0(GND_net), .I1(n16802[7]), .I2(n688_adj_4760), 
            .I3(n46296), .O(n16438[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_10 (.CI(n46296), .I0(n16802[7]), .I1(n688_adj_4760), 
            .CO(n46297));
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[20]), 
            .I3(n45737), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_4 (.CI(n46507), .I0(n17498[1]), .I1(n256_adj_4752), 
            .CO(n46508));
    SB_CARRY add_4451_7 (.CI(n46447), .I0(n12098[4]), .I1(n445_adj_4753), 
            .CO(n46448));
    SB_CARRY add_4568_3 (.CI(n46380), .I0(n14382[0]), .I1(n162_adj_4759), 
            .CO(n46381));
    SB_LUT4 add_4723_9_lut (.I0(GND_net), .I1(n16802[6]), .I2(n615_adj_4762), 
            .I3(n46295), .O(n16438[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n46198), .O(n51[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(n9_adj_1), 
            .I3(n45593), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_24 (.CI(n45593), .I0(setpoint[22]), .I1(n9_adj_1), 
            .CO(n45594));
    SB_CARRY unary_minus_26_add_3_22 (.CI(n45737), .I0(GND_net), .I1(n1_adj_4958[20]), 
            .CO(n45738));
    SB_CARRY add_4512_11 (.CI(n46666), .I0(n13337[8]), .I1(n740_adj_4757), 
            .CO(n46667));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[19]), 
            .I3(n45736), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n45736), .I0(GND_net), .I1(n1_adj_4958[19]), 
            .CO(n45737));
    SB_CARRY add_4652_6 (.CI(n46580), .I0(n15793[3]), .I1(n387_adj_4758), 
            .CO(n46581));
    SB_LUT4 add_4782_3_lut (.I0(GND_net), .I1(n17498[0]), .I2(n183_adj_4765), 
            .I3(n46506), .O(n17257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[18]), 
            .I3(n45735), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_6_lut (.I0(GND_net), .I1(n12098[3]), .I2(n372_adj_4768), 
            .I3(n46446), .O(n11174[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_20 (.CI(n45735), .I0(GND_net), .I1(n1_adj_4958[18]), 
            .CO(n45736));
    SB_CARRY add_4451_6 (.CI(n46446), .I0(n12098[3]), .I1(n372_adj_4768), 
            .CO(n46447));
    SB_LUT4 counter_1935_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n46197), .O(n51[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_5_lut (.I0(GND_net), .I1(n15793[2]), .I2(n314_adj_4769), 
            .I3(n46579), .O(n15282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_3 (.CI(n46506), .I0(n17498[0]), .I1(n183_adj_4765), 
            .CO(n46507));
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[17]), 
            .I3(n45734), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4451_5_lut (.I0(GND_net), .I1(n12098[2]), .I2(n299_adj_4771), 
            .I3(n46445), .O(n11174[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_5 (.CI(n46445), .I0(n12098[2]), .I1(n299_adj_4771), 
            .CO(n46446));
    SB_LUT4 add_4512_10_lut (.I0(GND_net), .I1(n13337[7]), .I2(n667_adj_4772), 
            .I3(n46665), .O(n12538[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_19 (.CI(n45734), .I0(GND_net), .I1(n1_adj_4958[17]), 
            .CO(n45735));
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[16]), 
            .I3(n45733), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_10 (.CI(n46665), .I0(n13337[7]), .I1(n667_adj_4772), 
            .CO(n46666));
    SB_CARRY unary_minus_26_add_3_18 (.CI(n45733), .I0(GND_net), .I1(n1_adj_4958[16]), 
            .CO(n45734));
    SB_CARRY add_4652_5 (.CI(n46579), .I0(n15793[2]), .I1(n314_adj_4769), 
            .CO(n46580));
    SB_LUT4 add_4782_2_lut (.I0(GND_net), .I1(n41_adj_4774), .I2(n110_adj_4775), 
            .I3(GND_net), .O(n17257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4782_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_9 (.CI(n46295), .I0(n16802[6]), .I1(n615_adj_4762), 
            .CO(n46296));
    SB_LUT4 add_4451_4_lut (.I0(GND_net), .I1(n12098[1]), .I2(n226_adj_4776), 
            .I3(n46444), .O(n11174[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_4 (.CI(n46444), .I0(n12098[1]), .I1(n226_adj_4776), 
            .CO(n46445));
    SB_CARRY counter_1935_add_4_32 (.CI(n46197), .I0(GND_net), .I1(counter[30]), 
            .CO(n46198));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[15]), 
            .I3(n45732), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n45732), .I0(GND_net), .I1(n1_adj_4958[15]), 
            .CO(n45733));
    SB_LUT4 add_4652_4_lut (.I0(GND_net), .I1(n15793[1]), .I2(n241_adj_4779), 
            .I3(n46578), .O(n15282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4782_2 (.CI(GND_net), .I0(n41_adj_4774), .I1(n110_adj_4775), 
            .CO(n46506));
    SB_LUT4 add_4451_3_lut (.I0(GND_net), .I1(n12098[0]), .I2(n153_adj_4780), 
            .I3(n46443), .O(n11174[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n46196), .O(n51[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4451_3 (.CI(n46443), .I0(n12098[0]), .I1(n153_adj_4780), 
            .CO(n46444));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[14]), 
            .I3(n45731), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_16 (.CI(n45731), .I0(GND_net), .I1(n1_adj_4958[14]), 
            .CO(n45732));
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[13]), 
            .I3(n45730), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_31 (.CI(n46196), .I0(GND_net), .I1(counter[29]), 
            .CO(n46197));
    SB_LUT4 add_4723_8_lut (.I0(GND_net), .I1(n16802[5]), .I2(n542_adj_4783), 
            .I3(n46294), .O(n16438[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n46195), .O(n51[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_15 (.CI(n45730), .I0(GND_net), .I1(n1_adj_4958[13]), 
            .CO(n45731));
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n45592), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_23 (.CI(n45592), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n45593));
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[12]), 
            .I3(n45729), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_30 (.CI(n46195), .I0(GND_net), .I1(counter[28]), 
            .CO(n46196));
    SB_LUT4 add_4568_2_lut (.I0(GND_net), .I1(n20_adj_4786), .I2(n89_adj_4787), 
            .I3(GND_net), .O(n13698[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_8 (.CI(n46294), .I0(n16802[5]), .I1(n542_adj_4783), 
            .CO(n46295));
    SB_LUT4 counter_1935_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n46194), .O(n51[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n45729), .I0(GND_net), .I1(n1_adj_4958[12]), 
            .CO(n45730));
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[11]), 
            .I3(n45728), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_29 (.CI(n46194), .I0(GND_net), .I1(counter[27]), 
            .CO(n46195));
    SB_LUT4 add_4723_7_lut (.I0(GND_net), .I1(n16802[4]), .I2(n469_adj_4789), 
            .I3(n46293), .O(n16438[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n46193), .O(n51[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_9_lut (.I0(GND_net), .I1(n13337[6]), .I2(n594_adj_4790), 
            .I3(n46664), .O(n12538[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_4 (.CI(n46578), .I0(n15793[1]), .I1(n241_adj_4779), 
            .CO(n46579));
    SB_LUT4 add_4451_2_lut (.I0(GND_net), .I1(n11_adj_4791), .I2(n80_adj_4792), 
            .I3(GND_net), .O(n11174[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4451_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4793));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3691[23] ), 
            .I1(n10158[21]), .I2(GND_net), .I3(n46505), .O(n9651[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4451_2 (.CI(GND_net), .I0(n11_adj_4791), .I1(n80_adj_4792), 
            .CO(n46443));
    SB_CARRY add_4568_2 (.CI(GND_net), .I0(n20_adj_4786), .I1(n89_adj_4787), 
            .CO(n46380));
    SB_CARRY add_4723_7 (.CI(n46293), .I0(n16802[4]), .I1(n469_adj_4789), 
            .CO(n46294));
    SB_CARRY unary_minus_26_add_3_13 (.CI(n45728), .I0(GND_net), .I1(n1_adj_4958[11]), 
            .CO(n45729));
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[10]), 
            .I3(n45727), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_28 (.CI(n46193), .I0(GND_net), .I1(counter[26]), 
            .CO(n46194));
    SB_CARRY unary_minus_26_add_3_12 (.CI(n45727), .I0(GND_net), .I1(n1_adj_4958[10]), 
            .CO(n45728));
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[9]), 
            .I3(n45726), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n45591), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_9 (.CI(n46664), .I0(n13337[6]), .I1(n594_adj_4790), 
            .CO(n46665));
    SB_LUT4 add_4652_3_lut (.I0(GND_net), .I1(n15793[0]), .I2(n168_adj_4797), 
            .I3(n46577), .O(n15282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4652_3 (.CI(n46577), .I0(n15793[0]), .I1(n168_adj_4797), 
            .CO(n46578));
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n356[15]), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4798));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4799));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n45726), .I0(GND_net), .I1(n1_adj_4958[9]), 
            .CO(n45727));
    SB_LUT4 counter_1935_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n46192), .O(n51[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[8]), 
            .I3(n45725), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n45725), .I0(GND_net), .I1(n1_adj_4958[8]), 
            .CO(n45726));
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4801));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4723_6_lut (.I0(GND_net), .I1(n16802[3]), .I2(n396_adj_4802), 
            .I3(n46292), .O(n16438[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4803));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4804));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[7]), 
            .I3(n45724), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_22 (.CI(n45591), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n45592));
    SB_CARRY unary_minus_26_add_3_9 (.CI(n45724), .I0(GND_net), .I1(n1_adj_4958[7]), 
            .CO(n45725));
    SB_CARRY counter_1935_add_4_27 (.CI(n46192), .I0(GND_net), .I1(counter[25]), 
            .CO(n46193));
    SB_LUT4 add_4512_8_lut (.I0(GND_net), .I1(n13337[5]), .I2(n521_adj_4806), 
            .I3(n46663), .O(n12538[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[6]), 
            .I3(n45723), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_8 (.CI(n45723), .I0(GND_net), .I1(n1_adj_4958[6]), 
            .CO(n45724));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[5]), 
            .I3(n45722), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_8 (.CI(n46663), .I0(n13337[5]), .I1(n521_adj_4806), 
            .CO(n46664));
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n45590), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_7_lut (.I0(GND_net), .I1(n13337[4]), .I2(n448_adj_4810), 
            .I3(n46662), .O(n12538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4652_2_lut (.I0(GND_net), .I1(n26_adj_4811), .I2(n95_adj_4812), 
            .I3(GND_net), .O(n15282[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4652_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n46191), .O(n51[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n45722), .I0(GND_net), .I1(n1_adj_4958[5]), 
            .CO(n45723));
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[4]), 
            .I3(n45721), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_7 (.CI(n46662), .I0(n13337[4]), .I1(n448_adj_4810), 
            .CO(n46663));
    SB_LUT4 add_4512_6_lut (.I0(GND_net), .I1(n13337[3]), .I2(n375_adj_4814), 
            .I3(n46661), .O(n12538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_6 (.CI(n46661), .I0(n13337[3]), .I1(n375_adj_4814), 
            .CO(n46662));
    SB_CARRY add_4652_2 (.CI(GND_net), .I0(n26_adj_4811), .I1(n95_adj_4812), 
            .CO(n46577));
    SB_LUT4 add_4682_16_lut (.I0(GND_net), .I1(n16242[13]), .I2(n1120_adj_4815), 
            .I3(n46576), .O(n15793[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4816));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4817));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4820_10_lut (.I0(GND_net), .I1(n17858[7]), .I2(n700_adj_4818), 
            .I3(n46379), .O(n17697[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_6 (.CI(n45721), .I0(GND_net), .I1(n1_adj_4958[4]), 
            .CO(n45722));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[3]), 
            .I3(n45720), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4821));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n45720), .I0(GND_net), .I1(n1_adj_4958[3]), 
            .CO(n45721));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[2]), 
            .I3(n45719), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n45719), .I0(GND_net), .I1(n1_adj_4958[2]), 
            .CO(n45720));
    SB_LUT4 add_4820_9_lut (.I0(GND_net), .I1(n17858[6]), .I2(n627_adj_4823), 
            .I3(n46378), .O(n17697[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4723_6 (.CI(n46292), .I0(n16802[3]), .I1(n396_adj_4802), 
            .CO(n46293));
    SB_CARRY counter_1935_add_4_26 (.CI(n46191), .I0(GND_net), .I1(counter[24]), 
            .CO(n46192));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[1]), 
            .I3(n45718), .O(n436[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n46190), .O(n51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4512_5_lut (.I0(GND_net), .I1(n13337[2]), .I2(n302_adj_4825), 
            .I3(n46660), .O(n12538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4826));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4682_15_lut (.I0(GND_net), .I1(n16242[12]), .I2(n1047_adj_4827), 
            .I3(n46575), .O(n15793[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n10158[20]), .I2(GND_net), 
            .I3(n46504), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_5 (.CI(n46660), .I0(n13337[2]), .I1(n302_adj_4825), 
            .CO(n46661));
    SB_LUT4 add_4512_4_lut (.I0(GND_net), .I1(n13337[1]), .I2(n229_adj_4828), 
            .I3(n46659), .O(n12538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_15 (.CI(n46575), .I0(n16242[12]), .I1(n1047_adj_4827), 
            .CO(n46576));
    SB_CARRY add_4512_4 (.CI(n46659), .I0(n13337[1]), .I1(n229_adj_4828), 
            .CO(n46660));
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4829));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4512_3_lut (.I0(GND_net), .I1(n13337[0]), .I2(n156_adj_4830), 
            .I3(n46658), .O(n12538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_25 (.CI(n46190), .I0(GND_net), .I1(counter[23]), 
            .CO(n46191));
    SB_CARRY mult_17_add_1225_23 (.CI(n46504), .I0(n10158[20]), .I1(GND_net), 
            .CO(n46505));
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n10158[19]), .I2(GND_net), 
            .I3(n46503), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_21_lut (.I0(GND_net), .I1(n12938[18]), .I2(GND_net), 
            .I3(n46442), .O(n12098[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4682_14_lut (.I0(GND_net), .I1(n16242[11]), .I2(n974_adj_4831), 
            .I3(n46574), .O(n15793[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n46503), .I0(n10158[19]), .I1(GND_net), 
            .CO(n46504));
    SB_LUT4 add_4492_20_lut (.I0(GND_net), .I1(n12938[17]), .I2(GND_net), 
            .I3(n46441), .O(n12098[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n45718), .I0(GND_net), .I1(n1_adj_4958[1]), 
            .CO(n45719));
    SB_LUT4 add_4723_5_lut (.I0(GND_net), .I1(n16802[2]), .I2(n323_adj_4832), 
            .I3(n46291), .O(n16438[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n46189), .O(n51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4958[0]), 
            .I3(VCC_net), .O(n436[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4835));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4958[0]), 
            .CO(n45718));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_4956[23]), 
            .I3(n45717), .O(n47_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4723_5 (.CI(n46291), .I0(n16802[2]), .I1(n323_adj_4832), 
            .CO(n46292));
    SB_CARRY counter_1935_add_4_24 (.CI(n46189), .I0(GND_net), .I1(counter[22]), 
            .CO(n46190));
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4837));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4682_14 (.CI(n46574), .I0(n16242[11]), .I1(n974_adj_4831), 
            .CO(n46575));
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n10158[18]), .I2(GND_net), 
            .I3(n46502), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4682_13_lut (.I0(GND_net), .I1(n16242[10]), .I2(n901_adj_4838), 
            .I3(n46573), .O(n15793[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n46502), .I0(n10158[18]), .I1(GND_net), 
            .CO(n46503));
    SB_CARRY add_4682_13 (.CI(n46573), .I0(n16242[10]), .I1(n901_adj_4838), 
            .CO(n46574));
    SB_LUT4 add_4682_12_lut (.I0(GND_net), .I1(n16242[9]), .I2(n828_adj_4839), 
            .I3(n46572), .O(n15793[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_3 (.CI(n46658), .I0(n13337[0]), .I1(n156_adj_4830), 
            .CO(n46659));
    SB_CARRY add_4682_12 (.CI(n46572), .I0(n16242[9]), .I1(n828_adj_4839), 
            .CO(n46573));
    SB_LUT4 add_4512_2_lut (.I0(GND_net), .I1(n14_adj_4840), .I2(n83_adj_4841), 
            .I3(GND_net), .O(n12538[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4512_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4682_11_lut (.I0(GND_net), .I1(n16242[8]), .I2(n755_adj_4842), 
            .I3(n46571), .O(n15793[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_11 (.CI(n46571), .I0(n16242[8]), .I1(n755_adj_4842), 
            .CO(n46572));
    SB_LUT4 add_4682_10_lut (.I0(GND_net), .I1(n16242[7]), .I2(n682_adj_4843), 
            .I3(n46570), .O(n15793[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n10158[17]), .I2(GND_net), 
            .I3(n46501), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4512_2 (.CI(GND_net), .I0(n14_adj_4840), .I1(n83_adj_4841), 
            .CO(n46658));
    SB_LUT4 add_4550_20_lut (.I0(GND_net), .I1(n14058[17]), .I2(GND_net), 
            .I3(n46657), .O(n13337[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n46501), .I0(n10158[17]), .I1(GND_net), 
            .CO(n46502));
    SB_CARRY add_4682_10 (.CI(n46570), .I0(n16242[7]), .I1(n682_adj_4843), 
            .CO(n46571));
    SB_LUT4 add_4550_19_lut (.I0(GND_net), .I1(n14058[16]), .I2(GND_net), 
            .I3(n46656), .O(n13337[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n10158[16]), .I2(GND_net), 
            .I3(n46500), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_20 (.CI(n46441), .I0(n12938[17]), .I1(GND_net), 
            .CO(n46442));
    SB_CARRY sub_8_add_2_21 (.CI(n45590), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n45591));
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4844));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4723_4_lut (.I0(GND_net), .I1(n16802[1]), .I2(n250_adj_4845), 
            .I3(n46290), .O(n16438[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n46188), .O(n51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[22]), 
            .I3(n45716), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1935_add_4_23 (.CI(n46188), .I0(GND_net), .I1(counter[21]), 
            .CO(n46189));
    SB_CARRY add_4550_19 (.CI(n46656), .I0(n14058[16]), .I1(GND_net), 
            .CO(n46657));
    SB_LUT4 add_4550_18_lut (.I0(GND_net), .I1(n14058[15]), .I2(GND_net), 
            .I3(n46655), .O(n13337[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4847));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n45716), .I0(GND_net), .I1(n1_adj_4956[22]), 
            .CO(n45717));
    SB_CARRY add_4820_9 (.CI(n46378), .I0(n17858[6]), .I1(n627_adj_4823), 
            .CO(n46379));
    SB_LUT4 add_4492_19_lut (.I0(GND_net), .I1(n12938[16]), .I2(GND_net), 
            .I3(n46440), .O(n12098[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_19 (.CI(n46440), .I0(n12938[16]), .I1(GND_net), 
            .CO(n46441));
    SB_LUT4 add_4682_9_lut (.I0(GND_net), .I1(n16242[6]), .I2(n609_adj_4848), 
            .I3(n46569), .O(n15793[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_18_lut (.I0(GND_net), .I1(n12938[15]), .I2(GND_net), 
            .I3(n46439), .O(n12098[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n46500), .I0(n10158[16]), .I1(GND_net), 
            .CO(n46501));
    SB_CARRY add_4682_9 (.CI(n46569), .I0(n16242[6]), .I1(n609_adj_4848), 
            .CO(n46570));
    SB_CARRY add_4550_18 (.CI(n46655), .I0(n14058[15]), .I1(GND_net), 
            .CO(n46656));
    SB_LUT4 add_4820_8_lut (.I0(GND_net), .I1(n17858[5]), .I2(n554_adj_4849), 
            .I3(n46377), .O(n17697[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4550_17_lut (.I0(GND_net), .I1(n14058[14]), .I2(GND_net), 
            .I3(n46654), .O(n13337[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n10158[15]), .I2(GND_net), 
            .I3(n46499), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4820_8 (.CI(n46377), .I0(n17858[5]), .I1(n554_adj_4849), 
            .CO(n46378));
    SB_CARRY add_4550_17 (.CI(n46654), .I0(n14058[14]), .I1(GND_net), 
            .CO(n46655));
    SB_CARRY add_4492_18 (.CI(n46439), .I0(n12938[15]), .I1(GND_net), 
            .CO(n46440));
    SB_CARRY mult_17_add_1225_18 (.CI(n46499), .I0(n10158[15]), .I1(GND_net), 
            .CO(n46500));
    SB_LUT4 add_4682_8_lut (.I0(GND_net), .I1(n16242[5]), .I2(n536_adj_4850), 
            .I3(n46568), .O(n15793[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4550_16_lut (.I0(GND_net), .I1(n14058[13]), .I2(n1108_adj_4851), 
            .I3(n46653), .O(n13337[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[21]), 
            .I3(n45715), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n45715), .I0(GND_net), .I1(n1_adj_4956[21]), 
            .CO(n45716));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[20]), 
            .I3(n45714), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31882_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n45445), 
            .I3(n18202[0]), .O(n4_adj_4475));   // verilog/motorControl.v(50[18:24])
    defparam i31882_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n45714), .I0(GND_net), .I1(n1_adj_4956[20]), 
            .CO(n45715));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[19]), 
            .I3(n45713), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n46187), .O(n51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n45713), .I0(GND_net), .I1(n1_adj_4956[19]), 
            .CO(n45714));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[18]), 
            .I3(n45712), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4492_17_lut (.I0(GND_net), .I1(n12938[14]), .I2(GND_net), 
            .I3(n46438), .O(n12098[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_16 (.CI(n46653), .I0(n14058[13]), .I1(n1108_adj_4851), 
            .CO(n46654));
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n10158[14]), .I2(GND_net), 
            .I3(n46498), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_17 (.CI(n46438), .I0(n12938[14]), .I1(GND_net), 
            .CO(n46439));
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4856));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_17_add_1225_17 (.CI(n46498), .I0(n10158[14]), .I1(GND_net), 
            .CO(n46499));
    SB_CARRY add_4682_8 (.CI(n46568), .I0(n16242[5]), .I1(n536_adj_4850), 
            .CO(n46569));
    SB_LUT4 add_4550_15_lut (.I0(GND_net), .I1(n14058[12]), .I2(n1035_adj_4857), 
            .I3(n46652), .O(n13337[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4858));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4682_7_lut (.I0(GND_net), .I1(n16242[4]), .I2(n463_adj_4859), 
            .I3(n46567), .O(n15793[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_15 (.CI(n46652), .I0(n14058[12]), .I1(n1035_adj_4857), 
            .CO(n46653));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n45712), .I0(GND_net), .I1(n1_adj_4956[18]), 
            .CO(n45713));
    SB_LUT4 add_4492_16_lut (.I0(GND_net), .I1(n12938[13]), .I2(n1105_adj_4860), 
            .I3(n46437), .O(n12098[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[17]), 
            .I3(n45711), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n45711), .I0(GND_net), .I1(n1_adj_4956[17]), 
            .CO(n45712));
    SB_LUT4 add_4550_14_lut (.I0(GND_net), .I1(n14058[11]), .I2(n962_adj_4862), 
            .I3(n46651), .O(n13337[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4820_7_lut (.I0(GND_net), .I1(n17858[4]), .I2(n481_adj_4863), 
            .I3(n46376), .O(n17697[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_14 (.CI(n46651), .I0(n14058[11]), .I1(n962_adj_4862), 
            .CO(n46652));
    SB_CARRY add_4820_7 (.CI(n46376), .I0(n17858[4]), .I1(n481_adj_4863), 
            .CO(n46377));
    SB_CARRY add_4682_7 (.CI(n46567), .I0(n16242[4]), .I1(n463_adj_4859), 
            .CO(n46568));
    SB_CARRY add_4723_4 (.CI(n46290), .I0(n16802[1]), .I1(n250_adj_4845), 
            .CO(n46291));
    SB_CARRY counter_1935_add_4_22 (.CI(n46187), .I0(GND_net), .I1(counter[20]), 
            .CO(n46188));
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4864));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n356[17]), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4865));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[16]), 
            .I3(n45710), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n45710), .I0(GND_net), .I1(n1_adj_4956[16]), 
            .CO(n45711));
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4867));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), .I3(GND_net), 
            .O(n9_adj_4868));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4869));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4870));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4550_13_lut (.I0(GND_net), .I1(n14058[10]), .I2(n889_adj_4871), 
            .I3(n46650), .O(n13337[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4872));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4550_13 (.CI(n46650), .I0(n14058[10]), .I1(n889_adj_4871), 
            .CO(n46651));
    SB_LUT4 add_4682_6_lut (.I0(GND_net), .I1(n16242[3]), .I2(n390_adj_4873), 
            .I3(n46566), .O(n15793[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45265_4_lut (.I0(n21_adj_4683), .I1(n19_adj_4867), .I2(n17_adj_4858), 
            .I3(n9_adj_4793), .O(n60165));
    defparam i45265_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4550_12_lut (.I0(GND_net), .I1(n14058[9]), .I2(n816_adj_4874), 
            .I3(n46649), .O(n13337[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n10158[13]), .I2(n1096_adj_4875), 
            .I3(n46497), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4820_6_lut (.I0(GND_net), .I1(n17858[3]), .I2(n408_adj_4876), 
            .I3(n46375), .O(n17697[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4820_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45248_4_lut (.I0(n27_adj_4648), .I1(n15_adj_4847), .I2(n13_adj_4816), 
            .I3(n11_adj_4801), .O(n60148));
    defparam i45248_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4550_12 (.CI(n46649), .I0(n14058[9]), .I1(n816_adj_4874), 
            .CO(n46650));
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4877));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4682_6 (.CI(n46566), .I0(n16242[3]), .I1(n390_adj_4873), 
            .CO(n46567));
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4682_5_lut (.I0(GND_net), .I1(n16242[2]), .I2(n317_adj_4878), 
            .I3(n46565), .O(n15793[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4682_5 (.CI(n46565), .I0(n16242[2]), .I1(n317_adj_4878), 
            .CO(n46566));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4956[15]), 
            .I3(n45709), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4550_11_lut (.I0(GND_net), .I1(n14058[8]), .I2(n743_adj_4879), 
            .I3(n46648), .O(n13337[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n46497), .I0(n10158[13]), .I1(n1096_adj_4875), 
            .CO(n46498));
    SB_CARRY add_4550_11 (.CI(n46648), .I0(n14058[8]), .I1(n743_adj_4879), 
            .CO(n46649));
    SB_LUT4 add_4682_4_lut (.I0(GND_net), .I1(n16242[1]), .I2(n244_adj_4880), 
            .I3(n46564), .O(n15793[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n10158[12]), .I2(n1023_adj_4881), 
            .I3(n46496), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_16 (.CI(n46437), .I0(n12938[13]), .I1(n1105_adj_4860), 
            .CO(n46438));
    SB_LUT4 add_4492_15_lut (.I0(GND_net), .I1(n12938[12]), .I2(n1032_adj_4882), 
            .I3(n46436), .O(n12098[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4492_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4492_15 (.CI(n46436), .I0(n12938[12]), .I1(n1032_adj_4882), 
            .CO(n46437));
    SB_LUT4 counter_1935_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n46186), .O(n51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_4817), 
            .I3(GND_net), .O(n12_adj_4883));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY counter_1935_add_4_21 (.CI(n46186), .I0(GND_net), .I1(counter[19]), 
            .CO(n46187));
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4682_4 (.CI(n46564), .I0(n16242[1]), .I1(n244_adj_4880), 
            .CO(n46565));
    SB_CARRY mult_17_add_1225_15 (.CI(n46496), .I0(n10158[12]), .I1(n1023_adj_4881), 
            .CO(n46497));
    SB_LUT4 add_4682_3_lut (.I0(GND_net), .I1(n16242[0]), .I2(n171_adj_4884), 
            .I3(n46563), .O(n15793[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4682_3 (.CI(n46563), .I0(n16242[0]), .I1(n171_adj_4884), 
            .CO(n46564));
    SB_CARRY add_4820_6 (.CI(n46375), .I0(n17858[3]), .I1(n408_adj_4876), 
            .CO(n46376));
    SB_LUT4 add_4550_10_lut (.I0(GND_net), .I1(n14058[7]), .I2(n670_adj_4885), 
            .I3(n46647), .O(n13337[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4682_2_lut (.I0(GND_net), .I1(n29_adj_4886), .I2(n98_adj_4887), 
            .I3(GND_net), .O(n15793[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4682_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4682_2 (.CI(GND_net), .I0(n29_adj_4886), .I1(n98_adj_4887), 
            .CO(n46563));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n10158[11]), .I2(n950_adj_4888), 
            .I3(n46495), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4843_8_lut (.I0(GND_net), .I1(n18034[5]), .I2(n560_adj_4889), 
            .I3(n46562), .O(n17922[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_10 (.CI(n46647), .I0(n14058[7]), .I1(n670_adj_4885), 
            .CO(n46648));
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4420));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_4816), 
            .I3(GND_net), .O(n10_adj_4890));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4891));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46576_3_lut (.I0(n4_adj_4892), .I1(n436[2]), .I2(n356[2]), 
            .I3(GND_net), .O(n61476));   // verilog/motorControl.v(54[23:39])
    defparam i46576_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46577_3_lut (.I0(n61476), .I1(n436[3]), .I2(n356[3]), .I3(GND_net), 
            .O(n8_adj_4893));   // verilog/motorControl.v(54[23:39])
    defparam i46577_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4894));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_17_add_1225_14 (.CI(n46495), .I0(n10158[11]), .I1(n950_adj_4888), 
            .CO(n46496));
    SB_LUT4 add_4550_9_lut (.I0(GND_net), .I1(n14058[6]), .I2(n597_adj_4895), 
            .I3(n46646), .O(n13337[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4723_3_lut (.I0(GND_net), .I1(n16802[0]), .I2(n177), .I3(n46289), 
            .O(n16438[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4723_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1935_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n46185), .O(n51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1935_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4843_7_lut (.I0(GND_net), .I1(n18034[4]), .I2(n487), .I3(n46561), 
            .O(n17922[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4843_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4550_9 (.CI(n46646), .I0(n14058[6]), .I1(n597_adj_4895), 
            .CO(n46647));
    SB_LUT4 add_4550_8_lut (.I0(GND_net), .I1(n14058[5]), .I2(n524), .I3(n46645), 
            .O(n13337[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4550_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n10158[10]), .I2(n877), 
            .I3(n46494), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_4883), .I1(n182[17]), .I2(n35_adj_4829), 
            .I3(GND_net), .O(n30_adj_4896));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44757_4_lut (.I0(n33_adj_4894), .I1(n21_adj_4869), .I2(n19_adj_4864), 
            .I3(n17_adj_4891), .O(n59657));
    defparam i44757_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46129_4_lut (.I0(n13_adj_4816), .I1(n11_adj_4801), .I2(n9_adj_4793), 
            .I3(n60212), .O(n61029));
    defparam i46129_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46123_4_lut (.I0(n19_adj_4867), .I1(n17_adj_4858), .I2(n15_adj_4847), 
            .I3(n61029), .O(n61023));
    defparam i46123_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i45779_4_lut (.I0(n15_adj_4826), .I1(n13_adj_4821), .I2(n375), 
            .I3(n436[5]), .O(n60679));
    defparam i45779_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i31869_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n18153[0]));   // verilog/motorControl.v(50[18:24])
    defparam i31869_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i47033_4_lut (.I0(n25_adj_4716), .I1(n23_adj_4715), .I2(n21_adj_4683), 
            .I3(n61023), .O(n61933));
    defparam i47033_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31793_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n18233[0]));   // verilog/motorControl.v(50[18:24])
    defparam i31793_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i46317_4_lut (.I0(n21_adj_4869), .I1(n19_adj_4864), .I2(n17_adj_4891), 
            .I3(n60679), .O(n61217));
    defparam i46317_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46479_4_lut (.I0(n31_adj_4668), .I1(n29_adj_4653), .I2(n27_adj_4648), 
            .I3(n61933), .O(n61379));
    defparam i46479_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31795_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n45363));   // verilog/motorControl.v(50[18:24])
    defparam i31795_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i47106_4_lut (.I0(n37_adj_4835), .I1(n35_adj_4829), .I2(n33_adj_4817), 
            .I3(n61379), .O(n62006));
    defparam i47106_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_4612), 
            .I3(GND_net), .O(n16_adj_4897));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46683_3_lut (.I0(n6), .I1(n182[10]), .I2(n21_adj_4683), .I3(GND_net), 
            .O(n61583));   // verilog/motorControl.v(47[21:44])
    defparam i46683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_2_lut_4_lut (.I0(control_update), .I1(n61965), .I2(PWMLimit[23]), 
            .I3(n356[23]), .O(n9611));
    defparam i4323_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 i46684_3_lut (.I0(n61583), .I1(n182[11]), .I2(n23_adj_4715), 
            .I3(GND_net), .O(n61584));   // verilog/motorControl.v(47[21:44])
    defparam i46684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4895));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_4858), 
            .I3(GND_net), .O(n8_adj_4899));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4888));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4887));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4886));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4885));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4884));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4882));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4881));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4880));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4879));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4878));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4876));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4875));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46293_4_lut (.I0(n27_adj_4803), .I1(n25_adj_4804), .I2(n23_adj_4837), 
            .I3(n61217), .O(n61193));
    defparam i46293_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4874));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4873));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4871));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[16]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4863));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4862));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31871_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n45445));   // verilog/motorControl.v(50[18:24])
    defparam i31871_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut_4_lut_adj_954 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n18233[0]), 
            .I3(n45395), .O(n18202[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_954.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[17]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4860));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4859));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4857));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[18]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[19]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[20]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_4897), .I1(n182[22]), .I2(n45_adj_4611), 
            .I3(GND_net), .O(n24_adj_4900));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[21]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4851));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4850));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4849));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4848));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[22]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4845));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4843));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4842));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4841));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4840));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44759_4_lut (.I0(n33_adj_4894), .I1(n31_adj_4798), .I2(n29_adj_4799), 
            .I3(n61193), .O(n59659));
    defparam i44759_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4839));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4838));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[23]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[0]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4832));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4831));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4830));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31836_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n45395), 
            .I3(n18233[0]), .O(n4_adj_4901));   // verilog/motorControl.v(50[18:24])
    defparam i31836_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4827));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4825));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[1]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4823));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[2]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[3]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4818));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4815));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4814));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[4]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4812));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20485_3_lut (.I0(n8_adj_4893), .I1(n356[4]), .I2(n436[4]), 
            .I3(GND_net), .O(n10_adj_4902));
    defparam i20485_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4811));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4810));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45199_4_lut (.I0(n43_adj_4612), .I1(n25_adj_4716), .I2(n23_adj_4715), 
            .I3(n60165), .O(n60099));
    defparam i45199_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46797_3_lut (.I0(n10_adj_4902), .I1(n436[16]), .I2(n33_adj_4894), 
            .I3(GND_net), .O(n61697));   // verilog/motorControl.v(54[23:39])
    defparam i46797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46267_4_lut (.I0(n24_adj_4900), .I1(n8_adj_4899), .I2(n45_adj_4611), 
            .I3(n60090), .O(n61167));   // verilog/motorControl.v(47[21:44])
    defparam i46267_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[5]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[6]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4806));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[7]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4802));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[8]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45597_3_lut (.I0(n61584), .I1(n182[12]), .I2(n25_adj_4716), 
            .I3(GND_net), .O(n60497));   // verilog/motorControl.v(47[21:44])
    defparam i45597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4797));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[9]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[10]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4792));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4791));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4790));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4789));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[11]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4787));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4786));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[12]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4783));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[13]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[14]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i18_3_lut (.I0(n436[10]), .I1(n436[19]), .I2(n39_adj_4872), 
            .I3(GND_net), .O(n18_adj_4903));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4780));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4779));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[15]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4776));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4775));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4774));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[16]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4772));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4771));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[17]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4769));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4768));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[18]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4765));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[19]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4762));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[20]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4760));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4759));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4757));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[21]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_4904));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4754));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4753));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4752));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[22]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46681_3_lut (.I0(n4_adj_4904), .I1(n182[13]), .I2(n27_adj_4648), 
            .I3(GND_net), .O(n61581));   // verilog/motorControl.v(47[21:44])
    defparam i46681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46682_3_lut (.I0(n61581), .I1(n182[14]), .I2(n29_adj_4653), 
            .I3(GND_net), .O(n61582));   // verilog/motorControl.v(47[21:44])
    defparam i46682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4750));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4748));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4958[23]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4746));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4745));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4744));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4742));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4741));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4740));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4739));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4738));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45240_4_lut (.I0(n33_adj_4817), .I1(n31_adj_4668), .I2(n29_adj_4653), 
            .I3(n60148), .O(n60140));
    defparam i45240_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46945_4_lut (.I0(n30_adj_4896), .I1(n10_adj_4890), .I2(n35_adj_4829), 
            .I3(n60132), .O(n61845));   // verilog/motorControl.v(47[21:44])
    defparam i46945_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4737));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4736));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4735));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4734));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4733));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4732));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4730));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4729));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4728));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4727));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4726));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4725));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4724));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4723));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4722));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4721));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4720));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4719));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4718));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45599_3_lut (.I0(n61582), .I1(n182[15]), .I2(n31_adj_4668), 
            .I3(GND_net), .O(n60499));   // verilog/motorControl.v(47[21:44])
    defparam i45599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4717));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4714));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47206_4_lut (.I0(n60499), .I1(n61845), .I2(n35_adj_4829), 
            .I3(n60140), .O(n62106));   // verilog/motorControl.v(47[21:44])
    defparam i47206_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4713));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47207_3_lut (.I0(n62106), .I1(n182[18]), .I2(n37_adj_4835), 
            .I3(GND_net), .O(n62107));   // verilog/motorControl.v(47[21:44])
    defparam i47207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4712));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4711));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4710));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4709));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4708));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[9]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4707));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4706));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4705));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[8]), .I1(n436[9]), .I2(n19_adj_4864), 
            .I3(GND_net), .O(n16_adj_4905));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4704));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4703));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4702));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47165_3_lut (.I0(n62107), .I1(n182[19]), .I2(n39_adj_4596), 
            .I3(GND_net), .O(n62065));   // verilog/motorControl.v(47[21:44])
    defparam i47165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4701));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45205_4_lut (.I0(n43_adj_4612), .I1(n41_adj_4600), .I2(n39_adj_4596), 
            .I3(n62006), .O(n60105));
    defparam i45205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4699));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4698));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4697));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4696));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4695));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4694));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4693));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4692));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46871_4_lut (.I0(n60497), .I1(n61167), .I2(n45_adj_4611), 
            .I3(n60099), .O(n61771));   // verilog/motorControl.v(47[21:44])
    defparam i46871_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4691));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4690));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4689));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4688));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4687));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4686));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4685));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4684));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4682));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4681));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4680));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4679));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4678));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i36_3_lut (.I0(n18_adj_4903), .I1(n436[20]), .I2(n41_adj_4856), 
            .I3(GND_net), .O(n36_adj_4906));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4677));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4676));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46798_3_lut (.I0(n61697), .I1(n436[17]), .I2(n35_adj_4865), 
            .I3(GND_net), .O(n61698));   // verilog/motorControl.v(54[23:39])
    defparam i46798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4675));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45605_3_lut (.I0(n62065), .I1(n182[20]), .I2(n41_adj_4600), 
            .I3(GND_net), .O(n60505));   // verilog/motorControl.v(47[21:44])
    defparam i45605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4674));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4673));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4672));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47059_4_lut (.I0(n60505), .I1(n61771), .I2(n45_adj_4611), 
            .I3(n60105), .O(n61959));   // verilog/motorControl.v(47[21:44])
    defparam i47059_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47060_3_lut (.I0(n61959), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(47[21:44])
    defparam i47060_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4671));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4670));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4669));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4667));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4666));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4665));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4664));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4663));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4662));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4661));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4660));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44704_4_lut (.I0(n39_adj_4872), .I1(n37_adj_4844), .I2(n35_adj_4865), 
            .I3(n59657), .O(n59604));
    defparam i44704_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4659));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4657));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4656));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4655));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4654));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[16] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4652));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4651));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4650));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4649));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11512_3_lut (.I0(n356[1]), .I1(n436[1]), .I2(n9613), .I3(GND_net), 
            .O(n25210));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24519_4_lut (.I0(PWMLimit[1]), .I1(n55139), .I2(n25210), 
            .I3(n9611), .O(n49[1]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24519_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4647));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4645));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4644));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4448));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4642));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4641));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11507_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n9613), .I3(GND_net), 
            .O(n25205));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47078_4_lut (.I0(n36_adj_4906), .I1(n16_adj_4905), .I2(n41_adj_4856), 
            .I3(n59592), .O(n61978));   // verilog/motorControl.v(54[23:39])
    defparam i47078_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4639));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4638));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4637));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46579_3_lut (.I0(n61698), .I1(n436[18]), .I2(n37_adj_4844), 
            .I3(GND_net), .O(n61479));   // verilog/motorControl.v(54[23:39])
    defparam i46579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4635));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4634));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4633));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4632));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24517_4_lut (.I0(PWMLimit[2]), .I1(n55139), .I2(n25205), 
            .I3(n9611), .O(n49[2]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24517_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n18178[2]), .I1(n6_adj_4907), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[18] ), .O(n18118[3]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h9666;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4630));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4629));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4628));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11502_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n9613), .I3(GND_net), 
            .O(n25200));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24516_4_lut (.I0(PWMLimit[3]), .I1(n55139), .I2(n25200), 
            .I3(n9611), .O(n49[3]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24516_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_956 (.I0(n18242[0]), .I1(n45231), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[20] ), .O(n18218[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h9666;
    SB_LUT4 i1_4_lut_adj_957 (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3691[23] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[22] ), .O(n56198));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_957.LUT_INIT = 16'h9c50;
    SB_LUT4 LessThan_25_i14_3_lut (.I0(n436[7]), .I1(n436[11]), .I2(n23_adj_4837), 
            .I3(GND_net), .O(n14_adj_4908));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_958 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[19] ), .O(n56202));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_959 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3691[20] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[21] ), .O(n56200));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_960 (.I0(n56200), .I1(n45429), .I2(n56202), .I3(n56198), 
            .O(n56208));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i20474_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n9613), .I3(GND_net), 
            .O(n34138));
    defparam i20474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31684_4_lut (.I0(n18242[0]), .I1(\Ki[2] ), .I2(n45231), .I3(\PID_CONTROLLER.integral_23__N_3691[20] ), 
            .O(n4_adj_4909));   // verilog/motorControl.v(50[27:38])
    defparam i31684_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i31776_4_lut (.I0(n18178[2]), .I1(\Ki[4] ), .I2(n6_adj_4907), 
            .I3(\PID_CONTROLLER.integral_23__N_3691[18] ), .O(n8_adj_4910));   // verilog/motorControl.v(50[27:38])
    defparam i31776_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_4821), 
            .I3(GND_net), .O(n12_adj_4911));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n6_adj_4912), .I1(n8_adj_4910), .I2(n4_adj_4909), 
            .I3(n56208), .O(n55037));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_962 (.I0(n55139), .I1(PWMLimit[4]), .I2(n34138), 
            .I3(n9611), .O(n49[4]));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'h5044;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4625));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4624));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4623));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4622));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4621));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4620));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11492_3_lut (.I0(n375), .I1(n436[5]), .I2(n9613), .I3(GND_net), 
            .O(n25190));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4619));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4618));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4617));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4616));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4615));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4614));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4613));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4610));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4609));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4608));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4607));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4606));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4605));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4604));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4603));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4602));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4601));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4599));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4598));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n55139), .I1(PWMLimit[5]), .I2(n25190), 
            .I3(n9611), .O(n49[5]));
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h5044;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4597));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4595));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4594));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4593));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4592));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4591));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i22_3_lut (.I0(n14_adj_4908), .I1(n436[12]), .I2(n25_adj_4804), 
            .I3(GND_net), .O(n22_adj_4913));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4590));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4589));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4588));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[10]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11487_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n9613), .I3(GND_net), 
            .O(n25185));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4587));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4586));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24515_4_lut (.I0(PWMLimit[6]), .I1(n55139), .I2(n25185), 
            .I3(n9611), .O(n49[6]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24515_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4583));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4582));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4581));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46893_4_lut (.I0(n22_adj_4913), .I1(n12_adj_4911), .I2(n25_adj_4804), 
            .I3(n59720), .O(n61793));   // verilog/motorControl.v(54[23:39])
    defparam i46893_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11482_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n9613), .I3(GND_net), 
            .O(n25180));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24514_4_lut (.I0(PWMLimit[7]), .I1(n55139), .I2(n25180), 
            .I3(n9611), .O(n49[7]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24514_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4579));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4576));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4575));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4574));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11477_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n9613), .I3(GND_net), 
            .O(n25175));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46894_3_lut (.I0(n61793), .I1(n436[13]), .I2(n27_adj_4803), 
            .I3(GND_net), .O(n61794));   // verilog/motorControl.v(54[23:39])
    defparam i46894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46593_3_lut (.I0(n61794), .I1(n436[14]), .I2(n29_adj_4799), 
            .I3(GND_net), .O(n61493));   // verilog/motorControl.v(54[23:39])
    defparam i46593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46558_4_lut (.I0(n39_adj_4872), .I1(n37_adj_4844), .I2(n35_adj_4865), 
            .I3(n59659), .O(n61458));
    defparam i46558_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24513_4_lut (.I0(PWMLimit[8]), .I1(n55139), .I2(n25175), 
            .I3(n9611), .O(n49[8]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24513_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i47210_4_lut (.I0(n61479), .I1(n61978), .I2(n41_adj_4856), 
            .I3(n59604), .O(n62110));   // verilog/motorControl.v(54[23:39])
    defparam i47210_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4568));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11472_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n9613), .I3(GND_net), 
            .O(n25170));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24512_4_lut (.I0(PWMLimit[9]), .I1(n55139), .I2(n25170), 
            .I3(n9611), .O(n49[9]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24512_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4567));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45639_3_lut (.I0(n61493), .I1(n436[15]), .I2(n31_adj_4798), 
            .I3(GND_net), .O(n60539));   // verilog/motorControl.v(54[23:39])
    defparam i45639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4566));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4565));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11467_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n9613), .I3(GND_net), 
            .O(n25165));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44894_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(PWMLimit[9]), 
            .I3(n356[9]), .O(n59794));
    defparam i44894_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4564));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24511_4_lut (.I0(PWMLimit[10]), .I1(n55139), .I2(n25165), 
            .I3(n9611), .O(n49[10]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24511_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i47250_4_lut (.I0(n60539), .I1(n62110), .I2(n41_adj_4856), 
            .I3(n61458), .O(n62150));   // verilog/motorControl.v(54[23:39])
    defparam i47250_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11462_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n9613), .I3(GND_net), 
            .O(n25160));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47251_3_lut (.I0(n62150), .I1(n436[21]), .I2(n356[21]), .I3(GND_net), 
            .O(n62151));   // verilog/motorControl.v(54[23:39])
    defparam i47251_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24510_4_lut (.I0(PWMLimit[11]), .I1(n55139), .I2(n25160), 
            .I3(n9611), .O(n49[11]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24510_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44934_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(PWMLimit[7]), 
            .I3(n356[7]), .O(n59834));
    defparam i44934_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i11457_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n9613), .I3(GND_net), 
            .O(n25155));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24509_4_lut (.I0(PWMLimit[12]), .I1(n55139), .I2(n25155), 
            .I3(n9611), .O(n49[12]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24509_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11452_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n9613), .I3(GND_net), 
            .O(n25150));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24508_4_lut (.I0(PWMLimit[13]), .I1(n55139), .I2(n25150), 
            .I3(n9611), .O(n49[13]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24508_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i47247_3_lut (.I0(n62151), .I1(n436[22]), .I2(n356[22]), .I3(GND_net), 
            .O(n62147));   // verilog/motorControl.v(54[23:39])
    defparam i47247_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11447_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n9613), .I3(GND_net), 
            .O(n25145));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24507_4_lut (.I0(PWMLimit[14]), .I1(n55139), .I2(n25145), 
            .I3(n9611), .O(n49[14]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24507_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11442_3_lut (.I0(n356[15]), .I1(n436[15]), .I2(n9613), .I3(GND_net), 
            .O(n25140));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24506_4_lut (.I0(PWMLimit[15]), .I1(n55139), .I2(n25140), 
            .I3(n9611), .O(n49[15]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24506_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_25_i48_3_lut (.I0(n62147), .I1(n356[23]), .I2(n436[23]), 
            .I3(GND_net), .O(n435));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11437_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n9613), .I3(GND_net), 
            .O(n25135));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24501_4_lut (.I0(PWMLimit[16]), .I1(n55139), .I2(n25135), 
            .I3(n9611), .O(n49[16]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24501_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11432_3_lut (.I0(n356[17]), .I1(n436[17]), .I2(n9613), .I3(GND_net), 
            .O(n25130));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24499_4_lut (.I0(PWMLimit[17]), .I1(n55139), .I2(n25130), 
            .I3(n9611), .O(n49[17]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24499_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11427_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n9613), .I3(GND_net), 
            .O(n25125));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4548));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24498_4_lut (.I0(PWMLimit[18]), .I1(n55139), .I2(n25125), 
            .I3(n9611), .O(n49[18]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24498_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i4325_3_lut (.I0(control_update), .I1(n409), .I2(n435), .I3(GND_net), 
            .O(n9613));   // verilog/motorControl.v(20[7:21])
    defparam i4325_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4914));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11422_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n9613), .I3(GND_net), 
            .O(n25120));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4915));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_964 (.I0(n55139), .I1(PWMLimit[19]), .I2(n25120), 
            .I3(n9611), .O(n49[19]));
    defparam i1_4_lut_adj_964.LUT_INIT = 16'h5044;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4916));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11417_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n9613), .I3(GND_net), 
            .O(n25115));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24497_4_lut (.I0(PWMLimit[20]), .I1(n55139), .I2(n25115), 
            .I3(n9611), .O(n49[20]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24497_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i35_2_lut (.I0(PWMLimit[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4917));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4547));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11412_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n9613), .I3(GND_net), 
            .O(n25110));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24496_4_lut (.I0(PWMLimit[21]), .I1(n55139), .I2(n25110), 
            .I3(n9611), .O(n49[21]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24496_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11273_3_lut (.I0(n356[0]), .I1(n436[0]), .I2(n9613), .I3(GND_net), 
            .O(n24971));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11407_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n9613), .I3(GND_net), 
            .O(n25105));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24495_4_lut (.I0(PWMLimit[22]), .I1(n55139), .I2(n25105), 
            .I3(n9611), .O(n49[22]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24495_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4918));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i31_2_lut (.I0(PWMLimit[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4919));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44820_2_lut_4_lut (.I0(n356[11]), .I1(n436[11]), .I2(n356[7]), 
            .I3(n436[7]), .O(n59720));
    defparam i44820_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i11402_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n9613), .I3(GND_net), 
            .O(n25100));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24494_4_lut (.I0(PWMLimit[23]), .I1(n55139), .I2(n25100), 
            .I3(n9611), .O(n49[23]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i24494_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4920));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4921));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4922));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4923));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i45_2_lut (.I0(PWMLimit[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4924));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44692_2_lut_4_lut (.I0(n356[19]), .I1(n436[19]), .I2(n356[10]), 
            .I3(n436[10]), .O(n59592));
    defparam i44692_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4925));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[11]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4926));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45190_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n60090));
    defparam i45190_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4546));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45232_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n60132));
    defparam i45232_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4927));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4928));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31825_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n45395));   // verilog/motorControl.v(50[18:24])
    defparam i31825_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[12]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(counter[17]), .I1(counter[18]), .I2(counter[21]), 
            .I3(counter[22]), .O(n55117));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45000_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(PWMLimit[2]), .O(n59900));   // verilog/motorControl.v(52[14:29])
    defparam i45000_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_4929));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i5_2_lut (.I0(counter[26]), .I1(counter[15]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4930));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut (.I0(counter[25]), .I1(counter[16]), .I2(counter[19]), 
            .I3(counter[14]), .O(n26_adj_4931));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_4932));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[5]), .I1(n12_adj_4932), .I2(counter[2]), 
            .I3(counter[0]), .O(n55108));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4933));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44973_4_lut (.I0(n21_adj_4928), .I1(n19_adj_4925), .I2(n17_adj_4922), 
            .I3(n9_adj_4868), .O(n59873));
    defparam i44973_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i3_4_lut_adj_965 (.I0(counter[12]), .I1(n55108), .I2(counter[8]), 
            .I3(counter[7]), .O(n9_adj_4934));
    defparam i3_4_lut_adj_965.LUT_INIT = 16'ha8a0;
    SB_LUT4 i9_4_lut_adj_966 (.I0(counter[24]), .I1(counter[28]), .I2(counter[29]), 
            .I3(n55117), .O(n24_adj_4935));
    defparam i9_4_lut_adj_966.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(counter[30]), .I1(n26_adj_4931), .I2(n20_adj_4930), 
            .I3(counter[27]), .O(n28_adj_4936));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_967 (.I0(counter[20]), .I1(counter[23]), .I2(n9_adj_4934), 
            .I3(n10_adj_4933), .O(n23_adj_4937));
    defparam i8_4_lut_adj_967.LUT_INIT = 16'hfeee;
    SB_LUT4 i24460_4_lut (.I0(n23_adj_4937), .I1(counter[31]), .I2(n28_adj_4936), 
            .I3(n24_adj_4935), .O(counter_31__N_3690));   // verilog/motorControl.v(26[8:41])
    defparam i24460_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i44956_4_lut (.I0(n27_adj_4921), .I1(n15_adj_4877), .I2(n13_adj_4870), 
            .I3(n11_adj_2), .O(n59856));
    defparam i44956_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_4920), 
            .I3(GND_net), .O(n12_adj_4939));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n375), .I1(n356[6]), .I2(n13_adj_4870), 
            .I3(GND_net), .O(n10_adj_4940));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i30_3_lut (.I0(n12_adj_4939), .I1(n356[17]), .I2(n35_adj_4917), 
            .I3(GND_net), .O(n30_adj_4941));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31854_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[21] ), .I3(\Ki[1] ), 
            .O(n18242[0]));   // verilog/motorControl.v(50[27:38])
    defparam i31854_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i31856_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[21] ), .I3(\Ki[1] ), 
            .O(n45429));   // verilog/motorControl.v(50[27:38])
    defparam i31856_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i31671_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[20] ), .I3(\Ki[1] ), 
            .O(n18218[0]));   // verilog/motorControl.v(50[27:38])
    defparam i31671_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i31673_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[20] ), .I3(\Ki[1] ), 
            .O(n45231));   // verilog/motorControl.v(50[27:38])
    defparam i31673_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i45873_4_lut (.I0(n13_adj_4870), .I1(n11_adj_2), .I2(n9_adj_4868), 
            .I3(n59900), .O(n60773));
    defparam i45873_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_3_lut_4_lut_adj_968 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(n4_adj_4942), .I3(n18218[1]), .O(n18178[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_968.LUT_INIT = 16'h8778;
    SB_LUT4 i31730_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(n4_adj_4942), .I3(n18218[1]), .O(n6_adj_4912));   // verilog/motorControl.v(50[27:38])
    defparam i31730_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i45861_4_lut (.I0(n19_adj_4925), .I1(n17_adj_4922), .I2(n15_adj_4877), 
            .I3(n60773), .O(n60761));
    defparam i45861_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i31722_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(n45272), .I3(n18218[0]), .O(n4_adj_4942));   // verilog/motorControl.v(50[27:38])
    defparam i31722_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_969 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(n45272), .I3(n18218[0]), .O(n18178[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_969.LUT_INIT = 16'h8778;
    SB_LUT4 i31709_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[20] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[19] ), .I3(\Ki[1] ), 
            .O(n18178[0]));   // verilog/motorControl.v(50[27:38])
    defparam i31709_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i31711_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[20] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[19] ), .I3(\Ki[1] ), 
            .O(n45272));   // verilog/motorControl.v(50[27:38])
    defparam i31711_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i46939_4_lut (.I0(n25_adj_4923), .I1(n23_adj_4927), .I2(n21_adj_4928), 
            .I3(n60761), .O(n61839));
    defparam i46939_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31768_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I2(n4_adj_4943), .I3(n18178[1]), .O(n6_adj_4907));   // verilog/motorControl.v(50[27:38])
    defparam i31768_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_970 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I2(n4_adj_4943), .I3(n18178[1]), .O(n18118[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_970.LUT_INIT = 16'h8778;
    SB_LUT4 i46355_4_lut (.I0(n31_adj_4919), .I1(n29_adj_4918), .I2(n27_adj_4921), 
            .I3(n61839), .O(n61255));
    defparam i46355_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_4_lut_adj_971 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I2(n45313), .I3(n18178[0]), .O(n18118[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_971.LUT_INIT = 16'h8778;
    SB_LUT4 i47082_4_lut (.I0(n37_adj_4914), .I1(n35_adj_4917), .I2(n33_adj_4920), 
            .I3(n61255), .O(n61982));
    defparam i47082_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31760_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3691[18] ), 
            .I2(n45313), .I3(n18178[0]), .O(n4_adj_4943));   // verilog/motorControl.v(50[27:38])
    defparam i31760_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_4926), 
            .I3(GND_net), .O(n16_adj_4944));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31747_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[18] ), .I3(\Ki[1] ), 
            .O(n18118[0]));   // verilog/motorControl.v(50[27:38])
    defparam i31747_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31749_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[19] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3691[18] ), .I3(\Ki[1] ), 
            .O(n45313));   // verilog/motorControl.v(50[27:38])
    defparam i31749_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_2_lut_3_lut (.I0(n4), .I1(n3), .I2(\data_in_frame[10][4] ), 
            .I3(GND_net), .O(n23375));   // verilog/coms.v(99[12:25])
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i46600_3_lut (.I0(n6_adj_4929), .I1(n356[10]), .I2(n21_adj_4928), 
            .I3(GND_net), .O(n61500));   // verilog/motorControl.v(52[14:29])
    defparam i46600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_4_lut (.I0(\data_in_frame[10][4] ), .I1(n22_adj_4569), 
            .I2(n23824), .I3(n53055), .O(n25_adj_4572));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i46601_3_lut (.I0(n61500), .I1(n356[11]), .I2(n23_adj_4927), 
            .I3(GND_net), .O(n61501));   // verilog/motorControl.v(52[14:29])
    defparam i46601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4922), 
            .I3(GND_net), .O(n8_adj_4947));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n16_adj_4944), .I1(n356[22]), .I2(n45_adj_4924), 
            .I3(GND_net), .O(n24_adj_4948));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44896_4_lut (.I0(n43_adj_4926), .I1(n25_adj_4923), .I2(n23_adj_4927), 
            .I3(n59873), .O(n59796));
    defparam i44896_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46273_4_lut (.I0(n24_adj_4948), .I1(n8_adj_4947), .I2(n45_adj_4924), 
            .I3(n59794), .O(n61173));   // verilog/motorControl.v(52[14:29])
    defparam i46273_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45627_3_lut (.I0(n61501), .I1(n356[12]), .I2(n25_adj_4923), 
            .I3(GND_net), .O(n60527));   // verilog/motorControl.v(52[14:29])
    defparam i45627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45315_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n60215));
    defparam i45315_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i4_4_lut (.I0(PWMLimit[0]), .I1(n356[1]), .I2(PWMLimit[1]), 
            .I3(n356[0]), .O(n4_adj_4949));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i45377_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n60277));
    defparam i45377_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46598_3_lut (.I0(n4_adj_4949), .I1(n356[13]), .I2(n27_adj_4921), 
            .I3(GND_net), .O(n61498));   // verilog/motorControl.v(52[14:29])
    defparam i46598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4501));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31823_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n18202[0]));   // verilog/motorControl.v(50[18:24])
    defparam i31823_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i46599_3_lut (.I0(n61498), .I1(n356[14]), .I2(n29_adj_4918), 
            .I3(GND_net), .O(n61499));   // verilog/motorControl.v(52[14:29])
    defparam i46599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44941_4_lut (.I0(n33_adj_4920), .I1(n31_adj_4919), .I2(n29_adj_4918), 
            .I3(n59856), .O(n59841));
    defparam i44941_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45188_3_lut_4_lut (.I0(deadband[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(deadband[2]), .O(n60088));   // verilog/motorControl.v(51[12:29])
    defparam i45188_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_4432));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i46971_4_lut (.I0(n30_adj_4941), .I1(n10_adj_4940), .I2(n35_adj_4917), 
            .I3(n59834), .O(n61871));   // verilog/motorControl.v(52[14:29])
    defparam i46971_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4500));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45629_3_lut (.I0(n61499), .I1(n356[15]), .I2(n31_adj_4919), 
            .I3(GND_net), .O(n60529));   // verilog/motorControl.v(52[14:29])
    defparam i45629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47150_4_lut (.I0(n60529), .I1(n61871), .I2(n35_adj_4917), 
            .I3(n59841), .O(n62050));   // verilog/motorControl.v(52[14:29])
    defparam i47150_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47151_3_lut (.I0(n62050), .I1(n356[18]), .I2(n37_adj_4914), 
            .I3(GND_net), .O(n62051));   // verilog/motorControl.v(52[14:29])
    defparam i47151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47136_3_lut (.I0(n62051), .I1(n356[19]), .I2(n39_adj_4916), 
            .I3(GND_net), .O(n62036));   // verilog/motorControl.v(52[14:29])
    defparam i47136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44902_4_lut (.I0(n43_adj_4926), .I1(n41_adj_4915), .I2(n39_adj_4916), 
            .I3(n61982), .O(n59802));
    defparam i44902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46877_4_lut (.I0(n60527), .I1(n61173), .I2(n45_adj_4924), 
            .I3(n59796), .O(n61777));   // verilog/motorControl.v(52[14:29])
    defparam i46877_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45635_3_lut (.I0(n62036), .I1(n356[20]), .I2(n41_adj_4915), 
            .I3(GND_net), .O(n60535));   // verilog/motorControl.v(52[14:29])
    defparam i45635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4499));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_2_lut_4_lut (.I0(n47989), .I1(\data_in_frame[9][5] ), .I2(\data_in_frame[11][6] ), 
            .I3(n47452), .O(n16));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut_adj_972 (.I0(n47989), .I1(\data_in_frame[9][5] ), 
            .I2(\data_in_frame[11][6] ), .I3(n52878), .O(n12_adj_4578));
    defparam i3_2_lut_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47065_4_lut (.I0(n60535), .I1(n61777), .I2(n45_adj_4924), 
            .I3(n59802), .O(n61965));   // verilog/motorControl.v(52[14:29])
    defparam i47065_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44615_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n151), .I2(n152), 
            .I3(IntegralLimit[2]), .O(n59515));   // verilog/motorControl.v(45[12:34])
    defparam i44615_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n151), 
            .I2(n152), .I3(GND_net), .O(n6_adj_4543));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47066_3_lut (.I0(n61965), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(52[14:29])
    defparam i47066_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[23] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(deadband[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(deadband[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3691[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[22] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[21] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(deadband[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[20] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(deadband[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4414));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3691[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4498));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3691[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i4_4_lut_4_lut (.I0(n356[0]), .I1(n356[1]), .I2(n436[1]), 
            .I3(n436[0]), .O(n4_adj_4892));   // verilog/motorControl.v(50[18:38])
    defparam LessThan_25_i4_4_lut_4_lut.LUT_INIT = 16'h7130;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4517));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4516));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n207[19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i20_3_lut (.I0(n207[19]), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[19] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4497));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n207[18]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i19_3_lut (.I0(n207[18]), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[18] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20482_3_lut_4_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10][4] ), 
            .I2(Kp_23__N_1724), .I3(n30905), .O(n27611));
    defparam i20482_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3691[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4515));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4514));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45076_4_lut (.I0(n356[6]), .I1(n375), .I2(n382[6]), .I3(n382[5]), 
            .O(n59976));
    defparam i45076_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4495));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45949_3_lut (.I0(n356[7]), .I1(n59976), .I2(n382[7]), .I3(GND_net), 
            .O(n60849));
    defparam i45949_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i27_rep_108_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n62926));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i27_rep_108_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45919_4_lut (.I0(n356[14]), .I1(n62926), .I2(n382[14]), .I3(n60849), 
            .O(n60819));
    defparam i45919_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_102_2_lut (.I0(n356[15]), .I1(n382[15]), 
            .I2(GND_net), .I3(GND_net), .O(n62920));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i31_rep_102_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45068_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n59968));
    defparam i45068_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut_4_lut_adj_973 (.I0(\Kp[3] ), .I1(n1[19]), .I2(n18233[1]), 
            .I3(n4_adj_4901), .O(n18202[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_973.LUT_INIT = 16'h8778;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31844_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n4_adj_4901), 
            .I3(n18233[1]), .O(n6_adj_4409));   // verilog/motorControl.v(50[18:24])
    defparam i31844_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[9] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[8] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[5] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45939_3_lut (.I0(n356[9]), .I1(n59968), .I2(n382[9]), .I3(GND_net), 
            .O(n60839));
    defparam i45939_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i45931_4_lut (.I0(n356[11]), .I1(n62942), .I2(n382[11]), .I3(n60839), 
            .O(n60831));
    defparam i45931_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3691[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_4954));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45004_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n59904));
    defparam i45004_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mux_14_i3_3_lut (.I0(n152), .I1(n204), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3691[2] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8_adj_4493));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45089_2_lut_4_lut (.I0(deadband[21]), .I1(n356[21]), .I2(deadband[9]), 
            .I3(n356[9]), .O(n59989));
    defparam i45089_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_4954), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24_adj_4492));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45085_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n59985));
    defparam i45085_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i9_rep_116_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n62934));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i9_rep_116_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45083_4_lut (.I0(n375), .I1(n62934), .I2(n382[5]), .I3(n59985), 
            .O(n59983));
    defparam i45083_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i13_rep_144_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n62962));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i13_rep_144_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45129_2_lut_4_lut (.I0(deadband[16]), .I1(n356[16]), .I2(deadband[7]), 
            .I3(n356[7]), .O(n60029));
    defparam i45129_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46411_4_lut (.I0(n356[7]), .I1(n62962), .I2(n382[7]), .I3(n59983), 
            .O(n61311));
    defparam i46411_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i31806_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n45363), 
            .I3(n18250[0]), .O(n4_c));   // verilog/motorControl.v(50[18:24])
    defparam i31806_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4956[13]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_21_i17_rep_141_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n62959));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i17_rep_141_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_974 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n18250[0]), 
            .I3(n45363), .O(n18233[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_974.LUT_INIT = 16'h8778;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (b_prev, GND_net, a_new, position_31__N_3803, 
            ENCODER1_B_N_keep, n1884, ENCODER1_A_N_keep, n27009, n1889, 
            \encoder1_position[0] , \encoder1_position[1] , \encoder1_position[2] , 
            \encoder1_position[3] , \encoder1_position[4] , \encoder1_position[5] , 
            \encoder1_position[6] , \encoder1_position[7] , \encoder1_position[8] , 
            \encoder1_position[9] , \encoder1_position[10] , \encoder1_position[11] , 
            \encoder1_position[12] , \encoder1_position[13] , \encoder1_position[14] , 
            \encoder1_position[15] , \encoder1_position[16] , \encoder1_position[17] , 
            \encoder1_position[18] , \encoder1_position[19] , \encoder1_position[20] , 
            \encoder1_position[21] , \encoder1_position[22] , \encoder1_position[23] , 
            n1905, n1903, n1901, n1899, n1897, n1895, n1893, n1891, 
            VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output position_31__N_3803;
    input ENCODER1_B_N_keep;
    input n1884;
    input ENCODER1_A_N_keep;
    input n27009;
    output n1889;
    output \encoder1_position[0] ;
    output \encoder1_position[1] ;
    output \encoder1_position[2] ;
    output \encoder1_position[3] ;
    output \encoder1_position[4] ;
    output \encoder1_position[5] ;
    output \encoder1_position[6] ;
    output \encoder1_position[7] ;
    output \encoder1_position[8] ;
    output \encoder1_position[9] ;
    output \encoder1_position[10] ;
    output \encoder1_position[11] ;
    output \encoder1_position[12] ;
    output \encoder1_position[13] ;
    output \encoder1_position[14] ;
    output \encoder1_position[15] ;
    output \encoder1_position[16] ;
    output \encoder1_position[17] ;
    output \encoder1_position[18] ;
    output \encoder1_position[19] ;
    output \encoder1_position[20] ;
    output \encoder1_position[21] ;
    output \encoder1_position[22] ;
    output \encoder1_position[23] ;
    output n1905;
    output n1903;
    output n1901;
    output n1899;
    output n1897;
    output n1895;
    output n1893;
    output n1891;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_3806, debounce_cnt, a_prev, direction_N_3808;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3811, n27008, n27004;
    wire [31:0]n133;
    
    wire n46229, n46228, n46227, n46226, n46225, n46224, n46223, 
        n46222, n46221, n46220, n46219, n46218, n46217, n46216, 
        n46215, n46214, n46213, n46212, n46211, n46210, n46209, 
        n46208, n46207, n46206, n46205, n46204, n46203, n46202, 
        n46201, n46200, n46199;
    
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3806));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3806), 
            .I3(a_new[1]), .O(position_31__N_3803));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3808));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i47316_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3811));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i47316_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1884), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1884), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1884), .D(a_prev_N_3811));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1889), .C(n1884), .D(n27009));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1884), .D(n27008));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1884), .D(n27004));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1936__i0 (.Q(\encoder1_position[0] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1884), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1884), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1936__i1 (.Q(\encoder1_position[1] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i2 (.Q(\encoder1_position[2] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i3 (.Q(\encoder1_position[3] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i4 (.Q(\encoder1_position[4] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i5 (.Q(\encoder1_position[5] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i6 (.Q(\encoder1_position[6] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i7 (.Q(\encoder1_position[7] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i8 (.Q(\encoder1_position[8] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i9 (.Q(\encoder1_position[9] ), .C(n1884), .E(position_31__N_3803), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i10 (.Q(\encoder1_position[10] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i11 (.Q(\encoder1_position[11] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i12 (.Q(\encoder1_position[12] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i13 (.Q(\encoder1_position[13] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i14 (.Q(\encoder1_position[14] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i15 (.Q(\encoder1_position[15] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i16 (.Q(\encoder1_position[16] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i17 (.Q(\encoder1_position[17] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i18 (.Q(\encoder1_position[18] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i19 (.Q(\encoder1_position[19] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i20 (.Q(\encoder1_position[20] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i21 (.Q(\encoder1_position[21] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i22 (.Q(\encoder1_position[22] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i23 (.Q(\encoder1_position[23] ), .C(n1884), 
            .E(position_31__N_3803), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i24 (.Q(n1905), .C(n1884), .E(position_31__N_3803), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i25 (.Q(n1903), .C(n1884), .E(position_31__N_3803), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i26 (.Q(n1901), .C(n1884), .E(position_31__N_3803), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i27 (.Q(n1899), .C(n1884), .E(position_31__N_3803), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i28 (.Q(n1897), .C(n1884), .E(position_31__N_3803), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i29 (.Q(n1895), .C(n1884), .E(position_31__N_3803), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i30 (.Q(n1893), .C(n1884), .E(position_31__N_3803), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i31 (.Q(n1891), .C(n1884), .E(position_31__N_3803), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1936_add_4_33_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1891), .I3(n46229), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1936_add_4_32_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1893), .I3(n46228), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_32 (.CI(n46228), .I0(direction_N_3808), 
            .I1(n1893), .CO(n46229));
    SB_LUT4 position_1936_add_4_31_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1895), .I3(n46227), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_31 (.CI(n46227), .I0(direction_N_3808), 
            .I1(n1895), .CO(n46228));
    SB_LUT4 position_1936_add_4_30_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1897), .I3(n46226), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_30 (.CI(n46226), .I0(direction_N_3808), 
            .I1(n1897), .CO(n46227));
    SB_LUT4 position_1936_add_4_29_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1899), .I3(n46225), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_29 (.CI(n46225), .I0(direction_N_3808), 
            .I1(n1899), .CO(n46226));
    SB_LUT4 position_1936_add_4_28_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1901), .I3(n46224), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_28 (.CI(n46224), .I0(direction_N_3808), 
            .I1(n1901), .CO(n46225));
    SB_LUT4 position_1936_add_4_27_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1903), .I3(n46223), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_27 (.CI(n46223), .I0(direction_N_3808), 
            .I1(n1903), .CO(n46224));
    SB_LUT4 position_1936_add_4_26_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(n1905), .I3(n46222), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_26 (.CI(n46222), .I0(direction_N_3808), 
            .I1(n1905), .CO(n46223));
    SB_LUT4 position_1936_add_4_25_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[23] ), .I3(n46221), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_25 (.CI(n46221), .I0(direction_N_3808), 
            .I1(\encoder1_position[23] ), .CO(n46222));
    SB_LUT4 position_1936_add_4_24_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[22] ), .I3(n46220), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_24 (.CI(n46220), .I0(direction_N_3808), 
            .I1(\encoder1_position[22] ), .CO(n46221));
    SB_LUT4 position_1936_add_4_23_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[21] ), .I3(n46219), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_23 (.CI(n46219), .I0(direction_N_3808), 
            .I1(\encoder1_position[21] ), .CO(n46220));
    SB_LUT4 position_1936_add_4_22_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[20] ), .I3(n46218), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_22 (.CI(n46218), .I0(direction_N_3808), 
            .I1(\encoder1_position[20] ), .CO(n46219));
    SB_LUT4 position_1936_add_4_21_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[19] ), .I3(n46217), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_21 (.CI(n46217), .I0(direction_N_3808), 
            .I1(\encoder1_position[19] ), .CO(n46218));
    SB_LUT4 position_1936_add_4_20_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[18] ), .I3(n46216), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_20 (.CI(n46216), .I0(direction_N_3808), 
            .I1(\encoder1_position[18] ), .CO(n46217));
    SB_LUT4 position_1936_add_4_19_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[17] ), .I3(n46215), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_19 (.CI(n46215), .I0(direction_N_3808), 
            .I1(\encoder1_position[17] ), .CO(n46216));
    SB_LUT4 position_1936_add_4_18_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[16] ), .I3(n46214), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_18 (.CI(n46214), .I0(direction_N_3808), 
            .I1(\encoder1_position[16] ), .CO(n46215));
    SB_LUT4 position_1936_add_4_17_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[15] ), .I3(n46213), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_17 (.CI(n46213), .I0(direction_N_3808), 
            .I1(\encoder1_position[15] ), .CO(n46214));
    SB_LUT4 position_1936_add_4_16_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[14] ), .I3(n46212), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_16 (.CI(n46212), .I0(direction_N_3808), 
            .I1(\encoder1_position[14] ), .CO(n46213));
    SB_LUT4 position_1936_add_4_15_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[13] ), .I3(n46211), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_15 (.CI(n46211), .I0(direction_N_3808), 
            .I1(\encoder1_position[13] ), .CO(n46212));
    SB_LUT4 position_1936_add_4_14_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[12] ), .I3(n46210), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_14 (.CI(n46210), .I0(direction_N_3808), 
            .I1(\encoder1_position[12] ), .CO(n46211));
    SB_LUT4 position_1936_add_4_13_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[11] ), .I3(n46209), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_13 (.CI(n46209), .I0(direction_N_3808), 
            .I1(\encoder1_position[11] ), .CO(n46210));
    SB_LUT4 position_1936_add_4_12_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[10] ), .I3(n46208), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_12 (.CI(n46208), .I0(direction_N_3808), 
            .I1(\encoder1_position[10] ), .CO(n46209));
    SB_LUT4 position_1936_add_4_11_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[9] ), .I3(n46207), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_11 (.CI(n46207), .I0(direction_N_3808), 
            .I1(\encoder1_position[9] ), .CO(n46208));
    SB_LUT4 position_1936_add_4_10_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[8] ), .I3(n46206), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_10 (.CI(n46206), .I0(direction_N_3808), 
            .I1(\encoder1_position[8] ), .CO(n46207));
    SB_LUT4 position_1936_add_4_9_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[7] ), .I3(n46205), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_9 (.CI(n46205), .I0(direction_N_3808), 
            .I1(\encoder1_position[7] ), .CO(n46206));
    SB_LUT4 position_1936_add_4_8_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[6] ), .I3(n46204), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_8 (.CI(n46204), .I0(direction_N_3808), 
            .I1(\encoder1_position[6] ), .CO(n46205));
    SB_LUT4 position_1936_add_4_7_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[5] ), .I3(n46203), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_7 (.CI(n46203), .I0(direction_N_3808), 
            .I1(\encoder1_position[5] ), .CO(n46204));
    SB_LUT4 position_1936_add_4_6_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[4] ), .I3(n46202), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_6 (.CI(n46202), .I0(direction_N_3808), 
            .I1(\encoder1_position[4] ), .CO(n46203));
    SB_LUT4 position_1936_add_4_5_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[3] ), .I3(n46201), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_5 (.CI(n46201), .I0(direction_N_3808), 
            .I1(\encoder1_position[3] ), .CO(n46202));
    SB_LUT4 position_1936_add_4_4_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[2] ), .I3(n46200), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_4 (.CI(n46200), .I0(direction_N_3808), 
            .I1(\encoder1_position[2] ), .CO(n46201));
    SB_LUT4 position_1936_add_4_3_lut (.I0(GND_net), .I1(direction_N_3808), 
            .I2(\encoder1_position[1] ), .I3(n46199), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_3 (.CI(n46199), .I0(direction_N_3808), 
            .I1(\encoder1_position[1] ), .CO(n46200));
    SB_LUT4 position_1936_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder1_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder1_position[0] ), 
            .CO(n46199));
    SB_LUT4 i13302_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3811), .I2(b_new[1]), 
            .I3(b_prev), .O(n27008));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13302_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13298_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3811), .I2(a_new[1]), 
            .I3(a_prev), .O(n27004));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13298_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2978, pwm_out, clk32MHz, pwm_setpoint, GND_net, reset, 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input n2978;
    output pwm_out;
    input clk32MHz;
    input [23:0]pwm_setpoint;
    input GND_net;
    input reset;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_553;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n41, n39, n45, n37, n43, n29, n31, n23, n25, n35, 
        n33, n9, n17, n19, n21, n11, n13, n15, n27, n59964, 
        n59922, n12, n30, n60053, n60915, n60903, n61879, n61285, 
        n61996, n6, n61593, n61594, n16, n24, n59863, n8, n59851, 
        n61147, n60469, n4, n61597, n61598, n59907, n10, n59898, 
        n61945, n60465, n62083, n62084, n62005, n59867, n61755, 
        n61457, n61951, n51903, n51911, n51913, n51915, n51771, 
        n51651, n51573, n51519, n51477, n51445, n51407, n51373, 
        n51347, n51321, n51283, n51213, n51177, n51155, n51123, 
        n51101, n51081, n51061, n51041, n51019, n46098, n48, n46097, 
        n46096, n46095, n46094, n46093, n46092, n46091, n46090, 
        n46089, n46088, n46087, n46086, n46085, n46084, n46083, 
        n46082, n46081, n46080, n46079, n46078, n46077, n46076, 
        n54830, n22, n15_adj_4404, n20, n24_adj_4405, n19_adj_4406;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2978), .D(pwm_out_N_553));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45064_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n59964));
    defparam i45064_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45022_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n59922));
    defparam i45022_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46015_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n60053), 
            .O(n60915));
    defparam i46015_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46003_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n60915), 
            .O(n60903));
    defparam i46003_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46979_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n60903), 
            .O(n61879));
    defparam i46979_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46385_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n61879), 
            .O(n61285));
    defparam i46385_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47096_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n61285), 
            .O(n61996));
    defparam i47096_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46693_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n61593));   // verilog/pwm.v(21[8:24])
    defparam i46693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46694_3_lut (.I0(n61593), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n61594));   // verilog/pwm.v(21[8:24])
    defparam i46694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44963_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n59964), 
            .O(n59863));
    defparam i44963_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46247_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n59851), 
            .O(n61147));   // verilog/pwm.v(21[8:24])
    defparam i46247_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45569_3_lut (.I0(n61594), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n60469));   // verilog/pwm.v(21[8:24])
    defparam i45569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i46697_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n61597));   // verilog/pwm.v(21[8:24])
    defparam i46697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46698_3_lut (.I0(n61597), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n61598));   // verilog/pwm.v(21[8:24])
    defparam i46698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45007_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n59922), 
            .O(n59907));
    defparam i45007_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47045_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n59898), 
            .O(n61945));   // verilog/pwm.v(21[8:24])
    defparam i47045_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45565_3_lut (.I0(n61598), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n60465));   // verilog/pwm.v(21[8:24])
    defparam i45565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47183_4_lut (.I0(n60465), .I1(n61945), .I2(n35), .I3(n59907), 
            .O(n62083));   // verilog/pwm.v(21[8:24])
    defparam i47183_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47184_3_lut (.I0(n62083), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n62084));   // verilog/pwm.v(21[8:24])
    defparam i47184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47105_3_lut (.I0(n62084), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n62005));   // verilog/pwm.v(21[8:24])
    defparam i47105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44967_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n61996), 
            .O(n59867));
    defparam i44967_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46855_4_lut (.I0(n60469), .I1(n61147), .I2(n45), .I3(n59863), 
            .O(n61755));   // verilog/pwm.v(21[8:24])
    defparam i46855_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46557_3_lut (.I0(n62005), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n61457));   // verilog/pwm.v(21[8:24])
    defparam i46557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47051_4_lut (.I0(n61457), .I1(n61755), .I2(n45), .I3(n59867), 
            .O(n61951));   // verilog/pwm.v(21[8:24])
    defparam i47051_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47052_3_lut (.I0(n61951), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_553));   // verilog/pwm.v(21[8:24])
    defparam i47052_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR pwm_counter_1930__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n51903), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n51911), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n51913), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n51915), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n51771), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n51651), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n51573), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n51519), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n51477), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n51445), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n51407), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n51373), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n51347), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n51321), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n51283), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n51213), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n51177), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n51155), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n51123), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n51101), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n51081), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n51061), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n51041), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1930__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n51019), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1930_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n46098), .O(n51019)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1930_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n46097), .O(n51041)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_24 (.CI(n46097), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n46098));
    SB_LUT4 pwm_counter_1930_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n46096), .O(n51061)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_23 (.CI(n46096), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n46097));
    SB_LUT4 pwm_counter_1930_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n46095), .O(n51081)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_22 (.CI(n46095), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n46096));
    SB_LUT4 pwm_counter_1930_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n46094), .O(n51101)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_21 (.CI(n46094), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n46095));
    SB_LUT4 pwm_counter_1930_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n46093), .O(n51123)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_20 (.CI(n46093), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n46094));
    SB_LUT4 pwm_counter_1930_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n46092), .O(n51155)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_19 (.CI(n46092), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n46093));
    SB_LUT4 pwm_counter_1930_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n46091), .O(n51177)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_18 (.CI(n46091), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n46092));
    SB_LUT4 pwm_counter_1930_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n46090), .O(n51213)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_17 (.CI(n46090), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n46091));
    SB_LUT4 pwm_counter_1930_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n46089), .O(n51283)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_16 (.CI(n46089), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n46090));
    SB_LUT4 pwm_counter_1930_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n46088), .O(n51321)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_15 (.CI(n46088), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n46089));
    SB_LUT4 pwm_counter_1930_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n46087), .O(n51347)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_14 (.CI(n46087), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n46088));
    SB_LUT4 pwm_counter_1930_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n46086), .O(n51373)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_13 (.CI(n46086), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n46087));
    SB_LUT4 pwm_counter_1930_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n46085), .O(n51407)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_12 (.CI(n46085), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n46086));
    SB_LUT4 pwm_counter_1930_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n46084), .O(n51445)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_11 (.CI(n46084), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n46085));
    SB_LUT4 pwm_counter_1930_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n46083), .O(n51477)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_10 (.CI(n46083), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n46084));
    SB_LUT4 pwm_counter_1930_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n46082), .O(n51519)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_9 (.CI(n46082), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n46083));
    SB_LUT4 pwm_counter_1930_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n46081), .O(n51573)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_8 (.CI(n46081), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n46082));
    SB_LUT4 pwm_counter_1930_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n46080), .O(n51651)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_7 (.CI(n46080), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n46081));
    SB_LUT4 pwm_counter_1930_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n46079), .O(n51771)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_6 (.CI(n46079), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n46080));
    SB_LUT4 pwm_counter_1930_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n46078), .O(n51915)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_5 (.CI(n46078), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n46079));
    SB_LUT4 pwm_counter_1930_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n46077), .O(n51913)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_4 (.CI(n46077), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n46078));
    SB_LUT4 pwm_counter_1930_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n46076), .O(n51911)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_3 (.CI(n46076), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n46077));
    SB_LUT4 pwm_counter_1930_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n51903)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1930_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1930_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n46076));
    SB_LUT4 i45153_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n60053));   // verilog/pwm.v(21[8:24])
    defparam i45153_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n54830));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[15]), .I1(pwm_counter[16]), .I2(pwm_counter[20]), 
            .I3(pwm_counter[19]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n54830), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4404));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[13]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4404), .I1(n22), .I2(pwm_counter[22]), 
            .I3(pwm_counter[18]), .O(n24_adj_4405));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[14]), .I1(pwm_counter[17]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4406));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4406), .I2(n24_adj_4405), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44951_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n59851));
    defparam i44951_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44998_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n59898));
    defparam i44998_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
